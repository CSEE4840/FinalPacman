0000
0000
0c30
1c1c
1e3c
3e3e
3f7e
3ffe
3ffe
1ffc
1ffc
0ff8
03e0
0000
0000
