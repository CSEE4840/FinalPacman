0F
30
40
47
88
90
90
90
FF
00
00
FF
00
00
00
00
FF
00
00
E0
10
08
08
08
FF
00
00
07
08
10
10
10
F0
0C
02
E2
11
09
09
09
09
09
09
11
E2
02
0C
F0
00
00
00
00
FF
00
00
00
00
00
00
07
08
10
10
10
00
00
00
E0
10
08
08
08
90
90
90
90
90
90
90
90
00
00
00
18
18
00
00
00
08
08
08
08
08
08
08
08
10
10
10
10
10
10
10
10
09
09
09
09
09
09
09
09
09
09
09
11
E1
01
01
01
90
90
90
88
87
80
80
80
00
00
00
FF
00
00
00
00
10
10
10
08
07
00
00
00
08
08
08
10
E0
00
00
00
90
90
90
88
47
40
30
0F
3C
7E
FF
FF
FF
FF
7E
3C
08
08
08
04
03
00
00
00
10
10
10
20
C0
00
00
00
00
00
00
00
0F
08
08
09
00
00
00
00
FF
01
01
FF
00
00
00
00
FF
80
80
FF
00
00
00
00
F0
10
10
90
00
00
00
00
03
04
08
08
00
00
00
00
FF
00
00
FF
00
00
00
00
C0
20
10
10
09
08
08
0F
00
00
00
00
00
00
00
00
00
FF
FF
00
90
10
10
F0
00
00
00
00
08
08
04
03
00
00
00
00
10
10
20
C0
00
00
00
00
80
80
80
87
88
90
90
90
01
01
01
E1
11
09
09
09
00
00
00
00
00
00
00
00
18
3C
66
C3
C3
FF
C3
C3
C3
C3
00
00
00
00
00
00
FE
66
66
66
7C
66
66
66
66
FE
00
00
00
00
00
00
3C
66
C2
C0
C0
C0
C0
C2
66
3C
00
00
00
00
00
00
FC
66
63
63
63
63
63
63
66
FC
00
00
00
00
00
00
FF
63
68
68
78
68
68
60
63
FF
00
00
00
00
00
00
FF
63
68
68
78
68
68
60
60
F0
00
00
00
00
00
00
3C
66
C2
C0
C0
CF
C3
C3
66
3C
00
00
00
00
00
00
C3
C3
C3
C3
FF
C3
C3
C3
C3
C3
00
00
00
00
00
00
3C
18
18
18
18
18
18
18
18
3C
00
00
00
00
00
00
1F
0C
0C
0C
0C
0C
CC
CC
78
30
00
00
00
00
00
00
E7
66
6C
78
70
78
6C
66
66
E7
00
00
00
00
00
00
F0
60
60
60
60
60
63
63
63
FF
00
00
00
00
00
00
C3
E7
FF
DB
C3
C3
C3
C3
C3
C3
00
00
00
00
00
00
C3
E3
F3
DB
CF
C7
C3
C3
C3
C3
00
00
00
00
00
00
3C
66
C3
C3
C3
C3
C3
C3
66
3C
00
00
00
00
00
00
FE
66
66
66
7E
60
60
60
60
F0
00
00
00
00
00
00
3C
66
C3
C3
C3
C3
CB
C7
66
3F
00
00
00
00
00
00
FE
66
66
66
7C
78
6C
66
66
E7
00
00
00
00
00
00
3E
66
C0
C0
7C
06
03
C3
66
3C
00
00
00
00
00
00
FF
DB
99
18
18
18
18
18
18
3C
00
00
00
00
00
00
C3
C3
C3
C3
C3
C3
C3
C3
66
3C
00
00
00
00
00
00
C3
C3
C3
C3
C3
C3
66
3C
18
18
00
00
00
00
00
00
C3
C3
C3
C3
C3
DB
FF
E7
C3
C3
00
00
00
00
00
00
C3
66
3C
18
18
3C
66
C3
C3
C3
00
00
00
00
00
00
C3
C3
66
3C
18
18
18
18
18
3C
00
00
00
00
00
00
FF
06
0C
18
30
60
C0
C0
C3
FF
00
00
00
00
00
00
3C
66
C3
C7
CF
DB
E3
C3
66
3C
00
00
00
00
00
00
18
38
78
18
18
18
18
18
18
7E
00
00
00
00
00
00
3C
66
C3
03
06
0C
18
30
60
FF
00
00
00
00
00
00
3C
66
C3
03
1E
03
03
C3
66
3C
00
00
00
00
00
00
06
0E
1E
36
66
FF
06
06
06
0F
00
00
00
00
00
00
FF
C0
C0
FC
06
03
03
C3
66
3C
00
00
00
00
00
00
3C
66
C0
C0
FC
C3
C3
C3
66
3C
00
00
00
00
00
00
FF
03
06
0C
18
30
60
60
60
60
00
00
00
00
00
00
3C
66
C3
66
3C
66
C3
C3
66
3C
00
00
00
00
00
00
3C
66
C3
C3
67
3F
03
03
66
3C
00
00
00
00
00
00
