    tile[0] = 6'd37;
    tile[1] = 6'd37;
    tile[2] = 6'd37;
    tile[3] = 6'd37;
    tile[4] = 6'd37;
    tile[5] = 6'd37;
    tile[6] = 6'd37;
    tile[7] = 6'd37;
    tile[8] = 6'd37;
    tile[9] = 6'd37;
    tile[10] = 6'd37;
    tile[11] = 6'd37;
    tile[12] = 6'd37;
    tile[13] = 6'd37;
    tile[14] = 6'd37;
    tile[15] = 6'd37;
    tile[16] = 6'd37;
    tile[17] = 6'd37;
    tile[18] = 6'd37;
    tile[19] = 6'd37;
    tile[20] = 6'd37;
    tile[21] = 6'd37;
    tile[22] = 6'd37;
    tile[23] = 6'd37;
    tile[24] = 6'd37;
    tile[25] = 6'd37;
    tile[26] = 6'd37;
    tile[27] = 6'd37;
    tile[28] = 6'd37;
    tile[29] = 6'd37;
    tile[30] = 6'd37;
    tile[31] = 6'd37;
    tile[32] = 6'd37;
    tile[33] = 6'd37;
    tile[34] = 6'd37;
    tile[35] = 6'd37;
    tile[36] = 6'd37;
    tile[37] = 6'd37;
    tile[38] = 6'd37;
    tile[39] = 6'd37;
    tile[40] = 6'd37;
    tile[41] = 6'd37;
    tile[42] = 6'd37;
    tile[43] = 6'd37;
    tile[44] = 6'd37;
    tile[45] = 6'd37;
    tile[46] = 6'd37;
    tile[47] = 6'd37;
    tile[48] = 6'd37;
    tile[49] = 6'd37;
    tile[50] = 6'd37;
    tile[51] = 6'd37;
    tile[52] = 6'd37;
    tile[53] = 6'd37;
    tile[54] = 6'd37;
    tile[55] = 6'd37;
    tile[56] = 6'd37;
    tile[57] = 6'd37;
    tile[58] = 6'd37;
    tile[59] = 6'd37;
    tile[60] = 6'd37;
    tile[61] = 6'd37;
    tile[62] = 6'd37;
    tile[63] = 6'd37;
    tile[64] = 6'd37;
    tile[65] = 6'd37;
    tile[66] = 6'd37;
    tile[67] = 6'd37;
    tile[68] = 6'd37;
    tile[69] = 6'd37;
    tile[70] = 6'd37;
    tile[71] = 6'd37;
    tile[72] = 6'd37;
    tile[73] = 6'd37;
    tile[74] = 6'd37;
    tile[75] = 6'd37;
    tile[76] = 6'd37;
    tile[77] = 6'd37;
    tile[78] = 6'd37;
    tile[79] = 6'd37;
    tile[80] = 6'd37;
    tile[81] = 6'd37;
    tile[82] = 6'd37;
    tile[83] = 6'd37;
    tile[84] = 6'd37;
    tile[85] = 6'd37;
    tile[86] = 6'd37;
    tile[87] = 6'd37;
    tile[88] = 6'd37;
    tile[89] = 6'd37;
    tile[90] = 6'd37;
    tile[91] = 6'd37;
    tile[92] = 6'd37;
    tile[93] = 6'd37;
    tile[94] = 6'd37;
    tile[95] = 6'd37;
    tile[96] = 6'd37;
    tile[97] = 6'd37;
    tile[98] = 6'd37;
    tile[99] = 6'd37;
    tile[100] = 6'd37;
    tile[101] = 6'd37;
    tile[102] = 6'd37;
    tile[103] = 6'd37;
    tile[104] = 6'd37;
    tile[105] = 6'd37;
    tile[106] = 6'd37;
    tile[107] = 6'd37;
    tile[108] = 6'd37;
    tile[109] = 6'd37;
    tile[110] = 6'd37;
    tile[111] = 6'd37;
    tile[112] = 6'd37;
    tile[113] = 6'd37;
    tile[114] = 6'd37;
    tile[115] = 6'd37;
    tile[116] = 6'd37;
    tile[117] = 6'd37;
    tile[118] = 6'd37;
    tile[119] = 6'd37;
    tile[120] = 6'd37;
    tile[121] = 6'd37;
    tile[122] = 6'd37;
    tile[123] = 6'd37;
    tile[124] = 6'd37;
    tile[125] = 6'd37;
    tile[126] = 6'd37;
    tile[127] = 6'd37;
    tile[128] = 6'd37;
    tile[129] = 6'd37;
    tile[130] = 6'd37;
    tile[131] = 6'd37;
    tile[132] = 6'd37;
    tile[133] = 6'd37;
    tile[134] = 6'd37;
    tile[135] = 6'd37;
    tile[136] = 6'd37;
    tile[137] = 6'd37;
    tile[138] = 6'd37;
    tile[139] = 6'd37;
    tile[140] = 6'd37;
    tile[141] = 6'd37;
    tile[142] = 6'd37;
    tile[143] = 6'd37;
    tile[144] = 6'd37;
    tile[145] = 6'd37;
    tile[146] = 6'd37;
    tile[147] = 6'd37;
    tile[148] = 6'd37;
    tile[149] = 6'd37;
    tile[150] = 6'd37;
    tile[151] = 6'd37;
    tile[152] = 6'd37;
    tile[153] = 6'd37;
    tile[154] = 6'd37;
    tile[155] = 6'd37;
    tile[156] = 6'd37;
    tile[157] = 6'd37;
    tile[158] = 6'd37;
    tile[159] = 6'd37;
    tile[160] = 6'd37;
    tile[161] = 6'd37;
    tile[162] = 6'd37;
    tile[163] = 6'd37;
    tile[164] = 6'd37;
    tile[165] = 6'd37;
    tile[166] = 6'd37;
    tile[167] = 6'd37;
    tile[168] = 6'd37;
    tile[169] = 6'd37;
    tile[170] = 6'd37;
    tile[171] = 6'd37;
    tile[172] = 6'd37;
    tile[173] = 6'd37;
    tile[174] = 6'd37;
    tile[175] = 6'd37;
    tile[176] = 6'd37;
    tile[177] = 6'd37;
    tile[178] = 6'd37;
    tile[179] = 6'd37;
    tile[180] = 6'd37;
    tile[181] = 6'd37;
    tile[182] = 6'd37;
    tile[183] = 6'd37;
    tile[184] = 6'd37;
    tile[185] = 6'd37;
    tile[186] = 6'd37;
    tile[187] = 6'd37;
    tile[188] = 6'd37;
    tile[189] = 6'd37;
    tile[190] = 6'd37;
    tile[191] = 6'd37;
    tile[192] = 6'd37;
    tile[193] = 6'd37;
    tile[194] = 6'd37;
    tile[195] = 6'd37;
    tile[196] = 6'd37;
    tile[197] = 6'd37;
    tile[198] = 6'd37;
    tile[199] = 6'd37;
    tile[200] = 6'd37;
    tile[201] = 6'd37;
    tile[202] = 6'd37;
    tile[203] = 6'd37;
    tile[204] = 6'd37;
    tile[205] = 6'd37;
    tile[206] = 6'd37;
    tile[207] = 6'd37;
    tile[208] = 6'd37;
    tile[209] = 6'd37;
    tile[210] = 6'd37;
    tile[211] = 6'd37;
    tile[212] = 6'd37;
    tile[213] = 6'd37;
    tile[214] = 6'd37;
    tile[215] = 6'd37;
    tile[216] = 6'd37;
    tile[217] = 6'd37;
    tile[218] = 6'd37;
    tile[219] = 6'd37;
    tile[220] = 6'd37;
    tile[221] = 6'd37;
    tile[222] = 6'd37;
    tile[223] = 6'd37;
    tile[224] = 6'd37;
    tile[225] = 6'd37;
    tile[226] = 6'd37;
    tile[227] = 6'd37;
    tile[228] = 6'd37;
    tile[229] = 6'd37;
    tile[230] = 6'd37;
    tile[231] = 6'd37;
    tile[232] = 6'd37;
    tile[233] = 6'd37;
    tile[234] = 6'd37;
    tile[235] = 6'd37;
    tile[236] = 6'd37;
    tile[237] = 6'd37;
    tile[238] = 6'd37;
    tile[239] = 6'd37;
    tile[240] = 6'd37;
    tile[241] = 6'd37;
    tile[242] = 6'd37;
    tile[243] = 6'd37;
    tile[244] = 6'd37;
    tile[245] = 6'd37;
    tile[246] = 6'd37;
    tile[247] = 6'd37;
    tile[248] = 6'd37;
    tile[249] = 6'd37;
    tile[250] = 6'd37;
    tile[251] = 6'd37;
    tile[252] = 6'd37;
    tile[253] = 6'd37;
    tile[254] = 6'd37;
    tile[255] = 6'd37;
    tile[256] = 6'd37;
    tile[257] = 6'd37;
    tile[258] = 6'd37;
    tile[259] = 6'd37;
    tile[260] = 6'd37;
    tile[261] = 6'd37;
    tile[262] = 6'd37;
    tile[263] = 6'd37;
    tile[264] = 6'd37;
    tile[265] = 6'd37;
    tile[266] = 6'd37;
    tile[267] = 6'd37;
    tile[268] = 6'd37;
    tile[269] = 6'd37;
    tile[270] = 6'd37;
    tile[271] = 6'd37;
    tile[272] = 6'd37;
    tile[273] = 6'd37;
    tile[274] = 6'd37;
    tile[275] = 6'd37;
    tile[276] = 6'd37;
    tile[277] = 6'd37;
    tile[278] = 6'd37;
    tile[279] = 6'd37;
    tile[280] = 6'd37;
    tile[281] = 6'd37;
    tile[282] = 6'd37;
    tile[283] = 6'd37;
    tile[284] = 6'd37;
    tile[285] = 6'd37;
    tile[286] = 6'd37;
    tile[287] = 6'd37;
    tile[288] = 6'd37;
    tile[289] = 6'd37;
    tile[290] = 6'd37;
    tile[291] = 6'd37;
    tile[292] = 6'd37;
    tile[293] = 6'd37;
    tile[294] = 6'd37;
    tile[295] = 6'd37;
    tile[296] = 6'd37;
    tile[297] = 6'd37;
    tile[298] = 6'd37;
    tile[299] = 6'd37;
    tile[300] = 6'd37;
    tile[301] = 6'd37;
    tile[302] = 6'd37;
    tile[303] = 6'd37;
    tile[304] = 6'd37;
    tile[305] = 6'd37;
    tile[306] = 6'd37;
    tile[307] = 6'd37;
    tile[308] = 6'd37;
    tile[309] = 6'd37;
    tile[310] = 6'd37;
    tile[311] = 6'd37;
    tile[312] = 6'd37;
    tile[313] = 6'd37;
    tile[314] = 6'd37;
    tile[315] = 6'd37;
    tile[316] = 6'd37;
    tile[317] = 6'd37;
    tile[318] = 6'd37;
    tile[319] = 6'd37;
    tile[320] = 6'd37;
    tile[321] = 6'd37;
    tile[322] = 6'd37;
    tile[323] = 6'd37;
    tile[324] = 6'd37;
    tile[325] = 6'd37;
    tile[326] = 6'd37;
    tile[327] = 6'd37;
    tile[328] = 6'd37;
    tile[329] = 6'd37;
    tile[330] = 6'd37;
    tile[331] = 6'd37;
    tile[332] = 6'd37;
    tile[333] = 6'd37;
    tile[334] = 6'd37;
    tile[335] = 6'd37;
    tile[336] = 6'd37;
    tile[337] = 6'd37;
    tile[338] = 6'd37;
    tile[339] = 6'd37;
    tile[340] = 6'd37;
    tile[341] = 6'd37;
    tile[342] = 6'd37;
    tile[343] = 6'd37;
    tile[344] = 6'd37;
    tile[345] = 6'd37;
    tile[346] = 6'd37;
    tile[347] = 6'd37;
    tile[348] = 6'd37;
    tile[349] = 6'd37;
    tile[350] = 6'd37;
    tile[351] = 6'd37;
    tile[352] = 6'd37;
    tile[353] = 6'd37;
    tile[354] = 6'd37;
    tile[355] = 6'd37;
    tile[356] = 6'd37;
    tile[357] = 6'd37;
    tile[358] = 6'd37;
    tile[359] = 6'd37;
    tile[360] = 6'd37;
    tile[361] = 6'd37;
    tile[362] = 6'd37;
    tile[363] = 6'd37;
    tile[364] = 6'd37;
    tile[365] = 6'd37;
    tile[366] = 6'd37;
    tile[367] = 6'd37;
    tile[368] = 6'd37;
    tile[369] = 6'd37;
    tile[370] = 6'd37;
    tile[371] = 6'd37;
    tile[372] = 6'd37;
    tile[373] = 6'd37;
    tile[374] = 6'd37;
    tile[375] = 6'd37;
    tile[376] = 6'd37;
    tile[377] = 6'd37;
    tile[378] = 6'd37;
    tile[379] = 6'd37;
    tile[380] = 6'd37;
    tile[381] = 6'd37;
    tile[382] = 6'd37;
    tile[383] = 6'd37;
    tile[384] = 6'd37;
    tile[385] = 6'd37;
    tile[386] = 6'd37;
    tile[387] = 6'd37;
    tile[388] = 6'd37;
    tile[389] = 6'd37;
    tile[390] = 6'd37;
    tile[391] = 6'd37;
    tile[392] = 6'd37;
    tile[393] = 6'd37;
    tile[394] = 6'd37;
    tile[395] = 6'd37;
    tile[396] = 6'd37;
    tile[397] = 6'd37;
    tile[398] = 6'd37;
    tile[399] = 6'd37;
    tile[400] = 6'd37;
    tile[401] = 6'd37;
    tile[402] = 6'd37;
    tile[403] = 6'd37;
    tile[404] = 6'd37;
    tile[405] = 6'd37;
    tile[406] = 6'd37;
    tile[407] = 6'd37;
    tile[408] = 6'd37;
    tile[409] = 6'd37;
    tile[410] = 6'd37;
    tile[411] = 6'd37;
    tile[412] = 6'd37;
    tile[413] = 6'd37;
    tile[414] = 6'd37;
    tile[415] = 6'd37;
    tile[416] = 6'd37;
    tile[417] = 6'd37;
    tile[418] = 6'd37;
    tile[419] = 6'd37;
    tile[420] = 6'd37;
    tile[421] = 6'd37;
    tile[422] = 6'd37;
    tile[423] = 6'd37;
    tile[424] = 6'd37;
    tile[425] = 6'd37;
    tile[426] = 6'd37;
    tile[427] = 6'd37;
    tile[428] = 6'd37;
    tile[429] = 6'd37;
    tile[430] = 6'd37;
    tile[431] = 6'd37;
    tile[432] = 6'd37;
    tile[433] = 6'd37;
    tile[434] = 6'd37;
    tile[435] = 6'd37;
    tile[436] = 6'd37;
    tile[437] = 6'd37;
    tile[438] = 6'd37;
    tile[439] = 6'd37;
    tile[440] = 6'd37;
    tile[441] = 6'd37;
    tile[442] = 6'd37;
    tile[443] = 6'd37;
    tile[444] = 6'd37;
    tile[445] = 6'd37;
    tile[446] = 6'd37;
    tile[447] = 6'd37;
    tile[448] = 6'd37;
    tile[449] = 6'd37;
    tile[450] = 6'd37;
    tile[451] = 6'd37;
    tile[452] = 6'd37;
    tile[453] = 6'd37;
    tile[454] = 6'd37;
    tile[455] = 6'd37;
    tile[456] = 6'd37;
    tile[457] = 6'd37;
    tile[458] = 6'd37;
    tile[459] = 6'd37;
    tile[460] = 6'd37;
    tile[461] = 6'd37;
    tile[462] = 6'd37;
    tile[463] = 6'd37;
    tile[464] = 6'd37;
    tile[465] = 6'd37;
    tile[466] = 6'd37;
    tile[467] = 6'd37;
    tile[468] = 6'd37;
    tile[469] = 6'd37;
    tile[470] = 6'd37;
    tile[471] = 6'd37;
    tile[472] = 6'd37;
    tile[473] = 6'd37;
    tile[474] = 6'd37;
    tile[475] = 6'd37;
    tile[476] = 6'd37;
    tile[477] = 6'd37;
    tile[478] = 6'd37;
    tile[479] = 6'd37;
    tile[480] = 6'd37;
    tile[481] = 6'd37;
    tile[482] = 6'd37;
    tile[483] = 6'd37;
    tile[484] = 6'd37;
    tile[485] = 6'd37;
    tile[486] = 6'd37;
    tile[487] = 6'd37;
    tile[488] = 6'd37;
    tile[489] = 6'd37;
    tile[490] = 6'd37;
    tile[491] = 6'd37;
    tile[492] = 6'd37;
    tile[493] = 6'd37;
    tile[494] = 6'd37;
    tile[495] = 6'd37;
    tile[496] = 6'd37;
    tile[497] = 6'd37;
    tile[498] = 6'd37;
    tile[499] = 6'd37;
    tile[500] = 6'd37;
    tile[501] = 6'd37;
    tile[502] = 6'd37;
    tile[503] = 6'd37;
    tile[504] = 6'd37;
    tile[505] = 6'd37;
    tile[506] = 6'd37;
    tile[507] = 6'd37;
    tile[508] = 6'd37;
    tile[509] = 6'd37;
    tile[510] = 6'd37;
    tile[511] = 6'd37;
    tile[512] = 6'd37;
    tile[513] = 6'd37;
    tile[514] = 6'd37;
    tile[515] = 6'd37;
    tile[516] = 6'd37;
    tile[517] = 6'd37;
    tile[518] = 6'd37;
    tile[519] = 6'd37;
    tile[520] = 6'd37;
    tile[521] = 6'd37;
    tile[522] = 6'd37;
    tile[523] = 6'd37;
    tile[524] = 6'd37;
    tile[525] = 6'd37;
    tile[526] = 6'd37;
    tile[527] = 6'd37;
    tile[528] = 6'd37;
    tile[529] = 6'd37;
    tile[530] = 6'd37;
    tile[531] = 6'd37;
    tile[532] = 6'd37;
    tile[533] = 6'd37;
    tile[534] = 6'd37;
    tile[535] = 6'd37;
    tile[536] = 6'd37;
    tile[537] = 6'd37;
    tile[538] = 6'd37;
    tile[539] = 6'd37;
    tile[540] = 6'd37;
    tile[541] = 6'd37;
    tile[542] = 6'd37;
    tile[543] = 6'd37;
    tile[544] = 6'd37;
    tile[545] = 6'd37;
    tile[546] = 6'd37;
    tile[547] = 6'd37;
    tile[548] = 6'd37;
    tile[549] = 6'd37;
    tile[550] = 6'd37;
    tile[551] = 6'd37;
    tile[552] = 6'd37;
    tile[553] = 6'd37;
    tile[554] = 6'd37;
    tile[555] = 6'd37;
    tile[556] = 6'd37;
    tile[557] = 6'd37;
    tile[558] = 6'd37;
    tile[559] = 6'd37;
    tile[560] = 6'd37;
    tile[561] = 6'd37;
    tile[562] = 6'd37;
    tile[563] = 6'd37;
    tile[564] = 6'd37;
    tile[565] = 6'd37;
    tile[566] = 6'd37;
    tile[567] = 6'd37;
    tile[568] = 6'd37;
    tile[569] = 6'd37;
    tile[570] = 6'd37;
    tile[571] = 6'd37;
    tile[572] = 6'd37;
    tile[573] = 6'd37;
    tile[574] = 6'd37;
    tile[575] = 6'd37;
    tile[576] = 6'd37;
    tile[577] = 6'd37;
    tile[578] = 6'd37;
    tile[579] = 6'd37;
    tile[580] = 6'd37;
    tile[581] = 6'd37;
    tile[582] = 6'd37;
    tile[583] = 6'd37;
    tile[584] = 6'd37;
    tile[585] = 6'd37;
    tile[586] = 6'd37;
    tile[587] = 6'd37;
    tile[588] = 6'd37;
    tile[589] = 6'd37;
    tile[590] = 6'd37;
    tile[591] = 6'd37;
    tile[592] = 6'd37;
    tile[593] = 6'd37;
    tile[594] = 6'd37;
    tile[595] = 6'd37;
    tile[596] = 6'd37;
    tile[597] = 6'd37;
    tile[598] = 6'd37;
    tile[599] = 6'd37;
    tile[600] = 6'd37;
    tile[601] = 6'd37;
    tile[602] = 6'd37;
    tile[603] = 6'd37;
    tile[604] = 6'd37;
    tile[605] = 6'd37;
    tile[606] = 6'd37;
    tile[607] = 6'd37;
    tile[608] = 6'd37;
    tile[609] = 6'd37;
    tile[610] = 6'd37;
    tile[611] = 6'd37;
    tile[612] = 6'd37;
    tile[613] = 6'd37;
    tile[614] = 6'd37;
    tile[615] = 6'd37;
    tile[616] = 6'd37;
    tile[617] = 6'd37;
    tile[618] = 6'd37;
    tile[619] = 6'd37;
    tile[620] = 6'd37;
    tile[621] = 6'd37;
    tile[622] = 6'd37;
    tile[623] = 6'd37;
    tile[624] = 6'd37;
    tile[625] = 6'd37;
    tile[626] = 6'd37;
    tile[627] = 6'd37;
    tile[628] = 6'd37;
    tile[629] = 6'd37;
    tile[630] = 6'd37;
    tile[631] = 6'd37;
    tile[632] = 6'd37;
    tile[633] = 6'd37;
    tile[634] = 6'd37;
    tile[635] = 6'd37;
    tile[636] = 6'd37;
    tile[637] = 6'd37;
    tile[638] = 6'd37;
    tile[639] = 6'd37;
    tile[640] = 6'd37;
    tile[641] = 6'd37;
    tile[642] = 6'd37;
    tile[643] = 6'd37;
    tile[644] = 6'd37;
    tile[645] = 6'd37;
    tile[646] = 6'd37;
    tile[647] = 6'd37;
    tile[648] = 6'd37;
    tile[649] = 6'd37;
    tile[650] = 6'd37;
    tile[651] = 6'd37;
    tile[652] = 6'd37;
    tile[653] = 6'd37;
    tile[654] = 6'd37;
    tile[655] = 6'd37;
    tile[656] = 6'd37;
    tile[657] = 6'd37;
    tile[658] = 6'd37;
    tile[659] = 6'd37;
    tile[660] = 6'd37;
    tile[661] = 6'd37;
    tile[662] = 6'd37;
    tile[663] = 6'd37;
    tile[664] = 6'd37;
    tile[665] = 6'd37;
    tile[666] = 6'd37;
    tile[667] = 6'd37;
    tile[668] = 6'd37;
    tile[669] = 6'd37;
    tile[670] = 6'd37;
    tile[671] = 6'd37;
    tile[672] = 6'd37;
    tile[673] = 6'd37;
    tile[674] = 6'd37;
    tile[675] = 6'd37;
    tile[676] = 6'd37;
    tile[677] = 6'd37;
    tile[678] = 6'd37;
    tile[679] = 6'd37;
    tile[680] = 6'd37;
    tile[681] = 6'd37;
    tile[682] = 6'd37;
    tile[683] = 6'd37;
    tile[684] = 6'd37;
    tile[685] = 6'd37;
    tile[686] = 6'd37;
    tile[687] = 6'd37;
    tile[688] = 6'd37;
    tile[689] = 6'd37;
    tile[690] = 6'd37;
    tile[691] = 6'd37;
    tile[692] = 6'd37;
    tile[693] = 6'd37;
    tile[694] = 6'd37;
    tile[695] = 6'd37;
    tile[696] = 6'd37;
    tile[697] = 6'd37;
    tile[698] = 6'd37;
    tile[699] = 6'd37;
    tile[700] = 6'd37;
    tile[701] = 6'd37;
    tile[702] = 6'd37;
    tile[703] = 6'd37;
    tile[704] = 6'd37;
    tile[705] = 6'd37;
    tile[706] = 6'd37;
    tile[707] = 6'd37;
    tile[708] = 6'd37;
    tile[709] = 6'd37;
    tile[710] = 6'd37;
    tile[711] = 6'd37;
    tile[712] = 6'd37;
    tile[713] = 6'd37;
    tile[714] = 6'd37;
    tile[715] = 6'd37;
    tile[716] = 6'd37;
    tile[717] = 6'd37;
    tile[718] = 6'd37;
    tile[719] = 6'd37;
    tile[720] = 6'd37;
    tile[721] = 6'd37;
    tile[722] = 6'd37;
    tile[723] = 6'd37;
    tile[724] = 6'd37;
    tile[725] = 6'd37;
    tile[726] = 6'd37;
    tile[727] = 6'd37;
    tile[728] = 6'd37;
    tile[729] = 6'd37;
    tile[730] = 6'd37;
    tile[731] = 6'd37;
    tile[732] = 6'd37;
    tile[733] = 6'd37;
    tile[734] = 6'd37;
    tile[735] = 6'd37;
    tile[736] = 6'd37;
    tile[737] = 6'd37;
    tile[738] = 6'd37;
    tile[739] = 6'd37;
    tile[740] = 6'd37;
    tile[741] = 6'd37;
    tile[742] = 6'd37;
    tile[743] = 6'd37;
    tile[744] = 6'd37;
    tile[745] = 6'd37;
    tile[746] = 6'd37;
    tile[747] = 6'd37;
    tile[748] = 6'd37;
    tile[749] = 6'd37;
    tile[750] = 6'd37;
    tile[751] = 6'd37;
    tile[752] = 6'd37;
    tile[753] = 6'd37;
    tile[754] = 6'd37;
    tile[755] = 6'd37;
    tile[756] = 6'd37;
    tile[757] = 6'd37;
    tile[758] = 6'd37;
    tile[759] = 6'd37;
    tile[760] = 6'd37;
    tile[761] = 6'd37;
    tile[762] = 6'd37;
    tile[763] = 6'd37;
    tile[764] = 6'd37;
    tile[765] = 6'd37;
    tile[766] = 6'd37;
    tile[767] = 6'd37;
    tile[768] = 6'd37;
    tile[769] = 6'd37;
    tile[770] = 6'd37;
    tile[771] = 6'd37;
    tile[772] = 6'd37;
    tile[773] = 6'd37;
    tile[774] = 6'd37;
    tile[775] = 6'd37;
    tile[776] = 6'd37;
    tile[777] = 6'd37;
    tile[778] = 6'd37;
    tile[779] = 6'd37;
    tile[780] = 6'd37;
    tile[781] = 6'd37;
    tile[782] = 6'd37;
    tile[783] = 6'd37;
    tile[784] = 6'd37;
    tile[785] = 6'd37;
    tile[786] = 6'd37;
    tile[787] = 6'd37;
    tile[788] = 6'd37;
    tile[789] = 6'd37;
    tile[790] = 6'd37;
    tile[791] = 6'd37;
    tile[792] = 6'd37;
    tile[793] = 6'd37;
    tile[794] = 6'd37;
    tile[795] = 6'd37;
    tile[796] = 6'd37;
    tile[797] = 6'd37;
    tile[798] = 6'd37;
    tile[799] = 6'd37;
    tile[800] = 6'd37;
    tile[801] = 6'd37;
    tile[802] = 6'd37;
    tile[803] = 6'd37;
    tile[804] = 6'd37;
    tile[805] = 6'd37;
    tile[806] = 6'd37;
    tile[807] = 6'd37;
    tile[808] = 6'd37;
    tile[809] = 6'd37;
    tile[810] = 6'd37;
    tile[811] = 6'd37;
    tile[812] = 6'd37;
    tile[813] = 6'd37;
    tile[814] = 6'd37;
    tile[815] = 6'd37;
    tile[816] = 6'd37;
    tile[817] = 6'd37;
    tile[818] = 6'd37;
    tile[819] = 6'd37;
    tile[820] = 6'd37;
    tile[821] = 6'd37;
    tile[822] = 6'd37;
    tile[823] = 6'd37;
    tile[824] = 6'd37;
    tile[825] = 6'd37;
    tile[826] = 6'd37;
    tile[827] = 6'd37;
    tile[828] = 6'd37;
    tile[829] = 6'd37;
    tile[830] = 6'd37;
    tile[831] = 6'd37;
    tile[832] = 6'd37;
    tile[833] = 6'd37;
    tile[834] = 6'd37;
    tile[835] = 6'd37;
    tile[836] = 6'd37;
    tile[837] = 6'd37;
    tile[838] = 6'd37;
    tile[839] = 6'd37;
    tile[840] = 6'd37;
    tile[841] = 6'd37;
    tile[842] = 6'd37;
    tile[843] = 6'd37;
    tile[844] = 6'd37;
    tile[845] = 6'd37;
    tile[846] = 6'd37;
    tile[847] = 6'd37;
    tile[848] = 6'd37;
    tile[849] = 6'd37;
    tile[850] = 6'd37;
    tile[851] = 6'd37;
    tile[852] = 6'd37;
    tile[853] = 6'd37;
    tile[854] = 6'd37;
    tile[855] = 6'd37;
    tile[856] = 6'd37;
    tile[857] = 6'd37;
    tile[858] = 6'd37;
    tile[859] = 6'd37;
    tile[860] = 6'd37;
    tile[861] = 6'd37;
    tile[862] = 6'd37;
    tile[863] = 6'd37;
    tile[864] = 6'd37;
    tile[865] = 6'd37;
    tile[866] = 6'd37;
    tile[867] = 6'd37;
    tile[868] = 6'd37;
    tile[869] = 6'd37;
    tile[870] = 6'd37;
    tile[871] = 6'd37;
    tile[872] = 6'd37;
    tile[873] = 6'd37;
    tile[874] = 6'd37;
    tile[875] = 6'd37;
    tile[876] = 6'd37;
    tile[877] = 6'd37;
    tile[878] = 6'd37;
    tile[879] = 6'd37;
    tile[880] = 6'd37;
    tile[881] = 6'd37;
    tile[882] = 6'd37;
    tile[883] = 6'd37;
    tile[884] = 6'd37;
    tile[885] = 6'd37;
    tile[886] = 6'd37;
    tile[887] = 6'd37;
    tile[888] = 6'd37;
    tile[889] = 6'd37;
    tile[890] = 6'd37;
    tile[891] = 6'd37;
    tile[892] = 6'd37;
    tile[893] = 6'd37;
    tile[894] = 6'd37;
    tile[895] = 6'd37;
    tile[896] = 6'd37;
    tile[897] = 6'd37;
    tile[898] = 6'd37;
    tile[899] = 6'd37;
    tile[900] = 6'd37;
    tile[901] = 6'd37;
    tile[902] = 6'd37;
    tile[903] = 6'd37;
    tile[904] = 6'd37;
    tile[905] = 6'd37;
    tile[906] = 6'd37;
    tile[907] = 6'd37;
    tile[908] = 6'd37;
    tile[909] = 6'd37;
    tile[910] = 6'd37;
    tile[911] = 6'd37;
    tile[912] = 6'd37;
    tile[913] = 6'd37;
    tile[914] = 6'd37;
    tile[915] = 6'd37;
    tile[916] = 6'd37;
    tile[917] = 6'd37;
    tile[918] = 6'd37;
    tile[919] = 6'd37;
    tile[920] = 6'd37;
    tile[921] = 6'd37;
    tile[922] = 6'd37;
    tile[923] = 6'd37;
    tile[924] = 6'd37;
    tile[925] = 6'd37;
    tile[926] = 6'd37;
    tile[927] = 6'd37;
    tile[928] = 6'd37;
    tile[929] = 6'd37;
    tile[930] = 6'd37;
    tile[931] = 6'd37;
    tile[932] = 6'd37;
    tile[933] = 6'd37;
    tile[934] = 6'd37;
    tile[935] = 6'd37;
    tile[936] = 6'd37;
    tile[937] = 6'd37;
    tile[938] = 6'd37;
    tile[939] = 6'd37;
    tile[940] = 6'd37;
    tile[941] = 6'd37;
    tile[942] = 6'd37;
    tile[943] = 6'd37;
    tile[944] = 6'd37;
    tile[945] = 6'd37;
    tile[946] = 6'd37;
    tile[947] = 6'd37;
    tile[948] = 6'd37;
    tile[949] = 6'd37;
    tile[950] = 6'd37;
    tile[951] = 6'd37;
    tile[952] = 6'd37;
    tile[953] = 6'd37;
    tile[954] = 6'd37;
    tile[955] = 6'd37;
    tile[956] = 6'd37;
    tile[957] = 6'd37;
    tile[958] = 6'd37;
    tile[959] = 6'd37;
    tile[960] = 6'd37;
    tile[961] = 6'd37;
    tile[962] = 6'd37;
    tile[963] = 6'd37;
    tile[964] = 6'd37;
    tile[965] = 6'd37;
    tile[966] = 6'd37;
    tile[967] = 6'd37;
    tile[968] = 6'd37;
    tile[969] = 6'd37;
    tile[970] = 6'd37;
    tile[971] = 6'd37;
    tile[972] = 6'd37;
    tile[973] = 6'd37;
    tile[974] = 6'd37;
    tile[975] = 6'd37;
    tile[976] = 6'd37;
    tile[977] = 6'd37;
    tile[978] = 6'd37;
    tile[979] = 6'd37;
    tile[980] = 6'd37;
    tile[981] = 6'd37;
    tile[982] = 6'd37;
    tile[983] = 6'd37;
    tile[984] = 6'd37;
    tile[985] = 6'd37;
    tile[986] = 6'd37;
    tile[987] = 6'd37;
    tile[988] = 6'd37;
    tile[989] = 6'd37;
    tile[990] = 6'd37;
    tile[991] = 6'd37;
    tile[992] = 6'd37;
    tile[993] = 6'd37;
    tile[994] = 6'd37;
    tile[995] = 6'd37;
    tile[996] = 6'd37;
    tile[997] = 6'd37;
    tile[998] = 6'd37;
    tile[999] = 6'd37;
    tile[1000] = 6'd37;
    tile[1001] = 6'd37;
    tile[1002] = 6'd37;
    tile[1003] = 6'd37;
    tile[1004] = 6'd37;
    tile[1005] = 6'd37;
    tile[1006] = 6'd37;
    tile[1007] = 6'd37;
    tile[1008] = 6'd37;
    tile[1009] = 6'd37;
    tile[1010] = 6'd37;
    tile[1011] = 6'd37;
    tile[1012] = 6'd37;
    tile[1013] = 6'd37;
    tile[1014] = 6'd37;
    tile[1015] = 6'd37;
    tile[1016] = 6'd37;
    tile[1017] = 6'd37;
    tile[1018] = 6'd37;
    tile[1019] = 6'd37;
    tile[1020] = 6'd37;
    tile[1021] = 6'd37;
    tile[1022] = 6'd37;
    tile[1023] = 6'd37;
    tile[1024] = 6'd37;
    tile[1025] = 6'd37;
    tile[1026] = 6'd37;
    tile[1027] = 6'd37;
    tile[1028] = 6'd37;
    tile[1029] = 6'd37;
    tile[1030] = 6'd37;
    tile[1031] = 6'd37;
    tile[1032] = 6'd37;
    tile[1033] = 6'd37;
    tile[1034] = 6'd37;
    tile[1035] = 6'd37;
    tile[1036] = 6'd37;
    tile[1037] = 6'd37;
    tile[1038] = 6'd37;
    tile[1039] = 6'd37;
    tile[1040] = 6'd37;
    tile[1041] = 6'd37;
    tile[1042] = 6'd37;
    tile[1043] = 6'd37;
    tile[1044] = 6'd37;
    tile[1045] = 6'd37;
    tile[1046] = 6'd37;
    tile[1047] = 6'd37;
    tile[1048] = 6'd37;
    tile[1049] = 6'd37;
    tile[1050] = 6'd37;
    tile[1051] = 6'd37;
    tile[1052] = 6'd37;
    tile[1053] = 6'd37;
    tile[1054] = 6'd37;
    tile[1055] = 6'd37;
    tile[1056] = 6'd37;
    tile[1057] = 6'd37;
    tile[1058] = 6'd37;
    tile[1059] = 6'd37;
    tile[1060] = 6'd37;
    tile[1061] = 6'd37;
    tile[1062] = 6'd37;
    tile[1063] = 6'd37;
    tile[1064] = 6'd37;
    tile[1065] = 6'd37;
    tile[1066] = 6'd37;
    tile[1067] = 6'd37;
    tile[1068] = 6'd37;
    tile[1069] = 6'd37;
    tile[1070] = 6'd37;
    tile[1071] = 6'd37;
    tile[1072] = 6'd37;
    tile[1073] = 6'd37;
    tile[1074] = 6'd37;
    tile[1075] = 6'd37;
    tile[1076] = 6'd37;
    tile[1077] = 6'd37;
    tile[1078] = 6'd37;
    tile[1079] = 6'd37;
    tile[1080] = 6'd37;
    tile[1081] = 6'd37;
    tile[1082] = 6'd37;
    tile[1083] = 6'd37;
    tile[1084] = 6'd37;
    tile[1085] = 6'd37;
    tile[1086] = 6'd37;
    tile[1087] = 6'd37;
    tile[1088] = 6'd37;
    tile[1089] = 6'd37;
    tile[1090] = 6'd37;
    tile[1091] = 6'd37;
    tile[1092] = 6'd37;
    tile[1093] = 6'd37;
    tile[1094] = 6'd37;
    tile[1095] = 6'd37;
    tile[1096] = 6'd37;
    tile[1097] = 6'd37;
    tile[1098] = 6'd37;
    tile[1099] = 6'd37;
    tile[1100] = 6'd37;
    tile[1101] = 6'd37;
    tile[1102] = 6'd37;
    tile[1103] = 6'd37;
    tile[1104] = 6'd37;
    tile[1105] = 6'd37;
    tile[1106] = 6'd37;
    tile[1107] = 6'd37;
    tile[1108] = 6'd37;
    tile[1109] = 6'd37;
    tile[1110] = 6'd37;
    tile[1111] = 6'd37;
    tile[1112] = 6'd37;
    tile[1113] = 6'd37;
    tile[1114] = 6'd37;
    tile[1115] = 6'd37;
    tile[1116] = 6'd37;
    tile[1117] = 6'd37;
    tile[1118] = 6'd37;
    tile[1119] = 6'd37;
    tile[1120] = 6'd37;
    tile[1121] = 6'd37;
    tile[1122] = 6'd37;
    tile[1123] = 6'd37;
    tile[1124] = 6'd37;
    tile[1125] = 6'd37;
    tile[1126] = 6'd37;
    tile[1127] = 6'd37;
    tile[1128] = 6'd37;
    tile[1129] = 6'd37;
    tile[1130] = 6'd37;
    tile[1131] = 6'd37;
    tile[1132] = 6'd37;
    tile[1133] = 6'd37;
    tile[1134] = 6'd37;
    tile[1135] = 6'd37;
    tile[1136] = 6'd37;
    tile[1137] = 6'd37;
    tile[1138] = 6'd37;
    tile[1139] = 6'd37;
    tile[1140] = 6'd37;
    tile[1141] = 6'd37;
    tile[1142] = 6'd37;
    tile[1143] = 6'd37;
    tile[1144] = 6'd37;
    tile[1145] = 6'd37;
    tile[1146] = 6'd37;
    tile[1147] = 6'd37;
    tile[1148] = 6'd37;
    tile[1149] = 6'd37;
    tile[1150] = 6'd37;
    tile[1151] = 6'd37;
    tile[1152] = 6'd37;
    tile[1153] = 6'd37;
    tile[1154] = 6'd37;
    tile[1155] = 6'd37;
    tile[1156] = 6'd37;
    tile[1157] = 6'd37;
    tile[1158] = 6'd37;
    tile[1159] = 6'd37;
    tile[1160] = 6'd37;
    tile[1161] = 6'd37;
    tile[1162] = 6'd37;
    tile[1163] = 6'd37;
    tile[1164] = 6'd37;
    tile[1165] = 6'd37;
    tile[1166] = 6'd37;
    tile[1167] = 6'd37;
    tile[1168] = 6'd37;
    tile[1169] = 6'd37;
    tile[1170] = 6'd37;
    tile[1171] = 6'd37;
    tile[1172] = 6'd37;
    tile[1173] = 6'd37;
    tile[1174] = 6'd37;
    tile[1175] = 6'd37;
    tile[1176] = 6'd37;
    tile[1177] = 6'd37;
    tile[1178] = 6'd37;
    tile[1179] = 6'd37;
    tile[1180] = 6'd37;
    tile[1181] = 6'd37;
    tile[1182] = 6'd37;
    tile[1183] = 6'd37;
    tile[1184] = 6'd37;
    tile[1185] = 6'd37;
    tile[1186] = 6'd37;
    tile[1187] = 6'd37;
    tile[1188] = 6'd37;
    tile[1189] = 6'd37;
    tile[1190] = 6'd37;
    tile[1191] = 6'd37;
    tile[1192] = 6'd37;
    tile[1193] = 6'd37;
    tile[1194] = 6'd37;
    tile[1195] = 6'd37;
    tile[1196] = 6'd37;
    tile[1197] = 6'd37;
    tile[1198] = 6'd37;
    tile[1199] = 6'd37;
    tile[1200] = 6'd37;
    tile[1201] = 6'd37;
    tile[1202] = 6'd37;
    tile[1203] = 6'd37;
    tile[1204] = 6'd37;
    tile[1205] = 6'd37;
    tile[1206] = 6'd37;
    tile[1207] = 6'd37;
    tile[1208] = 6'd37;
    tile[1209] = 6'd37;
    tile[1210] = 6'd37;
    tile[1211] = 6'd37;
    tile[1212] = 6'd37;
    tile[1213] = 6'd37;
    tile[1214] = 6'd37;
    tile[1215] = 6'd37;
    tile[1216] = 6'd37;
    tile[1217] = 6'd37;
    tile[1218] = 6'd37;
    tile[1219] = 6'd37;
    tile[1220] = 6'd37;
    tile[1221] = 6'd37;
    tile[1222] = 6'd37;
    tile[1223] = 6'd37;
    tile[1224] = 6'd37;
    tile[1225] = 6'd37;
    tile[1226] = 6'd0;
    tile[1227] = 6'd1;
    tile[1228] = 6'd1;
    tile[1229] = 6'd1;
    tile[1230] = 6'd1;
    tile[1231] = 6'd1;
    tile[1232] = 6'd1;
    tile[1233] = 6'd1;
    tile[1234] = 6'd1;
    tile[1235] = 6'd1;
    tile[1236] = 6'd1;
    tile[1237] = 6'd1;
    tile[1238] = 6'd1;
    tile[1239] = 6'd2;
    tile[1240] = 6'd3;
    tile[1241] = 6'd1;
    tile[1242] = 6'd1;
    tile[1243] = 6'd1;
    tile[1244] = 6'd1;
    tile[1245] = 6'd1;
    tile[1246] = 6'd1;
    tile[1247] = 6'd1;
    tile[1248] = 6'd1;
    tile[1249] = 6'd1;
    tile[1250] = 6'd1;
    tile[1251] = 6'd1;
    tile[1252] = 6'd1;
    tile[1253] = 6'd4;
    tile[1254] = 6'd37;
    tile[1255] = 6'd37;
    tile[1256] = 6'd37;
    tile[1257] = 6'd37;
    tile[1258] = 6'd37;
    tile[1259] = 6'd37;
    tile[1260] = 6'd37;
    tile[1261] = 6'd37;
    tile[1262] = 6'd37;
    tile[1263] = 6'd37;
    tile[1264] = 6'd37;
    tile[1265] = 6'd37;
    tile[1266] = 6'd37;
    tile[1267] = 6'd37;
    tile[1268] = 6'd37;
    tile[1269] = 6'd37;
    tile[1270] = 6'd37;
    tile[1271] = 6'd37;
    tile[1272] = 6'd37;
    tile[1273] = 6'd37;
    tile[1274] = 6'd37;
    tile[1275] = 6'd37;
    tile[1276] = 6'd37;
    tile[1277] = 6'd37;
    tile[1278] = 6'd37;
    tile[1279] = 6'd37;
    tile[1280] = 6'd37;
    tile[1281] = 6'd37;
    tile[1282] = 6'd37;
    tile[1283] = 6'd37;
    tile[1284] = 6'd37;
    tile[1285] = 6'd37;
    tile[1286] = 6'd37;
    tile[1287] = 6'd37;
    tile[1288] = 6'd37;
    tile[1289] = 6'd37;
    tile[1290] = 6'd37;
    tile[1291] = 6'd37;
    tile[1292] = 6'd37;
    tile[1293] = 6'd37;
    tile[1294] = 6'd37;
    tile[1295] = 6'd37;
    tile[1296] = 6'd37;
    tile[1297] = 6'd37;
    tile[1298] = 6'd37;
    tile[1299] = 6'd37;
    tile[1300] = 6'd37;
    tile[1301] = 6'd37;
    tile[1302] = 6'd37;
    tile[1303] = 6'd37;
    tile[1304] = 6'd37;
    tile[1305] = 6'd37;
    tile[1306] = 6'd9;
    tile[1307] = 6'd10;
    tile[1308] = 6'd10;
    tile[1309] = 6'd10;
    tile[1310] = 6'd10;
    tile[1311] = 6'd10;
    tile[1312] = 6'd10;
    tile[1313] = 6'd10;
    tile[1314] = 6'd10;
    tile[1315] = 6'd10;
    tile[1316] = 6'd10;
    tile[1317] = 6'd10;
    tile[1318] = 6'd10;
    tile[1319] = 6'd11;
    tile[1320] = 6'd12;
    tile[1321] = 6'd10;
    tile[1322] = 6'd10;
    tile[1323] = 6'd10;
    tile[1324] = 6'd10;
    tile[1325] = 6'd10;
    tile[1326] = 6'd10;
    tile[1327] = 6'd10;
    tile[1328] = 6'd10;
    tile[1329] = 6'd10;
    tile[1330] = 6'd10;
    tile[1331] = 6'd10;
    tile[1332] = 6'd10;
    tile[1333] = 6'd13;
    tile[1334] = 6'd37;
    tile[1335] = 6'd37;
    tile[1336] = 6'd37;
    tile[1337] = 6'd37;
    tile[1338] = 6'd37;
    tile[1339] = 6'd37;
    tile[1340] = 6'd37;
    tile[1341] = 6'd37;
    tile[1342] = 6'd37;
    tile[1343] = 6'd37;
    tile[1344] = 6'd37;
    tile[1345] = 6'd37;
    tile[1346] = 6'd37;
    tile[1347] = 6'd37;
    tile[1348] = 6'd37;
    tile[1349] = 6'd37;
    tile[1350] = 6'd37;
    tile[1351] = 6'd37;
    tile[1352] = 6'd37;
    tile[1353] = 6'd37;
    tile[1354] = 6'd37;
    tile[1355] = 6'd37;
    tile[1356] = 6'd37;
    tile[1357] = 6'd37;
    tile[1358] = 6'd37;
    tile[1359] = 6'd37;
    tile[1360] = 6'd37;
    tile[1361] = 6'd37;
    tile[1362] = 6'd37;
    tile[1363] = 6'd37;
    tile[1364] = 6'd37;
    tile[1365] = 6'd37;
    tile[1366] = 6'd37;
    tile[1367] = 6'd37;
    tile[1368] = 6'd37;
    tile[1369] = 6'd37;
    tile[1370] = 6'd37;
    tile[1371] = 6'd37;
    tile[1372] = 6'd37;
    tile[1373] = 6'd37;
    tile[1374] = 6'd37;
    tile[1375] = 6'd37;
    tile[1376] = 6'd37;
    tile[1377] = 6'd37;
    tile[1378] = 6'd37;
    tile[1379] = 6'd37;
    tile[1380] = 6'd37;
    tile[1381] = 6'd37;
    tile[1382] = 6'd37;
    tile[1383] = 6'd37;
    tile[1384] = 6'd37;
    tile[1385] = 6'd37;
    tile[1386] = 6'd9;
    tile[1387] = 6'd10;
    tile[1388] = 6'd7;
    tile[1389] = 6'd16;
    tile[1390] = 6'd16;
    tile[1391] = 6'd8;
    tile[1392] = 6'd10;
    tile[1393] = 6'd7;
    tile[1394] = 6'd16;
    tile[1395] = 6'd16;
    tile[1396] = 6'd16;
    tile[1397] = 6'd8;
    tile[1398] = 6'd10;
    tile[1399] = 6'd11;
    tile[1400] = 6'd12;
    tile[1401] = 6'd10;
    tile[1402] = 6'd7;
    tile[1403] = 6'd16;
    tile[1404] = 6'd16;
    tile[1405] = 6'd16;
    tile[1406] = 6'd8;
    tile[1407] = 6'd10;
    tile[1408] = 6'd7;
    tile[1409] = 6'd16;
    tile[1410] = 6'd16;
    tile[1411] = 6'd8;
    tile[1412] = 6'd10;
    tile[1413] = 6'd13;
    tile[1414] = 6'd37;
    tile[1415] = 6'd37;
    tile[1416] = 6'd37;
    tile[1417] = 6'd37;
    tile[1418] = 6'd37;
    tile[1419] = 6'd37;
    tile[1420] = 6'd37;
    tile[1421] = 6'd37;
    tile[1422] = 6'd37;
    tile[1423] = 6'd37;
    tile[1424] = 6'd37;
    tile[1425] = 6'd37;
    tile[1426] = 6'd37;
    tile[1427] = 6'd37;
    tile[1428] = 6'd37;
    tile[1429] = 6'd37;
    tile[1430] = 6'd37;
    tile[1431] = 6'd37;
    tile[1432] = 6'd37;
    tile[1433] = 6'd37;
    tile[1434] = 6'd37;
    tile[1435] = 6'd37;
    tile[1436] = 6'd37;
    tile[1437] = 6'd37;
    tile[1438] = 6'd37;
    tile[1439] = 6'd37;
    tile[1440] = 6'd37;
    tile[1441] = 6'd37;
    tile[1442] = 6'd37;
    tile[1443] = 6'd37;
    tile[1444] = 6'd37;
    tile[1445] = 6'd37;
    tile[1446] = 6'd37;
    tile[1447] = 6'd37;
    tile[1448] = 6'd37;
    tile[1449] = 6'd37;
    tile[1450] = 6'd37;
    tile[1451] = 6'd37;
    tile[1452] = 6'd37;
    tile[1453] = 6'd37;
    tile[1454] = 6'd37;
    tile[1455] = 6'd37;
    tile[1456] = 6'd37;
    tile[1457] = 6'd37;
    tile[1458] = 6'd37;
    tile[1459] = 6'd37;
    tile[1460] = 6'd37;
    tile[1461] = 6'd37;
    tile[1462] = 6'd37;
    tile[1463] = 6'd37;
    tile[1464] = 6'd37;
    tile[1465] = 6'd37;
    tile[1466] = 6'd9;
    tile[1467] = 6'd20;
    tile[1468] = 6'd12;
    tile[1469] = 6'd37;
    tile[1470] = 6'd37;
    tile[1471] = 6'd11;
    tile[1472] = 6'd10;
    tile[1473] = 6'd12;
    tile[1474] = 6'd37;
    tile[1475] = 6'd37;
    tile[1476] = 6'd37;
    tile[1477] = 6'd11;
    tile[1478] = 6'd10;
    tile[1479] = 6'd11;
    tile[1480] = 6'd13;
    tile[1481] = 6'd10;
    tile[1482] = 6'd12;
    tile[1483] = 6'd37;
    tile[1484] = 6'd37;
    tile[1485] = 6'd37;
    tile[1486] = 6'd11;
    tile[1487] = 6'd10;
    tile[1488] = 6'd12;
    tile[1489] = 6'd37;
    tile[1490] = 6'd37;
    tile[1491] = 6'd11;
    tile[1492] = 6'd10;
    tile[1493] = 6'd13;
    tile[1494] = 6'd37;
    tile[1495] = 6'd37;
    tile[1496] = 6'd37;
    tile[1497] = 6'd37;
    tile[1498] = 6'd37;
    tile[1499] = 6'd37;
    tile[1500] = 6'd37;
    tile[1501] = 6'd37;
    tile[1502] = 6'd37;
    tile[1503] = 6'd37;
    tile[1504] = 6'd37;
    tile[1505] = 6'd37;
    tile[1506] = 6'd37;
    tile[1507] = 6'd37;
    tile[1508] = 6'd37;
    tile[1509] = 6'd37;
    tile[1510] = 6'd37;
    tile[1511] = 6'd37;
    tile[1512] = 6'd37;
    tile[1513] = 6'd37;
    tile[1514] = 6'd37;
    tile[1515] = 6'd37;
    tile[1516] = 6'd37;
    tile[1517] = 6'd37;
    tile[1518] = 6'd37;
    tile[1519] = 6'd37;
    tile[1520] = 6'd37;
    tile[1521] = 6'd37;
    tile[1522] = 6'd37;
    tile[1523] = 6'd37;
    tile[1524] = 6'd37;
    tile[1525] = 6'd37;
    tile[1526] = 6'd37;
    tile[1527] = 6'd37;
    tile[1528] = 6'd37;
    tile[1529] = 6'd37;
    tile[1530] = 6'd37;
    tile[1531] = 6'd37;
    tile[1532] = 6'd37;
    tile[1533] = 6'd37;
    tile[1534] = 6'd37;
    tile[1535] = 6'd37;
    tile[1536] = 6'd37;
    tile[1537] = 6'd37;
    tile[1538] = 6'd37;
    tile[1539] = 6'd37;
    tile[1540] = 6'd37;
    tile[1541] = 6'd37;
    tile[1542] = 6'd37;
    tile[1543] = 6'd37;
    tile[1544] = 6'd37;
    tile[1545] = 6'd37;
    tile[1546] = 6'd9;
    tile[1547] = 6'd10;
    tile[1548] = 6'd17;
    tile[1549] = 6'd6;
    tile[1550] = 6'd6;
    tile[1551] = 6'd18;
    tile[1552] = 6'd10;
    tile[1553] = 6'd17;
    tile[1554] = 6'd6;
    tile[1555] = 6'd6;
    tile[1556] = 6'd6;
    tile[1557] = 6'd18;
    tile[1558] = 6'd10;
    tile[1559] = 6'd21;
    tile[1560] = 6'd22;
    tile[1561] = 6'd10;
    tile[1562] = 6'd17;
    tile[1563] = 6'd6;
    tile[1564] = 6'd6;
    tile[1565] = 6'd6;
    tile[1566] = 6'd18;
    tile[1567] = 6'd10;
    tile[1568] = 6'd17;
    tile[1569] = 6'd6;
    tile[1570] = 6'd6;
    tile[1571] = 6'd18;
    tile[1572] = 6'd10;
    tile[1573] = 6'd13;
    tile[1574] = 6'd37;
    tile[1575] = 6'd37;
    tile[1576] = 6'd37;
    tile[1577] = 6'd37;
    tile[1578] = 6'd37;
    tile[1579] = 6'd37;
    tile[1580] = 6'd37;
    tile[1581] = 6'd37;
    tile[1582] = 6'd37;
    tile[1583] = 6'd37;
    tile[1584] = 6'd37;
    tile[1585] = 6'd37;
    tile[1586] = 6'd37;
    tile[1587] = 6'd37;
    tile[1588] = 6'd37;
    tile[1589] = 6'd37;
    tile[1590] = 6'd37;
    tile[1591] = 6'd37;
    tile[1592] = 6'd37;
    tile[1593] = 6'd37;
    tile[1594] = 6'd37;
    tile[1595] = 6'd37;
    tile[1596] = 6'd37;
    tile[1597] = 6'd37;
    tile[1598] = 6'd37;
    tile[1599] = 6'd37;
    tile[1600] = 6'd37;
    tile[1601] = 6'd37;
    tile[1602] = 6'd37;
    tile[1603] = 6'd37;
    tile[1604] = 6'd37;
    tile[1605] = 6'd37;
    tile[1606] = 6'd37;
    tile[1607] = 6'd37;
    tile[1608] = 6'd37;
    tile[1609] = 6'd37;
    tile[1610] = 6'd37;
    tile[1611] = 6'd37;
    tile[1612] = 6'd37;
    tile[1613] = 6'd37;
    tile[1614] = 6'd37;
    tile[1615] = 6'd37;
    tile[1616] = 6'd37;
    tile[1617] = 6'd37;
    tile[1618] = 6'd37;
    tile[1619] = 6'd37;
    tile[1620] = 6'd37;
    tile[1621] = 6'd37;
    tile[1622] = 6'd37;
    tile[1623] = 6'd37;
    tile[1624] = 6'd37;
    tile[1625] = 6'd37;
    tile[1626] = 6'd9;
    tile[1627] = 6'd10;
    tile[1628] = 6'd10;
    tile[1629] = 6'd10;
    tile[1630] = 6'd10;
    tile[1631] = 6'd10;
    tile[1632] = 6'd10;
    tile[1633] = 6'd10;
    tile[1634] = 6'd10;
    tile[1635] = 6'd10;
    tile[1636] = 6'd10;
    tile[1637] = 6'd10;
    tile[1638] = 6'd10;
    tile[1639] = 6'd10;
    tile[1640] = 6'd10;
    tile[1641] = 6'd10;
    tile[1642] = 6'd10;
    tile[1643] = 6'd10;
    tile[1644] = 6'd10;
    tile[1645] = 6'd10;
    tile[1646] = 6'd10;
    tile[1647] = 6'd10;
    tile[1648] = 6'd10;
    tile[1649] = 6'd10;
    tile[1650] = 6'd10;
    tile[1651] = 6'd10;
    tile[1652] = 6'd10;
    tile[1653] = 6'd13;
    tile[1654] = 6'd37;
    tile[1655] = 6'd37;
    tile[1656] = 6'd37;
    tile[1657] = 6'd37;
    tile[1658] = 6'd37;
    tile[1659] = 6'd37;
    tile[1660] = 6'd37;
    tile[1661] = 6'd37;
    tile[1662] = 6'd37;
    tile[1663] = 6'd37;
    tile[1664] = 6'd37;
    tile[1665] = 6'd37;
    tile[1666] = 6'd37;
    tile[1667] = 6'd37;
    tile[1668] = 6'd37;
    tile[1669] = 6'd37;
    tile[1670] = 6'd37;
    tile[1671] = 6'd37;
    tile[1672] = 6'd37;
    tile[1673] = 6'd37;
    tile[1674] = 6'd37;
    tile[1675] = 6'd37;
    tile[1676] = 6'd37;
    tile[1677] = 6'd37;
    tile[1678] = 6'd37;
    tile[1679] = 6'd37;
    tile[1680] = 6'd37;
    tile[1681] = 6'd37;
    tile[1682] = 6'd37;
    tile[1683] = 6'd37;
    tile[1684] = 6'd37;
    tile[1685] = 6'd37;
    tile[1686] = 6'd37;
    tile[1687] = 6'd37;
    tile[1688] = 6'd37;
    tile[1689] = 6'd37;
    tile[1690] = 6'd37;
    tile[1691] = 6'd37;
    tile[1692] = 6'd37;
    tile[1693] = 6'd37;
    tile[1694] = 6'd37;
    tile[1695] = 6'd37;
    tile[1696] = 6'd37;
    tile[1697] = 6'd37;
    tile[1698] = 6'd37;
    tile[1699] = 6'd37;
    tile[1700] = 6'd37;
    tile[1701] = 6'd37;
    tile[1702] = 6'd37;
    tile[1703] = 6'd37;
    tile[1704] = 6'd37;
    tile[1705] = 6'd37;
    tile[1706] = 6'd9;
    tile[1707] = 6'd10;
    tile[1708] = 6'd7;
    tile[1709] = 6'd16;
    tile[1710] = 6'd16;
    tile[1711] = 6'd8;
    tile[1712] = 6'd10;
    tile[1713] = 6'd7;
    tile[1714] = 6'd8;
    tile[1715] = 6'd10;
    tile[1716] = 6'd7;
    tile[1717] = 6'd16;
    tile[1718] = 6'd16;
    tile[1719] = 6'd16;
    tile[1720] = 6'd16;
    tile[1721] = 6'd16;
    tile[1722] = 6'd16;
    tile[1723] = 6'd8;
    tile[1724] = 6'd10;
    tile[1725] = 6'd7;
    tile[1726] = 6'd8;
    tile[1727] = 6'd10;
    tile[1728] = 6'd7;
    tile[1729] = 6'd16;
    tile[1730] = 6'd16;
    tile[1731] = 6'd8;
    tile[1732] = 6'd10;
    tile[1733] = 6'd13;
    tile[1734] = 6'd37;
    tile[1735] = 6'd37;
    tile[1736] = 6'd37;
    tile[1737] = 6'd37;
    tile[1738] = 6'd37;
    tile[1739] = 6'd37;
    tile[1740] = 6'd37;
    tile[1741] = 6'd37;
    tile[1742] = 6'd37;
    tile[1743] = 6'd37;
    tile[1744] = 6'd37;
    tile[1745] = 6'd37;
    tile[1746] = 6'd37;
    tile[1747] = 6'd37;
    tile[1748] = 6'd37;
    tile[1749] = 6'd37;
    tile[1750] = 6'd37;
    tile[1751] = 6'd37;
    tile[1752] = 6'd37;
    tile[1753] = 6'd37;
    tile[1754] = 6'd37;
    tile[1755] = 6'd37;
    tile[1756] = 6'd37;
    tile[1757] = 6'd37;
    tile[1758] = 6'd37;
    tile[1759] = 6'd37;
    tile[1760] = 6'd37;
    tile[1761] = 6'd37;
    tile[1762] = 6'd37;
    tile[1763] = 6'd37;
    tile[1764] = 6'd37;
    tile[1765] = 6'd37;
    tile[1766] = 6'd37;
    tile[1767] = 6'd37;
    tile[1768] = 6'd37;
    tile[1769] = 6'd37;
    tile[1770] = 6'd37;
    tile[1771] = 6'd37;
    tile[1772] = 6'd37;
    tile[1773] = 6'd37;
    tile[1774] = 6'd37;
    tile[1775] = 6'd37;
    tile[1776] = 6'd37;
    tile[1777] = 6'd37;
    tile[1778] = 6'd37;
    tile[1779] = 6'd37;
    tile[1780] = 6'd37;
    tile[1781] = 6'd37;
    tile[1782] = 6'd37;
    tile[1783] = 6'd37;
    tile[1784] = 6'd37;
    tile[1785] = 6'd37;
    tile[1786] = 6'd9;
    tile[1787] = 6'd10;
    tile[1788] = 6'd17;
    tile[1789] = 6'd6;
    tile[1790] = 6'd6;
    tile[1791] = 6'd18;
    tile[1792] = 6'd10;
    tile[1793] = 6'd12;
    tile[1794] = 6'd11;
    tile[1795] = 6'd10;
    tile[1796] = 6'd7;
    tile[1797] = 6'd6;
    tile[1798] = 6'd6;
    tile[1799] = 6'd29;
    tile[1800] = 6'd27;
    tile[1801] = 6'd1;
    tile[1802] = 6'd2;
    tile[1803] = 6'd18;
    tile[1804] = 6'd10;
    tile[1805] = 6'd12;
    tile[1806] = 6'd11;
    tile[1807] = 6'd10;
    tile[1808] = 6'd17;
    tile[1809] = 6'd6;
    tile[1810] = 6'd6;
    tile[1811] = 6'd18;
    tile[1812] = 6'd10;
    tile[1813] = 6'd13;
    tile[1814] = 6'd37;
    tile[1815] = 6'd37;
    tile[1816] = 6'd37;
    tile[1817] = 6'd37;
    tile[1818] = 6'd37;
    tile[1819] = 6'd37;
    tile[1820] = 6'd37;
    tile[1821] = 6'd37;
    tile[1822] = 6'd37;
    tile[1823] = 6'd37;
    tile[1824] = 6'd37;
    tile[1825] = 6'd37;
    tile[1826] = 6'd37;
    tile[1827] = 6'd37;
    tile[1828] = 6'd37;
    tile[1829] = 6'd37;
    tile[1830] = 6'd37;
    tile[1831] = 6'd37;
    tile[1832] = 6'd37;
    tile[1833] = 6'd37;
    tile[1834] = 6'd37;
    tile[1835] = 6'd37;
    tile[1836] = 6'd37;
    tile[1837] = 6'd37;
    tile[1838] = 6'd37;
    tile[1839] = 6'd37;
    tile[1840] = 6'd37;
    tile[1841] = 6'd37;
    tile[1842] = 6'd37;
    tile[1843] = 6'd37;
    tile[1844] = 6'd37;
    tile[1845] = 6'd37;
    tile[1846] = 6'd37;
    tile[1847] = 6'd37;
    tile[1848] = 6'd37;
    tile[1849] = 6'd37;
    tile[1850] = 6'd37;
    tile[1851] = 6'd37;
    tile[1852] = 6'd37;
    tile[1853] = 6'd37;
    tile[1854] = 6'd37;
    tile[1855] = 6'd37;
    tile[1856] = 6'd37;
    tile[1857] = 6'd37;
    tile[1858] = 6'd37;
    tile[1859] = 6'd37;
    tile[1860] = 6'd37;
    tile[1861] = 6'd37;
    tile[1862] = 6'd37;
    tile[1863] = 6'd37;
    tile[1864] = 6'd37;
    tile[1865] = 6'd37;
    tile[1866] = 6'd9;
    tile[1867] = 6'd10;
    tile[1868] = 6'd10;
    tile[1869] = 6'd10;
    tile[1870] = 6'd10;
    tile[1871] = 6'd10;
    tile[1872] = 6'd10;
    tile[1873] = 6'd12;
    tile[1874] = 6'd11;
    tile[1875] = 6'd10;
    tile[1876] = 6'd10;
    tile[1877] = 6'd10;
    tile[1878] = 6'd10;
    tile[1879] = 6'd12;
    tile[1880] = 6'd11;
    tile[1881] = 6'd10;
    tile[1882] = 6'd10;
    tile[1883] = 6'd10;
    tile[1884] = 6'd10;
    tile[1885] = 6'd12;
    tile[1886] = 6'd11;
    tile[1887] = 6'd10;
    tile[1888] = 6'd10;
    tile[1889] = 6'd10;
    tile[1890] = 6'd10;
    tile[1891] = 6'd10;
    tile[1892] = 6'd10;
    tile[1893] = 6'd13;
    tile[1894] = 6'd37;
    tile[1895] = 6'd37;
    tile[1896] = 6'd37;
    tile[1897] = 6'd37;
    tile[1898] = 6'd37;
    tile[1899] = 6'd37;
    tile[1900] = 6'd37;
    tile[1901] = 6'd37;
    tile[1902] = 6'd37;
    tile[1903] = 6'd37;
    tile[1904] = 6'd37;
    tile[1905] = 6'd37;
    tile[1906] = 6'd37;
    tile[1907] = 6'd37;
    tile[1908] = 6'd37;
    tile[1909] = 6'd37;
    tile[1910] = 6'd37;
    tile[1911] = 6'd37;
    tile[1912] = 6'd37;
    tile[1913] = 6'd37;
    tile[1914] = 6'd37;
    tile[1915] = 6'd37;
    tile[1916] = 6'd37;
    tile[1917] = 6'd37;
    tile[1918] = 6'd37;
    tile[1919] = 6'd37;
    tile[1920] = 6'd37;
    tile[1921] = 6'd37;
    tile[1922] = 6'd37;
    tile[1923] = 6'd37;
    tile[1924] = 6'd37;
    tile[1925] = 6'd37;
    tile[1926] = 6'd37;
    tile[1927] = 6'd37;
    tile[1928] = 6'd37;
    tile[1929] = 6'd37;
    tile[1930] = 6'd37;
    tile[1931] = 6'd37;
    tile[1932] = 6'd37;
    tile[1933] = 6'd37;
    tile[1934] = 6'd37;
    tile[1935] = 6'd37;
    tile[1936] = 6'd37;
    tile[1937] = 6'd37;
    tile[1938] = 6'd37;
    tile[1939] = 6'd37;
    tile[1940] = 6'd37;
    tile[1941] = 6'd37;
    tile[1942] = 6'd37;
    tile[1943] = 6'd37;
    tile[1944] = 6'd37;
    tile[1945] = 6'd37;
    tile[1946] = 6'd19;
    tile[1947] = 6'd28;
    tile[1948] = 6'd28;
    tile[1949] = 6'd28;
    tile[1950] = 6'd28;
    tile[1951] = 6'd29;
    tile[1952] = 6'd10;
    tile[1953] = 6'd12;
    tile[1954] = 6'd33;
    tile[1955] = 6'd6;
    tile[1956] = 6'd6;
    tile[1957] = 6'd29;
    tile[1958] = 6'd10;
    tile[1959] = 6'd12;
    tile[1960] = 6'd11;
    tile[1961] = 6'd10;
    tile[1962] = 6'd7;
    tile[1963] = 6'd16;
    tile[1964] = 6'd16;
    tile[1965] = 6'd34;
    tile[1966] = 6'd11;
    tile[1967] = 6'd10;
    tile[1968] = 6'd27;
    tile[1969] = 6'd28;
    tile[1970] = 6'd28;
    tile[1971] = 6'd28;
    tile[1972] = 6'd25;
    tile[1973] = 6'd5;
    tile[1974] = 6'd37;
    tile[1975] = 6'd37;
    tile[1976] = 6'd37;
    tile[1977] = 6'd37;
    tile[1978] = 6'd37;
    tile[1979] = 6'd37;
    tile[1980] = 6'd37;
    tile[1981] = 6'd37;
    tile[1982] = 6'd37;
    tile[1983] = 6'd37;
    tile[1984] = 6'd37;
    tile[1985] = 6'd37;
    tile[1986] = 6'd37;
    tile[1987] = 6'd37;
    tile[1988] = 6'd37;
    tile[1989] = 6'd37;
    tile[1990] = 6'd37;
    tile[1991] = 6'd37;
    tile[1992] = 6'd37;
    tile[1993] = 6'd37;
    tile[1994] = 6'd37;
    tile[1995] = 6'd37;
    tile[1996] = 6'd37;
    tile[1997] = 6'd37;
    tile[1998] = 6'd37;
    tile[1999] = 6'd37;
    tile[2000] = 6'd37;
    tile[2001] = 6'd37;
    tile[2002] = 6'd37;
    tile[2003] = 6'd37;
    tile[2004] = 6'd37;
    tile[2005] = 6'd37;
    tile[2006] = 6'd37;
    tile[2007] = 6'd37;
    tile[2008] = 6'd37;
    tile[2009] = 6'd37;
    tile[2010] = 6'd37;
    tile[2011] = 6'd37;
    tile[2012] = 6'd37;
    tile[2013] = 6'd37;
    tile[2014] = 6'd37;
    tile[2015] = 6'd37;
    tile[2016] = 6'd37;
    tile[2017] = 6'd37;
    tile[2018] = 6'd37;
    tile[2019] = 6'd37;
    tile[2020] = 6'd37;
    tile[2021] = 6'd37;
    tile[2022] = 6'd37;
    tile[2023] = 6'd37;
    tile[2024] = 6'd37;
    tile[2025] = 6'd37;
    tile[2026] = 6'd37;
    tile[2027] = 6'd37;
    tile[2028] = 6'd37;
    tile[2029] = 6'd37;
    tile[2030] = 6'd37;
    tile[2031] = 6'd9;
    tile[2032] = 6'd10;
    tile[2033] = 6'd12;
    tile[2034] = 6'd27;
    tile[2035] = 6'd16;
    tile[2036] = 6'd16;
    tile[2037] = 6'd34;
    tile[2038] = 6'd10;
    tile[2039] = 6'd17;
    tile[2040] = 6'd18;
    tile[2041] = 6'd10;
    tile[2042] = 6'd17;
    tile[2043] = 6'd6;
    tile[2044] = 6'd6;
    tile[2045] = 6'd29;
    tile[2046] = 6'd11;
    tile[2047] = 6'd10;
    tile[2048] = 6'd13;
    tile[2049] = 6'd37;
    tile[2050] = 6'd37;
    tile[2051] = 6'd37;
    tile[2052] = 6'd37;
    tile[2053] = 6'd37;
    tile[2054] = 6'd37;
    tile[2055] = 6'd37;
    tile[2056] = 6'd37;
    tile[2057] = 6'd37;
    tile[2058] = 6'd37;
    tile[2059] = 6'd37;
    tile[2060] = 6'd37;
    tile[2061] = 6'd37;
    tile[2062] = 6'd37;
    tile[2063] = 6'd37;
    tile[2064] = 6'd37;
    tile[2065] = 6'd37;
    tile[2066] = 6'd37;
    tile[2067] = 6'd37;
    tile[2068] = 6'd37;
    tile[2069] = 6'd37;
    tile[2070] = 6'd37;
    tile[2071] = 6'd37;
    tile[2072] = 6'd37;
    tile[2073] = 6'd37;
    tile[2074] = 6'd37;
    tile[2075] = 6'd37;
    tile[2076] = 6'd37;
    tile[2077] = 6'd37;
    tile[2078] = 6'd37;
    tile[2079] = 6'd37;
    tile[2080] = 6'd37;
    tile[2081] = 6'd37;
    tile[2082] = 6'd37;
    tile[2083] = 6'd37;
    tile[2084] = 6'd37;
    tile[2085] = 6'd37;
    tile[2086] = 6'd37;
    tile[2087] = 6'd37;
    tile[2088] = 6'd37;
    tile[2089] = 6'd37;
    tile[2090] = 6'd37;
    tile[2091] = 6'd37;
    tile[2092] = 6'd37;
    tile[2093] = 6'd37;
    tile[2094] = 6'd37;
    tile[2095] = 6'd37;
    tile[2096] = 6'd37;
    tile[2097] = 6'd37;
    tile[2098] = 6'd37;
    tile[2099] = 6'd37;
    tile[2100] = 6'd37;
    tile[2101] = 6'd37;
    tile[2102] = 6'd37;
    tile[2103] = 6'd37;
    tile[2104] = 6'd37;
    tile[2105] = 6'd37;
    tile[2106] = 6'd37;
    tile[2107] = 6'd37;
    tile[2108] = 6'd37;
    tile[2109] = 6'd37;
    tile[2110] = 6'd37;
    tile[2111] = 6'd9;
    tile[2112] = 6'd10;
    tile[2113] = 6'd12;
    tile[2114] = 6'd11;
    tile[2115] = 6'd10;
    tile[2116] = 6'd10;
    tile[2117] = 6'd10;
    tile[2118] = 6'd10;
    tile[2119] = 6'd10;
    tile[2120] = 6'd10;
    tile[2121] = 6'd10;
    tile[2122] = 6'd10;
    tile[2123] = 6'd10;
    tile[2124] = 6'd10;
    tile[2125] = 6'd12;
    tile[2126] = 6'd11;
    tile[2127] = 6'd10;
    tile[2128] = 6'd13;
    tile[2129] = 6'd37;
    tile[2130] = 6'd37;
    tile[2131] = 6'd37;
    tile[2132] = 6'd37;
    tile[2133] = 6'd37;
    tile[2134] = 6'd37;
    tile[2135] = 6'd37;
    tile[2136] = 6'd37;
    tile[2137] = 6'd37;
    tile[2138] = 6'd37;
    tile[2139] = 6'd37;
    tile[2140] = 6'd37;
    tile[2141] = 6'd37;
    tile[2142] = 6'd37;
    tile[2143] = 6'd37;
    tile[2144] = 6'd37;
    tile[2145] = 6'd37;
    tile[2146] = 6'd37;
    tile[2147] = 6'd37;
    tile[2148] = 6'd37;
    tile[2149] = 6'd37;
    tile[2150] = 6'd37;
    tile[2151] = 6'd37;
    tile[2152] = 6'd37;
    tile[2153] = 6'd37;
    tile[2154] = 6'd37;
    tile[2155] = 6'd37;
    tile[2156] = 6'd37;
    tile[2157] = 6'd37;
    tile[2158] = 6'd37;
    tile[2159] = 6'd37;
    tile[2160] = 6'd37;
    tile[2161] = 6'd37;
    tile[2162] = 6'd37;
    tile[2163] = 6'd37;
    tile[2164] = 6'd37;
    tile[2165] = 6'd37;
    tile[2166] = 6'd37;
    tile[2167] = 6'd37;
    tile[2168] = 6'd37;
    tile[2169] = 6'd37;
    tile[2170] = 6'd37;
    tile[2171] = 6'd37;
    tile[2172] = 6'd37;
    tile[2173] = 6'd37;
    tile[2174] = 6'd37;
    tile[2175] = 6'd37;
    tile[2176] = 6'd37;
    tile[2177] = 6'd37;
    tile[2178] = 6'd37;
    tile[2179] = 6'd37;
    tile[2180] = 6'd37;
    tile[2181] = 6'd37;
    tile[2182] = 6'd37;
    tile[2183] = 6'd37;
    tile[2184] = 6'd37;
    tile[2185] = 6'd37;
    tile[2186] = 6'd37;
    tile[2187] = 6'd37;
    tile[2188] = 6'd37;
    tile[2189] = 6'd37;
    tile[2190] = 6'd37;
    tile[2191] = 6'd9;
    tile[2192] = 6'd10;
    tile[2193] = 6'd12;
    tile[2194] = 6'd11;
    tile[2195] = 6'd10;
    tile[2196] = 6'd23;
    tile[2197] = 6'd28;
    tile[2198] = 6'd24;
    tile[2199] = 6'd31;
    tile[2200] = 6'd31;
    tile[2201] = 6'd25;
    tile[2202] = 6'd28;
    tile[2203] = 6'd26;
    tile[2204] = 6'd10;
    tile[2205] = 6'd12;
    tile[2206] = 6'd11;
    tile[2207] = 6'd10;
    tile[2208] = 6'd13;
    tile[2209] = 6'd37;
    tile[2210] = 6'd37;
    tile[2211] = 6'd37;
    tile[2212] = 6'd37;
    tile[2213] = 6'd37;
    tile[2214] = 6'd37;
    tile[2215] = 6'd37;
    tile[2216] = 6'd37;
    tile[2217] = 6'd37;
    tile[2218] = 6'd37;
    tile[2219] = 6'd37;
    tile[2220] = 6'd37;
    tile[2221] = 6'd37;
    tile[2222] = 6'd37;
    tile[2223] = 6'd37;
    tile[2224] = 6'd37;
    tile[2225] = 6'd37;
    tile[2226] = 6'd37;
    tile[2227] = 6'd37;
    tile[2228] = 6'd37;
    tile[2229] = 6'd37;
    tile[2230] = 6'd37;
    tile[2231] = 6'd37;
    tile[2232] = 6'd37;
    tile[2233] = 6'd37;
    tile[2234] = 6'd37;
    tile[2235] = 6'd37;
    tile[2236] = 6'd37;
    tile[2237] = 6'd37;
    tile[2238] = 6'd37;
    tile[2239] = 6'd37;
    tile[2240] = 6'd37;
    tile[2241] = 6'd37;
    tile[2242] = 6'd37;
    tile[2243] = 6'd37;
    tile[2244] = 6'd37;
    tile[2245] = 6'd37;
    tile[2246] = 6'd37;
    tile[2247] = 6'd37;
    tile[2248] = 6'd37;
    tile[2249] = 6'd37;
    tile[2250] = 6'd37;
    tile[2251] = 6'd37;
    tile[2252] = 6'd37;
    tile[2253] = 6'd37;
    tile[2254] = 6'd37;
    tile[2255] = 6'd37;
    tile[2256] = 6'd37;
    tile[2257] = 6'd37;
    tile[2258] = 6'd37;
    tile[2259] = 6'd37;
    tile[2260] = 6'd37;
    tile[2261] = 6'd37;
    tile[2262] = 6'd37;
    tile[2263] = 6'd37;
    tile[2264] = 6'd37;
    tile[2265] = 6'd37;
    tile[2266] = 6'd1;
    tile[2267] = 6'd1;
    tile[2268] = 6'd1;
    tile[2269] = 6'd1;
    tile[2270] = 6'd1;
    tile[2271] = 6'd34;
    tile[2272] = 6'd10;
    tile[2273] = 6'd17;
    tile[2274] = 6'd18;
    tile[2275] = 6'd10;
    tile[2276] = 6'd13;
    tile[2277] = 6'd37;
    tile[2278] = 6'd37;
    tile[2279] = 6'd37;
    tile[2280] = 6'd37;
    tile[2281] = 6'd37;
    tile[2282] = 6'd37;
    tile[2283] = 6'd9;
    tile[2284] = 6'd10;
    tile[2285] = 6'd17;
    tile[2286] = 6'd18;
    tile[2287] = 6'd10;
    tile[2288] = 6'd33;
    tile[2289] = 6'd1;
    tile[2290] = 6'd1;
    tile[2291] = 6'd1;
    tile[2292] = 6'd1;
    tile[2293] = 6'd1;
    tile[2294] = 6'd37;
    tile[2295] = 6'd37;
    tile[2296] = 6'd37;
    tile[2297] = 6'd37;
    tile[2298] = 6'd37;
    tile[2299] = 6'd37;
    tile[2300] = 6'd37;
    tile[2301] = 6'd37;
    tile[2302] = 6'd37;
    tile[2303] = 6'd37;
    tile[2304] = 6'd37;
    tile[2305] = 6'd37;
    tile[2306] = 6'd37;
    tile[2307] = 6'd37;
    tile[2308] = 6'd37;
    tile[2309] = 6'd37;
    tile[2310] = 6'd37;
    tile[2311] = 6'd37;
    tile[2312] = 6'd37;
    tile[2313] = 6'd37;
    tile[2314] = 6'd37;
    tile[2315] = 6'd37;
    tile[2316] = 6'd37;
    tile[2317] = 6'd37;
    tile[2318] = 6'd37;
    tile[2319] = 6'd37;
    tile[2320] = 6'd37;
    tile[2321] = 6'd37;
    tile[2322] = 6'd37;
    tile[2323] = 6'd37;
    tile[2324] = 6'd37;
    tile[2325] = 6'd37;
    tile[2326] = 6'd37;
    tile[2327] = 6'd37;
    tile[2328] = 6'd37;
    tile[2329] = 6'd37;
    tile[2330] = 6'd37;
    tile[2331] = 6'd37;
    tile[2332] = 6'd37;
    tile[2333] = 6'd37;
    tile[2334] = 6'd37;
    tile[2335] = 6'd37;
    tile[2336] = 6'd37;
    tile[2337] = 6'd37;
    tile[2338] = 6'd37;
    tile[2339] = 6'd37;
    tile[2340] = 6'd37;
    tile[2341] = 6'd37;
    tile[2342] = 6'd37;
    tile[2343] = 6'd37;
    tile[2344] = 6'd37;
    tile[2345] = 6'd37;
    tile[2346] = 6'd37;
    tile[2347] = 6'd37;
    tile[2348] = 6'd37;
    tile[2349] = 6'd37;
    tile[2350] = 6'd37;
    tile[2351] = 6'd37;
    tile[2352] = 6'd37;
    tile[2353] = 6'd37;
    tile[2354] = 6'd37;
    tile[2355] = 6'd37;
    tile[2356] = 6'd13;
    tile[2357] = 6'd37;
    tile[2358] = 6'd37;
    tile[2359] = 6'd37;
    tile[2360] = 6'd37;
    tile[2361] = 6'd37;
    tile[2362] = 6'd37;
    tile[2363] = 6'd9;
    tile[2364] = 6'd37;
    tile[2365] = 6'd37;
    tile[2366] = 6'd37;
    tile[2367] = 6'd37;
    tile[2368] = 6'd37;
    tile[2369] = 6'd37;
    tile[2370] = 6'd37;
    tile[2371] = 6'd37;
    tile[2372] = 6'd37;
    tile[2373] = 6'd37;
    tile[2374] = 6'd37;
    tile[2375] = 6'd37;
    tile[2376] = 6'd37;
    tile[2377] = 6'd37;
    tile[2378] = 6'd37;
    tile[2379] = 6'd37;
    tile[2380] = 6'd37;
    tile[2381] = 6'd37;
    tile[2382] = 6'd37;
    tile[2383] = 6'd37;
    tile[2384] = 6'd37;
    tile[2385] = 6'd37;
    tile[2386] = 6'd37;
    tile[2387] = 6'd37;
    tile[2388] = 6'd37;
    tile[2389] = 6'd37;
    tile[2390] = 6'd37;
    tile[2391] = 6'd37;
    tile[2392] = 6'd37;
    tile[2393] = 6'd37;
    tile[2394] = 6'd37;
    tile[2395] = 6'd37;
    tile[2396] = 6'd37;
    tile[2397] = 6'd37;
    tile[2398] = 6'd37;
    tile[2399] = 6'd37;
    tile[2400] = 6'd37;
    tile[2401] = 6'd37;
    tile[2402] = 6'd37;
    tile[2403] = 6'd37;
    tile[2404] = 6'd37;
    tile[2405] = 6'd37;
    tile[2406] = 6'd37;
    tile[2407] = 6'd37;
    tile[2408] = 6'd37;
    tile[2409] = 6'd37;
    tile[2410] = 6'd37;
    tile[2411] = 6'd37;
    tile[2412] = 6'd37;
    tile[2413] = 6'd37;
    tile[2414] = 6'd37;
    tile[2415] = 6'd37;
    tile[2416] = 6'd37;
    tile[2417] = 6'd37;
    tile[2418] = 6'd37;
    tile[2419] = 6'd37;
    tile[2420] = 6'd37;
    tile[2421] = 6'd37;
    tile[2422] = 6'd37;
    tile[2423] = 6'd37;
    tile[2424] = 6'd37;
    tile[2425] = 6'd37;
    tile[2426] = 6'd28;
    tile[2427] = 6'd28;
    tile[2428] = 6'd28;
    tile[2429] = 6'd28;
    tile[2430] = 6'd28;
    tile[2431] = 6'd29;
    tile[2432] = 6'd10;
    tile[2433] = 6'd7;
    tile[2434] = 6'd8;
    tile[2435] = 6'd13;
    tile[2436] = 6'd37;
    tile[2437] = 6'd37;
    tile[2438] = 6'd37;
    tile[2439] = 6'd37;
    tile[2440] = 6'd37;
    tile[2441] = 6'd37;
    tile[2442] = 6'd37;
    tile[2443] = 6'd9;
    tile[2444] = 6'd10;
    tile[2445] = 6'd7;
    tile[2446] = 6'd8;
    tile[2447] = 6'd10;
    tile[2448] = 6'd27;
    tile[2449] = 6'd28;
    tile[2450] = 6'd28;
    tile[2451] = 6'd28;
    tile[2452] = 6'd28;
    tile[2453] = 6'd28;
    tile[2454] = 6'd37;
    tile[2455] = 6'd37;
    tile[2456] = 6'd37;
    tile[2457] = 6'd37;
    tile[2458] = 6'd37;
    tile[2459] = 6'd37;
    tile[2460] = 6'd37;
    tile[2461] = 6'd37;
    tile[2462] = 6'd37;
    tile[2463] = 6'd37;
    tile[2464] = 6'd37;
    tile[2465] = 6'd37;
    tile[2466] = 6'd37;
    tile[2467] = 6'd37;
    tile[2468] = 6'd37;
    tile[2469] = 6'd37;
    tile[2470] = 6'd37;
    tile[2471] = 6'd37;
    tile[2472] = 6'd37;
    tile[2473] = 6'd37;
    tile[2474] = 6'd37;
    tile[2475] = 6'd37;
    tile[2476] = 6'd37;
    tile[2477] = 6'd37;
    tile[2478] = 6'd37;
    tile[2479] = 6'd37;
    tile[2480] = 6'd37;
    tile[2481] = 6'd37;
    tile[2482] = 6'd37;
    tile[2483] = 6'd37;
    tile[2484] = 6'd37;
    tile[2485] = 6'd37;
    tile[2486] = 6'd37;
    tile[2487] = 6'd37;
    tile[2488] = 6'd37;
    tile[2489] = 6'd37;
    tile[2490] = 6'd37;
    tile[2491] = 6'd37;
    tile[2492] = 6'd37;
    tile[2493] = 6'd37;
    tile[2494] = 6'd37;
    tile[2495] = 6'd37;
    tile[2496] = 6'd37;
    tile[2497] = 6'd37;
    tile[2498] = 6'd37;
    tile[2499] = 6'd37;
    tile[2500] = 6'd37;
    tile[2501] = 6'd37;
    tile[2502] = 6'd37;
    tile[2503] = 6'd37;
    tile[2504] = 6'd37;
    tile[2505] = 6'd37;
    tile[2506] = 6'd37;
    tile[2507] = 6'd37;
    tile[2508] = 6'd37;
    tile[2509] = 6'd37;
    tile[2510] = 6'd37;
    tile[2511] = 6'd9;
    tile[2512] = 6'd10;
    tile[2513] = 6'd12;
    tile[2514] = 6'd11;
    tile[2515] = 6'd10;
    tile[2516] = 6'd30;
    tile[2517] = 6'd28;
    tile[2518] = 6'd28;
    tile[2519] = 6'd28;
    tile[2520] = 6'd28;
    tile[2521] = 6'd28;
    tile[2522] = 6'd28;
    tile[2523] = 6'd32;
    tile[2524] = 6'd10;
    tile[2525] = 6'd12;
    tile[2526] = 6'd11;
    tile[2527] = 6'd10;
    tile[2528] = 6'd13;
    tile[2529] = 6'd37;
    tile[2530] = 6'd37;
    tile[2531] = 6'd37;
    tile[2532] = 6'd37;
    tile[2533] = 6'd37;
    tile[2534] = 6'd37;
    tile[2535] = 6'd37;
    tile[2536] = 6'd37;
    tile[2537] = 6'd37;
    tile[2538] = 6'd37;
    tile[2539] = 6'd37;
    tile[2540] = 6'd37;
    tile[2541] = 6'd37;
    tile[2542] = 6'd37;
    tile[2543] = 6'd37;
    tile[2544] = 6'd37;
    tile[2545] = 6'd37;
    tile[2546] = 6'd37;
    tile[2547] = 6'd37;
    tile[2548] = 6'd37;
    tile[2549] = 6'd37;
    tile[2550] = 6'd37;
    tile[2551] = 6'd37;
    tile[2552] = 6'd37;
    tile[2553] = 6'd37;
    tile[2554] = 6'd37;
    tile[2555] = 6'd37;
    tile[2556] = 6'd37;
    tile[2557] = 6'd37;
    tile[2558] = 6'd37;
    tile[2559] = 6'd37;
    tile[2560] = 6'd37;
    tile[2561] = 6'd37;
    tile[2562] = 6'd37;
    tile[2563] = 6'd37;
    tile[2564] = 6'd37;
    tile[2565] = 6'd37;
    tile[2566] = 6'd37;
    tile[2567] = 6'd37;
    tile[2568] = 6'd37;
    tile[2569] = 6'd37;
    tile[2570] = 6'd37;
    tile[2571] = 6'd37;
    tile[2572] = 6'd37;
    tile[2573] = 6'd37;
    tile[2574] = 6'd37;
    tile[2575] = 6'd37;
    tile[2576] = 6'd37;
    tile[2577] = 6'd37;
    tile[2578] = 6'd37;
    tile[2579] = 6'd37;
    tile[2580] = 6'd37;
    tile[2581] = 6'd37;
    tile[2582] = 6'd37;
    tile[2583] = 6'd37;
    tile[2584] = 6'd37;
    tile[2585] = 6'd37;
    tile[2586] = 6'd37;
    tile[2587] = 6'd37;
    tile[2588] = 6'd37;
    tile[2589] = 6'd37;
    tile[2590] = 6'd37;
    tile[2591] = 6'd9;
    tile[2592] = 6'd10;
    tile[2593] = 6'd12;
    tile[2594] = 6'd11;
    tile[2595] = 6'd10;
    tile[2596] = 6'd37;
    tile[2597] = 6'd37;
    tile[2598] = 6'd37;
    tile[2599] = 6'd37;
    tile[2600] = 6'd37;
    tile[2601] = 6'd37;
    tile[2602] = 6'd37;
    tile[2603] = 6'd37;
    tile[2604] = 6'd10;
    tile[2605] = 6'd12;
    tile[2606] = 6'd11;
    tile[2607] = 6'd10;
    tile[2608] = 6'd13;
    tile[2609] = 6'd37;
    tile[2610] = 6'd37;
    tile[2611] = 6'd37;
    tile[2612] = 6'd37;
    tile[2613] = 6'd37;
    tile[2614] = 6'd37;
    tile[2615] = 6'd37;
    tile[2616] = 6'd37;
    tile[2617] = 6'd37;
    tile[2618] = 6'd37;
    tile[2619] = 6'd37;
    tile[2620] = 6'd37;
    tile[2621] = 6'd37;
    tile[2622] = 6'd37;
    tile[2623] = 6'd37;
    tile[2624] = 6'd37;
    tile[2625] = 6'd37;
    tile[2626] = 6'd37;
    tile[2627] = 6'd37;
    tile[2628] = 6'd37;
    tile[2629] = 6'd37;
    tile[2630] = 6'd37;
    tile[2631] = 6'd37;
    tile[2632] = 6'd37;
    tile[2633] = 6'd37;
    tile[2634] = 6'd37;
    tile[2635] = 6'd37;
    tile[2636] = 6'd37;
    tile[2637] = 6'd37;
    tile[2638] = 6'd37;
    tile[2639] = 6'd37;
    tile[2640] = 6'd37;
    tile[2641] = 6'd37;
    tile[2642] = 6'd37;
    tile[2643] = 6'd37;
    tile[2644] = 6'd37;
    tile[2645] = 6'd37;
    tile[2646] = 6'd37;
    tile[2647] = 6'd37;
    tile[2648] = 6'd37;
    tile[2649] = 6'd37;
    tile[2650] = 6'd37;
    tile[2651] = 6'd37;
    tile[2652] = 6'd37;
    tile[2653] = 6'd37;
    tile[2654] = 6'd37;
    tile[2655] = 6'd37;
    tile[2656] = 6'd37;
    tile[2657] = 6'd37;
    tile[2658] = 6'd37;
    tile[2659] = 6'd37;
    tile[2660] = 6'd37;
    tile[2661] = 6'd37;
    tile[2662] = 6'd37;
    tile[2663] = 6'd37;
    tile[2664] = 6'd37;
    tile[2665] = 6'd37;
    tile[2666] = 6'd37;
    tile[2667] = 6'd37;
    tile[2668] = 6'd37;
    tile[2669] = 6'd37;
    tile[2670] = 6'd37;
    tile[2671] = 6'd9;
    tile[2672] = 6'd10;
    tile[2673] = 6'd12;
    tile[2674] = 6'd11;
    tile[2675] = 6'd10;
    tile[2676] = 6'd7;
    tile[2677] = 6'd16;
    tile[2678] = 6'd16;
    tile[2679] = 6'd16;
    tile[2680] = 6'd16;
    tile[2681] = 6'd16;
    tile[2682] = 6'd16;
    tile[2683] = 6'd8;
    tile[2684] = 6'd10;
    tile[2685] = 6'd12;
    tile[2686] = 6'd11;
    tile[2687] = 6'd10;
    tile[2688] = 6'd13;
    tile[2689] = 6'd37;
    tile[2690] = 6'd37;
    tile[2691] = 6'd37;
    tile[2692] = 6'd37;
    tile[2693] = 6'd37;
    tile[2694] = 6'd37;
    tile[2695] = 6'd37;
    tile[2696] = 6'd37;
    tile[2697] = 6'd37;
    tile[2698] = 6'd37;
    tile[2699] = 6'd37;
    tile[2700] = 6'd37;
    tile[2701] = 6'd37;
    tile[2702] = 6'd37;
    tile[2703] = 6'd37;
    tile[2704] = 6'd37;
    tile[2705] = 6'd37;
    tile[2706] = 6'd37;
    tile[2707] = 6'd37;
    tile[2708] = 6'd37;
    tile[2709] = 6'd37;
    tile[2710] = 6'd37;
    tile[2711] = 6'd37;
    tile[2712] = 6'd37;
    tile[2713] = 6'd37;
    tile[2714] = 6'd37;
    tile[2715] = 6'd37;
    tile[2716] = 6'd37;
    tile[2717] = 6'd37;
    tile[2718] = 6'd37;
    tile[2719] = 6'd37;
    tile[2720] = 6'd37;
    tile[2721] = 6'd37;
    tile[2722] = 6'd37;
    tile[2723] = 6'd37;
    tile[2724] = 6'd37;
    tile[2725] = 6'd37;
    tile[2726] = 6'd37;
    tile[2727] = 6'd37;
    tile[2728] = 6'd37;
    tile[2729] = 6'd37;
    tile[2730] = 6'd37;
    tile[2731] = 6'd37;
    tile[2732] = 6'd37;
    tile[2733] = 6'd37;
    tile[2734] = 6'd37;
    tile[2735] = 6'd37;
    tile[2736] = 6'd37;
    tile[2737] = 6'd37;
    tile[2738] = 6'd37;
    tile[2739] = 6'd37;
    tile[2740] = 6'd37;
    tile[2741] = 6'd37;
    tile[2742] = 6'd37;
    tile[2743] = 6'd37;
    tile[2744] = 6'd37;
    tile[2745] = 6'd37;
    tile[2746] = 6'd0;
    tile[2747] = 6'd1;
    tile[2748] = 6'd1;
    tile[2749] = 6'd1;
    tile[2750] = 6'd1;
    tile[2751] = 6'd34;
    tile[2752] = 6'd10;
    tile[2753] = 6'd17;
    tile[2754] = 6'd18;
    tile[2755] = 6'd10;
    tile[2756] = 6'd17;
    tile[2757] = 6'd6;
    tile[2758] = 6'd6;
    tile[2759] = 6'd29;
    tile[2760] = 6'd27;
    tile[2761] = 6'd6;
    tile[2762] = 6'd6;
    tile[2763] = 6'd18;
    tile[2764] = 6'd10;
    tile[2765] = 6'd17;
    tile[2766] = 6'd18;
    tile[2767] = 6'd10;
    tile[2768] = 6'd33;
    tile[2769] = 6'd1;
    tile[2770] = 6'd1;
    tile[2771] = 6'd1;
    tile[2772] = 6'd1;
    tile[2773] = 6'd4;
    tile[2774] = 6'd37;
    tile[2775] = 6'd37;
    tile[2776] = 6'd37;
    tile[2777] = 6'd37;
    tile[2778] = 6'd37;
    tile[2779] = 6'd37;
    tile[2780] = 6'd37;
    tile[2781] = 6'd37;
    tile[2782] = 6'd37;
    tile[2783] = 6'd37;
    tile[2784] = 6'd37;
    tile[2785] = 6'd37;
    tile[2786] = 6'd37;
    tile[2787] = 6'd37;
    tile[2788] = 6'd37;
    tile[2789] = 6'd37;
    tile[2790] = 6'd37;
    tile[2791] = 6'd37;
    tile[2792] = 6'd37;
    tile[2793] = 6'd37;
    tile[2794] = 6'd37;
    tile[2795] = 6'd37;
    tile[2796] = 6'd37;
    tile[2797] = 6'd37;
    tile[2798] = 6'd37;
    tile[2799] = 6'd37;
    tile[2800] = 6'd37;
    tile[2801] = 6'd37;
    tile[2802] = 6'd37;
    tile[2803] = 6'd37;
    tile[2804] = 6'd37;
    tile[2805] = 6'd37;
    tile[2806] = 6'd37;
    tile[2807] = 6'd37;
    tile[2808] = 6'd37;
    tile[2809] = 6'd37;
    tile[2810] = 6'd37;
    tile[2811] = 6'd37;
    tile[2812] = 6'd37;
    tile[2813] = 6'd37;
    tile[2814] = 6'd37;
    tile[2815] = 6'd37;
    tile[2816] = 6'd37;
    tile[2817] = 6'd37;
    tile[2818] = 6'd37;
    tile[2819] = 6'd37;
    tile[2820] = 6'd37;
    tile[2821] = 6'd37;
    tile[2822] = 6'd37;
    tile[2823] = 6'd37;
    tile[2824] = 6'd37;
    tile[2825] = 6'd37;
    tile[2826] = 6'd9;
    tile[2827] = 6'd10;
    tile[2828] = 6'd10;
    tile[2829] = 6'd10;
    tile[2830] = 6'd10;
    tile[2831] = 6'd10;
    tile[2832] = 6'd10;
    tile[2833] = 6'd10;
    tile[2834] = 6'd10;
    tile[2835] = 6'd10;
    tile[2836] = 6'd10;
    tile[2837] = 6'd10;
    tile[2838] = 6'd10;
    tile[2839] = 6'd11;
    tile[2840] = 6'd12;
    tile[2841] = 6'd10;
    tile[2842] = 6'd10;
    tile[2843] = 6'd10;
    tile[2844] = 6'd10;
    tile[2845] = 6'd10;
    tile[2846] = 6'd10;
    tile[2847] = 6'd10;
    tile[2848] = 6'd10;
    tile[2849] = 6'd10;
    tile[2850] = 6'd10;
    tile[2851] = 6'd10;
    tile[2852] = 6'd10;
    tile[2853] = 6'd13;
    tile[2854] = 6'd37;
    tile[2855] = 6'd37;
    tile[2856] = 6'd37;
    tile[2857] = 6'd37;
    tile[2858] = 6'd37;
    tile[2859] = 6'd37;
    tile[2860] = 6'd37;
    tile[2861] = 6'd37;
    tile[2862] = 6'd37;
    tile[2863] = 6'd37;
    tile[2864] = 6'd37;
    tile[2865] = 6'd37;
    tile[2866] = 6'd37;
    tile[2867] = 6'd37;
    tile[2868] = 6'd37;
    tile[2869] = 6'd37;
    tile[2870] = 6'd37;
    tile[2871] = 6'd37;
    tile[2872] = 6'd37;
    tile[2873] = 6'd37;
    tile[2874] = 6'd37;
    tile[2875] = 6'd37;
    tile[2876] = 6'd37;
    tile[2877] = 6'd37;
    tile[2878] = 6'd37;
    tile[2879] = 6'd37;
    tile[2880] = 6'd37;
    tile[2881] = 6'd37;
    tile[2882] = 6'd37;
    tile[2883] = 6'd37;
    tile[2884] = 6'd37;
    tile[2885] = 6'd37;
    tile[2886] = 6'd37;
    tile[2887] = 6'd37;
    tile[2888] = 6'd37;
    tile[2889] = 6'd37;
    tile[2890] = 6'd37;
    tile[2891] = 6'd37;
    tile[2892] = 6'd37;
    tile[2893] = 6'd37;
    tile[2894] = 6'd37;
    tile[2895] = 6'd37;
    tile[2896] = 6'd37;
    tile[2897] = 6'd37;
    tile[2898] = 6'd37;
    tile[2899] = 6'd37;
    tile[2900] = 6'd37;
    tile[2901] = 6'd37;
    tile[2902] = 6'd37;
    tile[2903] = 6'd37;
    tile[2904] = 6'd37;
    tile[2905] = 6'd37;
    tile[2906] = 6'd9;
    tile[2907] = 6'd10;
    tile[2908] = 6'd7;
    tile[2909] = 6'd16;
    tile[2910] = 6'd16;
    tile[2911] = 6'd8;
    tile[2912] = 6'd10;
    tile[2913] = 6'd7;
    tile[2914] = 6'd16;
    tile[2915] = 6'd16;
    tile[2916] = 6'd16;
    tile[2917] = 6'd8;
    tile[2918] = 6'd10;
    tile[2919] = 6'd11;
    tile[2920] = 6'd12;
    tile[2921] = 6'd10;
    tile[2922] = 6'd7;
    tile[2923] = 6'd16;
    tile[2924] = 6'd16;
    tile[2925] = 6'd16;
    tile[2926] = 6'd8;
    tile[2927] = 6'd10;
    tile[2928] = 6'd7;
    tile[2929] = 6'd16;
    tile[2930] = 6'd16;
    tile[2931] = 6'd8;
    tile[2932] = 6'd10;
    tile[2933] = 6'd13;
    tile[2934] = 6'd37;
    tile[2935] = 6'd37;
    tile[2936] = 6'd37;
    tile[2937] = 6'd37;
    tile[2938] = 6'd37;
    tile[2939] = 6'd37;
    tile[2940] = 6'd37;
    tile[2941] = 6'd37;
    tile[2942] = 6'd37;
    tile[2943] = 6'd37;
    tile[2944] = 6'd37;
    tile[2945] = 6'd37;
    tile[2946] = 6'd37;
    tile[2947] = 6'd37;
    tile[2948] = 6'd37;
    tile[2949] = 6'd37;
    tile[2950] = 6'd37;
    tile[2951] = 6'd37;
    tile[2952] = 6'd37;
    tile[2953] = 6'd37;
    tile[2954] = 6'd37;
    tile[2955] = 6'd37;
    tile[2956] = 6'd37;
    tile[2957] = 6'd37;
    tile[2958] = 6'd37;
    tile[2959] = 6'd37;
    tile[2960] = 6'd37;
    tile[2961] = 6'd37;
    tile[2962] = 6'd37;
    tile[2963] = 6'd37;
    tile[2964] = 6'd37;
    tile[2965] = 6'd37;
    tile[2966] = 6'd37;
    tile[2967] = 6'd37;
    tile[2968] = 6'd37;
    tile[2969] = 6'd37;
    tile[2970] = 6'd37;
    tile[2971] = 6'd37;
    tile[2972] = 6'd37;
    tile[2973] = 6'd37;
    tile[2974] = 6'd37;
    tile[2975] = 6'd37;
    tile[2976] = 6'd37;
    tile[2977] = 6'd37;
    tile[2978] = 6'd37;
    tile[2979] = 6'd37;
    tile[2980] = 6'd37;
    tile[2981] = 6'd37;
    tile[2982] = 6'd37;
    tile[2983] = 6'd37;
    tile[2984] = 6'd37;
    tile[2985] = 6'd37;
    tile[2986] = 6'd9;
    tile[2987] = 6'd10;
    tile[2988] = 6'd17;
    tile[2989] = 6'd6;
    tile[2990] = 6'd29;
    tile[2991] = 6'd11;
    tile[2992] = 6'd10;
    tile[2993] = 6'd17;
    tile[2994] = 6'd6;
    tile[2995] = 6'd6;
    tile[2996] = 6'd6;
    tile[2997] = 6'd18;
    tile[2998] = 6'd10;
    tile[2999] = 6'd33;
    tile[3000] = 6'd34;
    tile[3001] = 6'd10;
    tile[3002] = 6'd17;
    tile[3003] = 6'd6;
    tile[3004] = 6'd6;
    tile[3005] = 6'd6;
    tile[3006] = 6'd18;
    tile[3007] = 6'd10;
    tile[3008] = 6'd12;
    tile[3009] = 6'd27;
    tile[3010] = 6'd6;
    tile[3011] = 6'd18;
    tile[3012] = 6'd10;
    tile[3013] = 6'd13;
    tile[3014] = 6'd37;
    tile[3015] = 6'd37;
    tile[3016] = 6'd37;
    tile[3017] = 6'd37;
    tile[3018] = 6'd37;
    tile[3019] = 6'd37;
    tile[3020] = 6'd37;
    tile[3021] = 6'd37;
    tile[3022] = 6'd37;
    tile[3023] = 6'd37;
    tile[3024] = 6'd37;
    tile[3025] = 6'd37;
    tile[3026] = 6'd37;
    tile[3027] = 6'd37;
    tile[3028] = 6'd37;
    tile[3029] = 6'd37;
    tile[3030] = 6'd37;
    tile[3031] = 6'd37;
    tile[3032] = 6'd37;
    tile[3033] = 6'd37;
    tile[3034] = 6'd37;
    tile[3035] = 6'd37;
    tile[3036] = 6'd37;
    tile[3037] = 6'd37;
    tile[3038] = 6'd37;
    tile[3039] = 6'd37;
    tile[3040] = 6'd37;
    tile[3041] = 6'd37;
    tile[3042] = 6'd37;
    tile[3043] = 6'd37;
    tile[3044] = 6'd37;
    tile[3045] = 6'd37;
    tile[3046] = 6'd37;
    tile[3047] = 6'd37;
    tile[3048] = 6'd37;
    tile[3049] = 6'd37;
    tile[3050] = 6'd37;
    tile[3051] = 6'd37;
    tile[3052] = 6'd37;
    tile[3053] = 6'd37;
    tile[3054] = 6'd37;
    tile[3055] = 6'd37;
    tile[3056] = 6'd37;
    tile[3057] = 6'd37;
    tile[3058] = 6'd37;
    tile[3059] = 6'd37;
    tile[3060] = 6'd37;
    tile[3061] = 6'd37;
    tile[3062] = 6'd37;
    tile[3063] = 6'd37;
    tile[3064] = 6'd37;
    tile[3065] = 6'd37;
    tile[3066] = 6'd9;
    tile[3067] = 6'd10;
    tile[3068] = 6'd10;
    tile[3069] = 6'd10;
    tile[3070] = 6'd12;
    tile[3071] = 6'd11;
    tile[3072] = 6'd10;
    tile[3073] = 6'd10;
    tile[3074] = 6'd10;
    tile[3075] = 6'd10;
    tile[3076] = 6'd10;
    tile[3077] = 6'd10;
    tile[3078] = 6'd10;
    tile[3079] = 6'd10;
    tile[3080] = 6'd10;
    tile[3081] = 6'd10;
    tile[3082] = 6'd10;
    tile[3083] = 6'd10;
    tile[3084] = 6'd10;
    tile[3085] = 6'd10;
    tile[3086] = 6'd10;
    tile[3087] = 6'd10;
    tile[3088] = 6'd12;
    tile[3089] = 6'd11;
    tile[3090] = 6'd10;
    tile[3091] = 6'd10;
    tile[3092] = 6'd10;
    tile[3093] = 6'd13;
    tile[3094] = 6'd37;
    tile[3095] = 6'd37;
    tile[3096] = 6'd37;
    tile[3097] = 6'd37;
    tile[3098] = 6'd37;
    tile[3099] = 6'd37;
    tile[3100] = 6'd37;
    tile[3101] = 6'd37;
    tile[3102] = 6'd37;
    tile[3103] = 6'd37;
    tile[3104] = 6'd37;
    tile[3105] = 6'd37;
    tile[3106] = 6'd37;
    tile[3107] = 6'd37;
    tile[3108] = 6'd37;
    tile[3109] = 6'd37;
    tile[3110] = 6'd37;
    tile[3111] = 6'd37;
    tile[3112] = 6'd37;
    tile[3113] = 6'd37;
    tile[3114] = 6'd37;
    tile[3115] = 6'd37;
    tile[3116] = 6'd37;
    tile[3117] = 6'd37;
    tile[3118] = 6'd37;
    tile[3119] = 6'd37;
    tile[3120] = 6'd37;
    tile[3121] = 6'd37;
    tile[3122] = 6'd37;
    tile[3123] = 6'd37;
    tile[3124] = 6'd37;
    tile[3125] = 6'd37;
    tile[3126] = 6'd37;
    tile[3127] = 6'd37;
    tile[3128] = 6'd37;
    tile[3129] = 6'd37;
    tile[3130] = 6'd37;
    tile[3131] = 6'd37;
    tile[3132] = 6'd37;
    tile[3133] = 6'd37;
    tile[3134] = 6'd37;
    tile[3135] = 6'd37;
    tile[3136] = 6'd37;
    tile[3137] = 6'd37;
    tile[3138] = 6'd37;
    tile[3139] = 6'd37;
    tile[3140] = 6'd37;
    tile[3141] = 6'd37;
    tile[3142] = 6'd37;
    tile[3143] = 6'd37;
    tile[3144] = 6'd37;
    tile[3145] = 6'd37;
    tile[3146] = 6'd15;
    tile[3147] = 6'd6;
    tile[3148] = 6'd8;
    tile[3149] = 6'd10;
    tile[3150] = 6'd12;
    tile[3151] = 6'd11;
    tile[3152] = 6'd10;
    tile[3153] = 6'd7;
    tile[3154] = 6'd8;
    tile[3155] = 6'd10;
    tile[3156] = 6'd7;
    tile[3157] = 6'd10;
    tile[3158] = 6'd10;
    tile[3159] = 6'd10;
    tile[3160] = 6'd10;
    tile[3161] = 6'd10;
    tile[3162] = 6'd10;
    tile[3163] = 6'd8;
    tile[3164] = 6'd10;
    tile[3165] = 6'd7;
    tile[3166] = 6'd8;
    tile[3167] = 6'd10;
    tile[3168] = 6'd12;
    tile[3169] = 6'd11;
    tile[3170] = 6'd10;
    tile[3171] = 6'd27;
    tile[3172] = 6'd6;
    tile[3173] = 6'd14;
    tile[3174] = 6'd37;
    tile[3175] = 6'd37;
    tile[3176] = 6'd37;
    tile[3177] = 6'd37;
    tile[3178] = 6'd37;
    tile[3179] = 6'd37;
    tile[3180] = 6'd37;
    tile[3181] = 6'd37;
    tile[3182] = 6'd37;
    tile[3183] = 6'd37;
    tile[3184] = 6'd37;
    tile[3185] = 6'd37;
    tile[3186] = 6'd37;
    tile[3187] = 6'd37;
    tile[3188] = 6'd37;
    tile[3189] = 6'd37;
    tile[3190] = 6'd37;
    tile[3191] = 6'd37;
    tile[3192] = 6'd37;
    tile[3193] = 6'd37;
    tile[3194] = 6'd37;
    tile[3195] = 6'd37;
    tile[3196] = 6'd37;
    tile[3197] = 6'd37;
    tile[3198] = 6'd37;
    tile[3199] = 6'd37;
    tile[3200] = 6'd37;
    tile[3201] = 6'd37;
    tile[3202] = 6'd37;
    tile[3203] = 6'd37;
    tile[3204] = 6'd37;
    tile[3205] = 6'd37;
    tile[3206] = 6'd37;
    tile[3207] = 6'd37;
    tile[3208] = 6'd37;
    tile[3209] = 6'd37;
    tile[3210] = 6'd37;
    tile[3211] = 6'd37;
    tile[3212] = 6'd37;
    tile[3213] = 6'd37;
    tile[3214] = 6'd37;
    tile[3215] = 6'd37;
    tile[3216] = 6'd37;
    tile[3217] = 6'd37;
    tile[3218] = 6'd37;
    tile[3219] = 6'd37;
    tile[3220] = 6'd37;
    tile[3221] = 6'd37;
    tile[3222] = 6'd37;
    tile[3223] = 6'd37;
    tile[3224] = 6'd37;
    tile[3225] = 6'd37;
    tile[3226] = 6'd35;
    tile[3227] = 6'd16;
    tile[3228] = 6'd18;
    tile[3229] = 6'd10;
    tile[3230] = 6'd17;
    tile[3231] = 6'd18;
    tile[3232] = 6'd10;
    tile[3233] = 6'd12;
    tile[3234] = 6'd11;
    tile[3235] = 6'd10;
    tile[3236] = 6'd17;
    tile[3237] = 6'd6;
    tile[3238] = 6'd6;
    tile[3239] = 6'd29;
    tile[3240] = 6'd27;
    tile[3241] = 6'd6;
    tile[3242] = 6'd6;
    tile[3243] = 6'd18;
    tile[3244] = 6'd10;
    tile[3245] = 6'd12;
    tile[3246] = 6'd11;
    tile[3247] = 6'd10;
    tile[3248] = 6'd17;
    tile[3249] = 6'd18;
    tile[3250] = 6'd10;
    tile[3251] = 6'd33;
    tile[3252] = 6'd16;
    tile[3253] = 6'd36;
    tile[3254] = 6'd37;
    tile[3255] = 6'd37;
    tile[3256] = 6'd37;
    tile[3257] = 6'd37;
    tile[3258] = 6'd37;
    tile[3259] = 6'd37;
    tile[3260] = 6'd37;
    tile[3261] = 6'd37;
    tile[3262] = 6'd37;
    tile[3263] = 6'd37;
    tile[3264] = 6'd37;
    tile[3265] = 6'd37;
    tile[3266] = 6'd37;
    tile[3267] = 6'd37;
    tile[3268] = 6'd37;
    tile[3269] = 6'd37;
    tile[3270] = 6'd37;
    tile[3271] = 6'd37;
    tile[3272] = 6'd37;
    tile[3273] = 6'd37;
    tile[3274] = 6'd37;
    tile[3275] = 6'd37;
    tile[3276] = 6'd37;
    tile[3277] = 6'd37;
    tile[3278] = 6'd37;
    tile[3279] = 6'd37;
    tile[3280] = 6'd37;
    tile[3281] = 6'd37;
    tile[3282] = 6'd37;
    tile[3283] = 6'd37;
    tile[3284] = 6'd37;
    tile[3285] = 6'd37;
    tile[3286] = 6'd37;
    tile[3287] = 6'd37;
    tile[3288] = 6'd37;
    tile[3289] = 6'd37;
    tile[3290] = 6'd37;
    tile[3291] = 6'd37;
    tile[3292] = 6'd37;
    tile[3293] = 6'd37;
    tile[3294] = 6'd37;
    tile[3295] = 6'd37;
    tile[3296] = 6'd37;
    tile[3297] = 6'd37;
    tile[3298] = 6'd37;
    tile[3299] = 6'd37;
    tile[3300] = 6'd37;
    tile[3301] = 6'd37;
    tile[3302] = 6'd37;
    tile[3303] = 6'd37;
    tile[3304] = 6'd37;
    tile[3305] = 6'd37;
    tile[3306] = 6'd9;
    tile[3307] = 6'd10;
    tile[3308] = 6'd10;
    tile[3309] = 6'd10;
    tile[3310] = 6'd10;
    tile[3311] = 6'd10;
    tile[3312] = 6'd10;
    tile[3313] = 6'd12;
    tile[3314] = 6'd11;
    tile[3315] = 6'd10;
    tile[3316] = 6'd10;
    tile[3317] = 6'd10;
    tile[3318] = 6'd10;
    tile[3319] = 6'd11;
    tile[3320] = 6'd12;
    tile[3321] = 6'd10;
    tile[3322] = 6'd10;
    tile[3323] = 6'd10;
    tile[3324] = 6'd10;
    tile[3325] = 6'd12;
    tile[3326] = 6'd11;
    tile[3327] = 6'd10;
    tile[3328] = 6'd10;
    tile[3329] = 6'd10;
    tile[3330] = 6'd10;
    tile[3331] = 6'd10;
    tile[3332] = 6'd10;
    tile[3333] = 6'd13;
    tile[3334] = 6'd37;
    tile[3335] = 6'd37;
    tile[3336] = 6'd37;
    tile[3337] = 6'd37;
    tile[3338] = 6'd37;
    tile[3339] = 6'd37;
    tile[3340] = 6'd37;
    tile[3341] = 6'd37;
    tile[3342] = 6'd37;
    tile[3343] = 6'd37;
    tile[3344] = 6'd37;
    tile[3345] = 6'd37;
    tile[3346] = 6'd37;
    tile[3347] = 6'd37;
    tile[3348] = 6'd37;
    tile[3349] = 6'd37;
    tile[3350] = 6'd37;
    tile[3351] = 6'd37;
    tile[3352] = 6'd37;
    tile[3353] = 6'd37;
    tile[3354] = 6'd37;
    tile[3355] = 6'd37;
    tile[3356] = 6'd37;
    tile[3357] = 6'd37;
    tile[3358] = 6'd37;
    tile[3359] = 6'd37;
    tile[3360] = 6'd37;
    tile[3361] = 6'd37;
    tile[3362] = 6'd37;
    tile[3363] = 6'd37;
    tile[3364] = 6'd37;
    tile[3365] = 6'd37;
    tile[3366] = 6'd37;
    tile[3367] = 6'd37;
    tile[3368] = 6'd37;
    tile[3369] = 6'd37;
    tile[3370] = 6'd37;
    tile[3371] = 6'd37;
    tile[3372] = 6'd37;
    tile[3373] = 6'd37;
    tile[3374] = 6'd37;
    tile[3375] = 6'd37;
    tile[3376] = 6'd37;
    tile[3377] = 6'd37;
    tile[3378] = 6'd37;
    tile[3379] = 6'd37;
    tile[3380] = 6'd37;
    tile[3381] = 6'd37;
    tile[3382] = 6'd37;
    tile[3383] = 6'd37;
    tile[3384] = 6'd37;
    tile[3385] = 6'd37;
    tile[3386] = 6'd9;
    tile[3387] = 6'd10;
    tile[3388] = 6'd7;
    tile[3389] = 6'd16;
    tile[3390] = 6'd16;
    tile[3391] = 6'd16;
    tile[3392] = 6'd16;
    tile[3393] = 6'd34;
    tile[3394] = 6'd33;
    tile[3395] = 6'd16;
    tile[3396] = 6'd16;
    tile[3397] = 6'd8;
    tile[3398] = 6'd10;
    tile[3399] = 6'd11;
    tile[3400] = 6'd12;
    tile[3401] = 6'd10;
    tile[3402] = 6'd7;
    tile[3403] = 6'd16;
    tile[3404] = 6'd16;
    tile[3405] = 6'd34;
    tile[3406] = 6'd33;
    tile[3407] = 6'd16;
    tile[3408] = 6'd16;
    tile[3409] = 6'd16;
    tile[3410] = 6'd16;
    tile[3411] = 6'd8;
    tile[3412] = 6'd10;
    tile[3413] = 6'd13;
    tile[3414] = 6'd37;
    tile[3415] = 6'd37;
    tile[3416] = 6'd37;
    tile[3417] = 6'd37;
    tile[3418] = 6'd37;
    tile[3419] = 6'd37;
    tile[3420] = 6'd37;
    tile[3421] = 6'd37;
    tile[3422] = 6'd37;
    tile[3423] = 6'd37;
    tile[3424] = 6'd37;
    tile[3425] = 6'd37;
    tile[3426] = 6'd37;
    tile[3427] = 6'd37;
    tile[3428] = 6'd37;
    tile[3429] = 6'd37;
    tile[3430] = 6'd37;
    tile[3431] = 6'd37;
    tile[3432] = 6'd37;
    tile[3433] = 6'd37;
    tile[3434] = 6'd37;
    tile[3435] = 6'd37;
    tile[3436] = 6'd37;
    tile[3437] = 6'd37;
    tile[3438] = 6'd37;
    tile[3439] = 6'd37;
    tile[3440] = 6'd37;
    tile[3441] = 6'd37;
    tile[3442] = 6'd37;
    tile[3443] = 6'd37;
    tile[3444] = 6'd37;
    tile[3445] = 6'd37;
    tile[3446] = 6'd37;
    tile[3447] = 6'd37;
    tile[3448] = 6'd37;
    tile[3449] = 6'd37;
    tile[3450] = 6'd37;
    tile[3451] = 6'd37;
    tile[3452] = 6'd37;
    tile[3453] = 6'd37;
    tile[3454] = 6'd37;
    tile[3455] = 6'd37;
    tile[3456] = 6'd37;
    tile[3457] = 6'd37;
    tile[3458] = 6'd37;
    tile[3459] = 6'd37;
    tile[3460] = 6'd37;
    tile[3461] = 6'd37;
    tile[3462] = 6'd37;
    tile[3463] = 6'd37;
    tile[3464] = 6'd37;
    tile[3465] = 6'd37;
    tile[3466] = 6'd9;
    tile[3467] = 6'd10;
    tile[3468] = 6'd17;
    tile[3469] = 6'd6;
    tile[3470] = 6'd6;
    tile[3471] = 6'd6;
    tile[3472] = 6'd6;
    tile[3473] = 6'd6;
    tile[3474] = 6'd6;
    tile[3475] = 6'd6;
    tile[3476] = 6'd6;
    tile[3477] = 6'd18;
    tile[3478] = 6'd10;
    tile[3479] = 6'd33;
    tile[3480] = 6'd34;
    tile[3481] = 6'd10;
    tile[3482] = 6'd17;
    tile[3483] = 6'd6;
    tile[3484] = 6'd6;
    tile[3485] = 6'd6;
    tile[3486] = 6'd6;
    tile[3487] = 6'd6;
    tile[3488] = 6'd6;
    tile[3489] = 6'd6;
    tile[3490] = 6'd6;
    tile[3491] = 6'd18;
    tile[3492] = 6'd10;
    tile[3493] = 6'd13;
    tile[3494] = 6'd37;
    tile[3495] = 6'd37;
    tile[3496] = 6'd37;
    tile[3497] = 6'd37;
    tile[3498] = 6'd37;
    tile[3499] = 6'd37;
    tile[3500] = 6'd37;
    tile[3501] = 6'd37;
    tile[3502] = 6'd37;
    tile[3503] = 6'd37;
    tile[3504] = 6'd37;
    tile[3505] = 6'd37;
    tile[3506] = 6'd37;
    tile[3507] = 6'd37;
    tile[3508] = 6'd37;
    tile[3509] = 6'd37;
    tile[3510] = 6'd37;
    tile[3511] = 6'd37;
    tile[3512] = 6'd37;
    tile[3513] = 6'd37;
    tile[3514] = 6'd37;
    tile[3515] = 6'd37;
    tile[3516] = 6'd37;
    tile[3517] = 6'd37;
    tile[3518] = 6'd37;
    tile[3519] = 6'd37;
    tile[3520] = 6'd37;
    tile[3521] = 6'd37;
    tile[3522] = 6'd37;
    tile[3523] = 6'd37;
    tile[3524] = 6'd37;
    tile[3525] = 6'd37;
    tile[3526] = 6'd37;
    tile[3527] = 6'd37;
    tile[3528] = 6'd37;
    tile[3529] = 6'd37;
    tile[3530] = 6'd37;
    tile[3531] = 6'd37;
    tile[3532] = 6'd37;
    tile[3533] = 6'd37;
    tile[3534] = 6'd37;
    tile[3535] = 6'd37;
    tile[3536] = 6'd37;
    tile[3537] = 6'd37;
    tile[3538] = 6'd37;
    tile[3539] = 6'd37;
    tile[3540] = 6'd37;
    tile[3541] = 6'd37;
    tile[3542] = 6'd37;
    tile[3543] = 6'd37;
    tile[3544] = 6'd37;
    tile[3545] = 6'd37;
    tile[3546] = 6'd9;
    tile[3547] = 6'd10;
    tile[3548] = 6'd10;
    tile[3549] = 6'd10;
    tile[3550] = 6'd10;
    tile[3551] = 6'd10;
    tile[3552] = 6'd10;
    tile[3553] = 6'd10;
    tile[3554] = 6'd10;
    tile[3555] = 6'd10;
    tile[3556] = 6'd10;
    tile[3557] = 6'd10;
    tile[3558] = 6'd10;
    tile[3559] = 6'd10;
    tile[3560] = 6'd10;
    tile[3561] = 6'd10;
    tile[3562] = 6'd10;
    tile[3563] = 6'd10;
    tile[3564] = 6'd10;
    tile[3565] = 6'd10;
    tile[3566] = 6'd10;
    tile[3567] = 6'd10;
    tile[3568] = 6'd10;
    tile[3569] = 6'd10;
    tile[3570] = 6'd10;
    tile[3571] = 6'd10;
    tile[3572] = 6'd10;
    tile[3573] = 6'd13;
    tile[3574] = 6'd37;
    tile[3575] = 6'd37;
    tile[3576] = 6'd37;
    tile[3577] = 6'd37;
    tile[3578] = 6'd37;
    tile[3579] = 6'd37;
    tile[3580] = 6'd37;
    tile[3581] = 6'd37;
    tile[3582] = 6'd37;
    tile[3583] = 6'd37;
    tile[3584] = 6'd37;
    tile[3585] = 6'd37;
    tile[3586] = 6'd37;
    tile[3587] = 6'd37;
    tile[3588] = 6'd37;
    tile[3589] = 6'd37;
    tile[3590] = 6'd37;
    tile[3591] = 6'd37;
    tile[3592] = 6'd37;
    tile[3593] = 6'd37;
    tile[3594] = 6'd37;
    tile[3595] = 6'd37;
    tile[3596] = 6'd37;
    tile[3597] = 6'd37;
    tile[3598] = 6'd37;
    tile[3599] = 6'd37;
    tile[3600] = 6'd37;
    tile[3601] = 6'd37;
    tile[3602] = 6'd37;
    tile[3603] = 6'd37;
    tile[3604] = 6'd37;
    tile[3605] = 6'd37;
    tile[3606] = 6'd37;
    tile[3607] = 6'd37;
    tile[3608] = 6'd37;
    tile[3609] = 6'd37;
    tile[3610] = 6'd37;
    tile[3611] = 6'd37;
    tile[3612] = 6'd37;
    tile[3613] = 6'd37;
    tile[3614] = 6'd37;
    tile[3615] = 6'd37;
    tile[3616] = 6'd37;
    tile[3617] = 6'd37;
    tile[3618] = 6'd37;
    tile[3619] = 6'd37;
    tile[3620] = 6'd37;
    tile[3621] = 6'd37;
    tile[3622] = 6'd37;
    tile[3623] = 6'd37;
    tile[3624] = 6'd37;
    tile[3625] = 6'd37;
    tile[3626] = 6'd19;
    tile[3627] = 6'd1;
    tile[3628] = 6'd1;
    tile[3629] = 6'd1;
    tile[3630] = 6'd1;
    tile[3631] = 6'd1;
    tile[3632] = 6'd1;
    tile[3633] = 6'd1;
    tile[3634] = 6'd1;
    tile[3635] = 6'd1;
    tile[3636] = 6'd1;
    tile[3637] = 6'd1;
    tile[3638] = 6'd1;
    tile[3639] = 6'd1;
    tile[3640] = 6'd1;
    tile[3641] = 6'd1;
    tile[3642] = 6'd1;
    tile[3643] = 6'd1;
    tile[3644] = 6'd1;
    tile[3645] = 6'd1;
    tile[3646] = 6'd1;
    tile[3647] = 6'd1;
    tile[3648] = 6'd1;
    tile[3649] = 6'd1;
    tile[3650] = 6'd1;
    tile[3651] = 6'd1;
    tile[3652] = 6'd1;
    tile[3653] = 6'd5;
    tile[3654] = 6'd37;
    tile[3655] = 6'd37;
    tile[3656] = 6'd37;
    tile[3657] = 6'd37;
    tile[3658] = 6'd37;
    tile[3659] = 6'd37;
    tile[3660] = 6'd37;
    tile[3661] = 6'd37;
    tile[3662] = 6'd37;
    tile[3663] = 6'd37;
    tile[3664] = 6'd37;
    tile[3665] = 6'd37;
    tile[3666] = 6'd37;
    tile[3667] = 6'd37;
    tile[3668] = 6'd37;
    tile[3669] = 6'd37;
    tile[3670] = 6'd37;
    tile[3671] = 6'd37;
    tile[3672] = 6'd37;
    tile[3673] = 6'd37;
    tile[3674] = 6'd37;
    tile[3675] = 6'd37;
    tile[3676] = 6'd37;
    tile[3677] = 6'd37;
    tile[3678] = 6'd37;
    tile[3679] = 6'd37;
    tile[3680] = 6'd37;
    tile[3681] = 6'd37;
    tile[3682] = 6'd37;
    tile[3683] = 6'd37;
    tile[3684] = 6'd37;
    tile[3685] = 6'd37;
    tile[3686] = 6'd37;
    tile[3687] = 6'd37;
    tile[3688] = 6'd37;
    tile[3689] = 6'd37;
    tile[3690] = 6'd37;
    tile[3691] = 6'd37;
    tile[3692] = 6'd37;
    tile[3693] = 6'd37;
    tile[3694] = 6'd37;
    tile[3695] = 6'd37;
    tile[3696] = 6'd37;
    tile[3697] = 6'd37;
    tile[3698] = 6'd37;
    tile[3699] = 6'd37;
    tile[3700] = 6'd37;
    tile[3701] = 6'd37;
    tile[3702] = 6'd37;
    tile[3703] = 6'd37;
    tile[3704] = 6'd37;
    tile[3705] = 6'd37;
    tile[3706] = 6'd37;
    tile[3707] = 6'd37;
    tile[3708] = 6'd37;
    tile[3709] = 6'd37;
    tile[3710] = 6'd37;
    tile[3711] = 6'd37;
    tile[3712] = 6'd37;
    tile[3713] = 6'd37;
    tile[3714] = 6'd37;
    tile[3715] = 6'd37;
    tile[3716] = 6'd37;
    tile[3717] = 6'd37;
    tile[3718] = 6'd37;
    tile[3719] = 6'd37;
    tile[3720] = 6'd37;
    tile[3721] = 6'd37;
    tile[3722] = 6'd37;
    tile[3723] = 6'd37;
    tile[3724] = 6'd37;
    tile[3725] = 6'd37;
    tile[3726] = 6'd37;
    tile[3727] = 6'd37;
    tile[3728] = 6'd37;
    tile[3729] = 6'd37;
    tile[3730] = 6'd37;
    tile[3731] = 6'd37;
    tile[3732] = 6'd37;
    tile[3733] = 6'd37;
    tile[3734] = 6'd37;
    tile[3735] = 6'd37;
    tile[3736] = 6'd37;
    tile[3737] = 6'd37;
    tile[3738] = 6'd37;
    tile[3739] = 6'd37;
    tile[3740] = 6'd37;
    tile[3741] = 6'd37;
    tile[3742] = 6'd37;
    tile[3743] = 6'd37;
    tile[3744] = 6'd37;
    tile[3745] = 6'd37;
    tile[3746] = 6'd37;
    tile[3747] = 6'd37;
    tile[3748] = 6'd37;
    tile[3749] = 6'd37;
    tile[3750] = 6'd37;
    tile[3751] = 6'd37;
    tile[3752] = 6'd37;
    tile[3753] = 6'd37;
    tile[3754] = 6'd37;
    tile[3755] = 6'd37;
    tile[3756] = 6'd37;
    tile[3757] = 6'd37;
    tile[3758] = 6'd37;
    tile[3759] = 6'd37;
    tile[3760] = 6'd37;
    tile[3761] = 6'd37;
    tile[3762] = 6'd37;
    tile[3763] = 6'd37;
    tile[3764] = 6'd37;
    tile[3765] = 6'd37;
    tile[3766] = 6'd37;
    tile[3767] = 6'd37;
    tile[3768] = 6'd37;
    tile[3769] = 6'd37;
    tile[3770] = 6'd37;
    tile[3771] = 6'd37;
    tile[3772] = 6'd37;
    tile[3773] = 6'd37;
    tile[3774] = 6'd37;
    tile[3775] = 6'd37;
    tile[3776] = 6'd37;
    tile[3777] = 6'd37;
    tile[3778] = 6'd37;
    tile[3779] = 6'd37;
    tile[3780] = 6'd37;
    tile[3781] = 6'd37;
    tile[3782] = 6'd37;
    tile[3783] = 6'd37;
    tile[3784] = 6'd37;
    tile[3785] = 6'd37;
    tile[3786] = 6'd37;
    tile[3787] = 6'd37;
    tile[3788] = 6'd37;
    tile[3789] = 6'd37;
    tile[3790] = 6'd37;
    tile[3791] = 6'd37;
    tile[3792] = 6'd37;
    tile[3793] = 6'd37;
    tile[3794] = 6'd37;
    tile[3795] = 6'd37;
    tile[3796] = 6'd37;
    tile[3797] = 6'd37;
    tile[3798] = 6'd37;
    tile[3799] = 6'd37;
    tile[3800] = 6'd37;
    tile[3801] = 6'd37;
    tile[3802] = 6'd37;
    tile[3803] = 6'd37;
    tile[3804] = 6'd37;
    tile[3805] = 6'd37;
    tile[3806] = 6'd37;
    tile[3807] = 6'd37;
    tile[3808] = 6'd37;
    tile[3809] = 6'd37;
    tile[3810] = 6'd37;
    tile[3811] = 6'd37;
    tile[3812] = 6'd37;
    tile[3813] = 6'd37;
    tile[3814] = 6'd37;
    tile[3815] = 6'd37;
    tile[3816] = 6'd37;
    tile[3817] = 6'd37;
    tile[3818] = 6'd37;
    tile[3819] = 6'd37;
    tile[3820] = 6'd37;
    tile[3821] = 6'd37;
    tile[3822] = 6'd37;
    tile[3823] = 6'd37;
    tile[3824] = 6'd37;
    tile[3825] = 6'd37;
    tile[3826] = 6'd37;
    tile[3827] = 6'd37;
    tile[3828] = 6'd37;
    tile[3829] = 6'd37;
    tile[3830] = 6'd37;
    tile[3831] = 6'd37;
    tile[3832] = 6'd37;
    tile[3833] = 6'd37;
    tile[3834] = 6'd37;
    tile[3835] = 6'd37;
    tile[3836] = 6'd37;
    tile[3837] = 6'd37;
    tile[3838] = 6'd37;
    tile[3839] = 6'd37;
    tile[3840] = 6'd37;
    tile[3841] = 6'd37;
    tile[3842] = 6'd37;
    tile[3843] = 6'd37;
    tile[3844] = 6'd37;
    tile[3845] = 6'd37;
    tile[3846] = 6'd37;
    tile[3847] = 6'd37;
    tile[3848] = 6'd37;
    tile[3849] = 6'd37;
    tile[3850] = 6'd37;
    tile[3851] = 6'd37;
    tile[3852] = 6'd37;
    tile[3853] = 6'd37;
    tile[3854] = 6'd37;
    tile[3855] = 6'd37;
    tile[3856] = 6'd37;
    tile[3857] = 6'd37;
    tile[3858] = 6'd37;
    tile[3859] = 6'd37;
    tile[3860] = 6'd37;
    tile[3861] = 6'd37;
    tile[3862] = 6'd37;
    tile[3863] = 6'd37;
    tile[3864] = 6'd37;
    tile[3865] = 6'd37;
    tile[3866] = 6'd37;
    tile[3867] = 6'd37;
    tile[3868] = 6'd37;
    tile[3869] = 6'd37;
    tile[3870] = 6'd37;
    tile[3871] = 6'd37;
    tile[3872] = 6'd37;
    tile[3873] = 6'd37;
    tile[3874] = 6'd37;
    tile[3875] = 6'd37;
    tile[3876] = 6'd37;
    tile[3877] = 6'd37;
    tile[3878] = 6'd37;
    tile[3879] = 6'd37;
    tile[3880] = 6'd37;
    tile[3881] = 6'd37;
    tile[3882] = 6'd37;
    tile[3883] = 6'd37;
    tile[3884] = 6'd37;
    tile[3885] = 6'd37;
    tile[3886] = 6'd37;
    tile[3887] = 6'd37;
    tile[3888] = 6'd37;
    tile[3889] = 6'd37;
    tile[3890] = 6'd37;
    tile[3891] = 6'd37;
    tile[3892] = 6'd37;
    tile[3893] = 6'd37;
    tile[3894] = 6'd37;
    tile[3895] = 6'd37;
    tile[3896] = 6'd37;
    tile[3897] = 6'd37;
    tile[3898] = 6'd37;
    tile[3899] = 6'd37;
    tile[3900] = 6'd37;
    tile[3901] = 6'd37;
    tile[3902] = 6'd37;
    tile[3903] = 6'd37;
    tile[3904] = 6'd37;
    tile[3905] = 6'd37;
    tile[3906] = 6'd37;
    tile[3907] = 6'd37;
    tile[3908] = 6'd37;
    tile[3909] = 6'd37;
    tile[3910] = 6'd37;
    tile[3911] = 6'd37;
    tile[3912] = 6'd37;
    tile[3913] = 6'd37;
    tile[3914] = 6'd37;
    tile[3915] = 6'd37;
    tile[3916] = 6'd37;
    tile[3917] = 6'd37;
    tile[3918] = 6'd37;
    tile[3919] = 6'd37;
    tile[3920] = 6'd37;
    tile[3921] = 6'd37;
    tile[3922] = 6'd37;
    tile[3923] = 6'd37;
    tile[3924] = 6'd37;
    tile[3925] = 6'd37;
    tile[3926] = 6'd37;
    tile[3927] = 6'd37;
    tile[3928] = 6'd37;
    tile[3929] = 6'd37;
    tile[3930] = 6'd37;
    tile[3931] = 6'd37;
    tile[3932] = 6'd37;
    tile[3933] = 6'd37;
    tile[3934] = 6'd37;
    tile[3935] = 6'd37;
    tile[3936] = 6'd37;
    tile[3937] = 6'd37;
    tile[3938] = 6'd37;
    tile[3939] = 6'd37;
    tile[3940] = 6'd37;
    tile[3941] = 6'd37;
    tile[3942] = 6'd37;
    tile[3943] = 6'd37;
    tile[3944] = 6'd37;
    tile[3945] = 6'd37;
    tile[3946] = 6'd37;
    tile[3947] = 6'd37;
    tile[3948] = 6'd37;
    tile[3949] = 6'd37;
    tile[3950] = 6'd37;
    tile[3951] = 6'd37;
    tile[3952] = 6'd37;
    tile[3953] = 6'd37;
    tile[3954] = 6'd37;
    tile[3955] = 6'd37;
    tile[3956] = 6'd37;
    tile[3957] = 6'd37;
    tile[3958] = 6'd37;
    tile[3959] = 6'd37;
    tile[3960] = 6'd37;
    tile[3961] = 6'd37;
    tile[3962] = 6'd37;
    tile[3963] = 6'd37;
    tile[3964] = 6'd37;
    tile[3965] = 6'd37;
    tile[3966] = 6'd37;
    tile[3967] = 6'd37;
    tile[3968] = 6'd37;
    tile[3969] = 6'd37;
    tile[3970] = 6'd37;
    tile[3971] = 6'd37;
    tile[3972] = 6'd37;
    tile[3973] = 6'd37;
    tile[3974] = 6'd37;
    tile[3975] = 6'd37;
    tile[3976] = 6'd37;
    tile[3977] = 6'd37;
    tile[3978] = 6'd37;
    tile[3979] = 6'd37;
    tile[3980] = 6'd37;
    tile[3981] = 6'd37;
    tile[3982] = 6'd37;
    tile[3983] = 6'd37;
    tile[3984] = 6'd37;
    tile[3985] = 6'd37;
    tile[3986] = 6'd37;
    tile[3987] = 6'd37;
    tile[3988] = 6'd37;
    tile[3989] = 6'd37;
    tile[3990] = 6'd37;
    tile[3991] = 6'd37;
    tile[3992] = 6'd37;
    tile[3993] = 6'd37;
    tile[3994] = 6'd37;
    tile[3995] = 6'd37;
    tile[3996] = 6'd37;
    tile[3997] = 6'd37;
    tile[3998] = 6'd37;
    tile[3999] = 6'd37;
    tile[4000] = 6'd37;
    tile[4001] = 6'd37;
    tile[4002] = 6'd37;
    tile[4003] = 6'd37;
    tile[4004] = 6'd37;
    tile[4005] = 6'd37;
    tile[4006] = 6'd37;
    tile[4007] = 6'd37;
    tile[4008] = 6'd37;
    tile[4009] = 6'd37;
    tile[4010] = 6'd37;
    tile[4011] = 6'd37;
    tile[4012] = 6'd37;
    tile[4013] = 6'd37;
    tile[4014] = 6'd37;
    tile[4015] = 6'd37;
    tile[4016] = 6'd37;
    tile[4017] = 6'd37;
    tile[4018] = 6'd37;
    tile[4019] = 6'd37;
    tile[4020] = 6'd37;
    tile[4021] = 6'd37;
    tile[4022] = 6'd37;
    tile[4023] = 6'd37;
    tile[4024] = 6'd37;
    tile[4025] = 6'd37;
    tile[4026] = 6'd37;
    tile[4027] = 6'd37;
    tile[4028] = 6'd37;
    tile[4029] = 6'd37;
    tile[4030] = 6'd37;
    tile[4031] = 6'd37;
    tile[4032] = 6'd37;
    tile[4033] = 6'd37;
    tile[4034] = 6'd37;
    tile[4035] = 6'd37;
    tile[4036] = 6'd37;
    tile[4037] = 6'd37;
    tile[4038] = 6'd37;
    tile[4039] = 6'd37;
    tile[4040] = 6'd37;
    tile[4041] = 6'd37;
    tile[4042] = 6'd37;
    tile[4043] = 6'd37;
    tile[4044] = 6'd37;
    tile[4045] = 6'd37;
    tile[4046] = 6'd37;
    tile[4047] = 6'd37;
    tile[4048] = 6'd37;
    tile[4049] = 6'd37;
    tile[4050] = 6'd37;
    tile[4051] = 6'd37;
    tile[4052] = 6'd37;
    tile[4053] = 6'd37;
    tile[4054] = 6'd37;
    tile[4055] = 6'd37;
    tile[4056] = 6'd37;
    tile[4057] = 6'd37;
    tile[4058] = 6'd37;
    tile[4059] = 6'd37;
    tile[4060] = 6'd37;
    tile[4061] = 6'd37;
    tile[4062] = 6'd37;
    tile[4063] = 6'd37;
    tile[4064] = 6'd37;
    tile[4065] = 6'd37;
    tile[4066] = 6'd37;
    tile[4067] = 6'd37;
    tile[4068] = 6'd37;
    tile[4069] = 6'd37;
    tile[4070] = 6'd37;
    tile[4071] = 6'd37;
    tile[4072] = 6'd37;
    tile[4073] = 6'd37;
    tile[4074] = 6'd37;
    tile[4075] = 6'd37;
    tile[4076] = 6'd37;
    tile[4077] = 6'd37;
    tile[4078] = 6'd37;
    tile[4079] = 6'd37;
    tile[4080] = 6'd37;
    tile[4081] = 6'd37;
    tile[4082] = 6'd37;
    tile[4083] = 6'd37;
    tile[4084] = 6'd37;
    tile[4085] = 6'd37;
    tile[4086] = 6'd37;
    tile[4087] = 6'd37;
    tile[4088] = 6'd37;
    tile[4089] = 6'd37;
    tile[4090] = 6'd37;
    tile[4091] = 6'd37;
    tile[4092] = 6'd37;
    tile[4093] = 6'd37;
    tile[4094] = 6'd37;
    tile[4095] = 6'd37;
    tile[4096] = 6'd37;
    tile[4097] = 6'd37;
    tile[4098] = 6'd37;
    tile[4099] = 6'd37;
    tile[4100] = 6'd37;
    tile[4101] = 6'd37;
    tile[4102] = 6'd37;
    tile[4103] = 6'd37;
    tile[4104] = 6'd37;
    tile[4105] = 6'd37;
    tile[4106] = 6'd37;
    tile[4107] = 6'd37;
    tile[4108] = 6'd37;
    tile[4109] = 6'd37;
    tile[4110] = 6'd37;
    tile[4111] = 6'd37;
    tile[4112] = 6'd37;
    tile[4113] = 6'd37;
    tile[4114] = 6'd37;
    tile[4115] = 6'd37;
    tile[4116] = 6'd37;
    tile[4117] = 6'd37;
    tile[4118] = 6'd37;
    tile[4119] = 6'd37;
    tile[4120] = 6'd37;
    tile[4121] = 6'd37;
    tile[4122] = 6'd37;
    tile[4123] = 6'd37;
    tile[4124] = 6'd37;
    tile[4125] = 6'd37;
    tile[4126] = 6'd37;
    tile[4127] = 6'd37;
    tile[4128] = 6'd37;
    tile[4129] = 6'd37;
    tile[4130] = 6'd37;
    tile[4131] = 6'd37;
    tile[4132] = 6'd37;
    tile[4133] = 6'd37;
    tile[4134] = 6'd37;
    tile[4135] = 6'd37;
    tile[4136] = 6'd37;
    tile[4137] = 6'd37;
    tile[4138] = 6'd37;
    tile[4139] = 6'd37;
    tile[4140] = 6'd37;
    tile[4141] = 6'd37;
    tile[4142] = 6'd37;
    tile[4143] = 6'd37;
    tile[4144] = 6'd37;
    tile[4145] = 6'd37;
    tile[4146] = 6'd37;
    tile[4147] = 6'd37;
    tile[4148] = 6'd37;
    tile[4149] = 6'd37;
    tile[4150] = 6'd37;
    tile[4151] = 6'd37;
    tile[4152] = 6'd37;
    tile[4153] = 6'd37;
    tile[4154] = 6'd37;
    tile[4155] = 6'd37;
    tile[4156] = 6'd37;
    tile[4157] = 6'd37;
    tile[4158] = 6'd37;
    tile[4159] = 6'd37;
    tile[4160] = 6'd37;
    tile[4161] = 6'd37;
    tile[4162] = 6'd37;
    tile[4163] = 6'd37;
    tile[4164] = 6'd37;
    tile[4165] = 6'd37;
    tile[4166] = 6'd37;
    tile[4167] = 6'd37;
    tile[4168] = 6'd37;
    tile[4169] = 6'd37;
    tile[4170] = 6'd37;
    tile[4171] = 6'd37;
    tile[4172] = 6'd37;
    tile[4173] = 6'd37;
    tile[4174] = 6'd37;
    tile[4175] = 6'd37;
    tile[4176] = 6'd37;
    tile[4177] = 6'd37;
    tile[4178] = 6'd37;
    tile[4179] = 6'd37;
    tile[4180] = 6'd37;
    tile[4181] = 6'd37;
    tile[4182] = 6'd37;
    tile[4183] = 6'd37;
    tile[4184] = 6'd37;
    tile[4185] = 6'd37;
    tile[4186] = 6'd37;
    tile[4187] = 6'd37;
    tile[4188] = 6'd37;
    tile[4189] = 6'd37;
    tile[4190] = 6'd37;
    tile[4191] = 6'd37;
    tile[4192] = 6'd37;
    tile[4193] = 6'd37;
    tile[4194] = 6'd37;
    tile[4195] = 6'd37;
    tile[4196] = 6'd37;
    tile[4197] = 6'd37;
    tile[4198] = 6'd37;
    tile[4199] = 6'd37;
    tile[4200] = 6'd37;
    tile[4201] = 6'd37;
    tile[4202] = 6'd37;
    tile[4203] = 6'd37;
    tile[4204] = 6'd37;
    tile[4205] = 6'd37;
    tile[4206] = 6'd37;
    tile[4207] = 6'd37;
    tile[4208] = 6'd37;
    tile[4209] = 6'd37;
    tile[4210] = 6'd37;
    tile[4211] = 6'd37;
    tile[4212] = 6'd37;
    tile[4213] = 6'd37;
    tile[4214] = 6'd37;
    tile[4215] = 6'd37;
    tile[4216] = 6'd37;
    tile[4217] = 6'd37;
    tile[4218] = 6'd37;
    tile[4219] = 6'd37;
    tile[4220] = 6'd37;
    tile[4221] = 6'd37;
    tile[4222] = 6'd37;
    tile[4223] = 6'd37;
    tile[4224] = 6'd37;
    tile[4225] = 6'd37;
    tile[4226] = 6'd37;
    tile[4227] = 6'd37;
    tile[4228] = 6'd37;
    tile[4229] = 6'd37;
    tile[4230] = 6'd37;
    tile[4231] = 6'd37;
    tile[4232] = 6'd37;
    tile[4233] = 6'd37;
    tile[4234] = 6'd37;
    tile[4235] = 6'd37;
    tile[4236] = 6'd37;
    tile[4237] = 6'd37;
    tile[4238] = 6'd37;
    tile[4239] = 6'd37;
    tile[4240] = 6'd37;
    tile[4241] = 6'd37;
    tile[4242] = 6'd37;
    tile[4243] = 6'd37;
    tile[4244] = 6'd37;
    tile[4245] = 6'd37;
    tile[4246] = 6'd37;
    tile[4247] = 6'd37;
    tile[4248] = 6'd37;
    tile[4249] = 6'd37;
    tile[4250] = 6'd37;
    tile[4251] = 6'd37;
    tile[4252] = 6'd37;
    tile[4253] = 6'd37;
    tile[4254] = 6'd37;
    tile[4255] = 6'd37;
    tile[4256] = 6'd37;
    tile[4257] = 6'd37;
    tile[4258] = 6'd37;
    tile[4259] = 6'd37;
    tile[4260] = 6'd37;
    tile[4261] = 6'd37;
    tile[4262] = 6'd37;
    tile[4263] = 6'd37;
    tile[4264] = 6'd37;
    tile[4265] = 6'd37;
    tile[4266] = 6'd37;
    tile[4267] = 6'd37;
    tile[4268] = 6'd37;
    tile[4269] = 6'd37;
    tile[4270] = 6'd37;
    tile[4271] = 6'd37;
    tile[4272] = 6'd37;
    tile[4273] = 6'd37;
    tile[4274] = 6'd37;
    tile[4275] = 6'd37;
    tile[4276] = 6'd37;
    tile[4277] = 6'd37;
    tile[4278] = 6'd37;
    tile[4279] = 6'd37;
    tile[4280] = 6'd37;
    tile[4281] = 6'd37;
    tile[4282] = 6'd37;
    tile[4283] = 6'd37;
    tile[4284] = 6'd37;
    tile[4285] = 6'd37;
    tile[4286] = 6'd37;
    tile[4287] = 6'd37;
    tile[4288] = 6'd37;
    tile[4289] = 6'd37;
    tile[4290] = 6'd37;
    tile[4291] = 6'd37;
    tile[4292] = 6'd37;
    tile[4293] = 6'd37;
    tile[4294] = 6'd37;
    tile[4295] = 6'd37;
    tile[4296] = 6'd37;
    tile[4297] = 6'd37;
    tile[4298] = 6'd37;
    tile[4299] = 6'd37;
    tile[4300] = 6'd37;
    tile[4301] = 6'd37;
    tile[4302] = 6'd37;
    tile[4303] = 6'd37;
    tile[4304] = 6'd37;
    tile[4305] = 6'd37;
    tile[4306] = 6'd37;
    tile[4307] = 6'd37;
    tile[4308] = 6'd37;
    tile[4309] = 6'd37;
    tile[4310] = 6'd37;
    tile[4311] = 6'd37;
    tile[4312] = 6'd37;
    tile[4313] = 6'd37;
    tile[4314] = 6'd37;
    tile[4315] = 6'd37;
    tile[4316] = 6'd37;
    tile[4317] = 6'd37;
    tile[4318] = 6'd37;
    tile[4319] = 6'd37;
    tile[4320] = 6'd37;
    tile[4321] = 6'd37;
    tile[4322] = 6'd37;
    tile[4323] = 6'd37;
    tile[4324] = 6'd37;
    tile[4325] = 6'd37;
    tile[4326] = 6'd37;
    tile[4327] = 6'd37;
    tile[4328] = 6'd37;
    tile[4329] = 6'd37;
    tile[4330] = 6'd37;
    tile[4331] = 6'd37;
    tile[4332] = 6'd37;
    tile[4333] = 6'd37;
    tile[4334] = 6'd37;
    tile[4335] = 6'd37;
    tile[4336] = 6'd37;
    tile[4337] = 6'd37;
    tile[4338] = 6'd37;
    tile[4339] = 6'd37;
    tile[4340] = 6'd37;
    tile[4341] = 6'd37;
    tile[4342] = 6'd37;
    tile[4343] = 6'd37;
    tile[4344] = 6'd37;
    tile[4345] = 6'd37;
    tile[4346] = 6'd37;
    tile[4347] = 6'd37;
    tile[4348] = 6'd37;
    tile[4349] = 6'd37;
    tile[4350] = 6'd37;
    tile[4351] = 6'd37;
    tile[4352] = 6'd37;
    tile[4353] = 6'd37;
    tile[4354] = 6'd37;
    tile[4355] = 6'd37;
    tile[4356] = 6'd37;
    tile[4357] = 6'd37;
    tile[4358] = 6'd37;
    tile[4359] = 6'd37;
    tile[4360] = 6'd37;
    tile[4361] = 6'd37;
    tile[4362] = 6'd37;
    tile[4363] = 6'd37;
    tile[4364] = 6'd37;
    tile[4365] = 6'd37;
    tile[4366] = 6'd37;
    tile[4367] = 6'd37;
    tile[4368] = 6'd37;
    tile[4369] = 6'd37;
    tile[4370] = 6'd37;
    tile[4371] = 6'd37;
    tile[4372] = 6'd37;
    tile[4373] = 6'd37;
    tile[4374] = 6'd37;
    tile[4375] = 6'd37;
    tile[4376] = 6'd37;
    tile[4377] = 6'd37;
    tile[4378] = 6'd37;
    tile[4379] = 6'd37;
    tile[4380] = 6'd37;
    tile[4381] = 6'd37;
    tile[4382] = 6'd37;
    tile[4383] = 6'd37;
    tile[4384] = 6'd37;
    tile[4385] = 6'd37;
    tile[4386] = 6'd37;
    tile[4387] = 6'd37;
    tile[4388] = 6'd37;
    tile[4389] = 6'd37;
    tile[4390] = 6'd37;
    tile[4391] = 6'd37;
    tile[4392] = 6'd37;
    tile[4393] = 6'd37;
    tile[4394] = 6'd37;
    tile[4395] = 6'd37;
    tile[4396] = 6'd37;
    tile[4397] = 6'd37;
    tile[4398] = 6'd37;
    tile[4399] = 6'd37;
    tile[4400] = 6'd37;
    tile[4401] = 6'd37;
    tile[4402] = 6'd37;
    tile[4403] = 6'd37;
    tile[4404] = 6'd37;
    tile[4405] = 6'd37;
    tile[4406] = 6'd37;
    tile[4407] = 6'd37;
    tile[4408] = 6'd37;
    tile[4409] = 6'd37;
    tile[4410] = 6'd37;
    tile[4411] = 6'd37;
    tile[4412] = 6'd37;
    tile[4413] = 6'd37;
    tile[4414] = 6'd37;
    tile[4415] = 6'd37;
    tile[4416] = 6'd37;
    tile[4417] = 6'd37;
    tile[4418] = 6'd37;
    tile[4419] = 6'd37;
    tile[4420] = 6'd37;
    tile[4421] = 6'd37;
    tile[4422] = 6'd37;
    tile[4423] = 6'd37;
    tile[4424] = 6'd37;
    tile[4425] = 6'd37;
    tile[4426] = 6'd37;
    tile[4427] = 6'd37;
    tile[4428] = 6'd37;
    tile[4429] = 6'd37;
    tile[4430] = 6'd37;
    tile[4431] = 6'd37;
    tile[4432] = 6'd37;
    tile[4433] = 6'd37;
    tile[4434] = 6'd37;
    tile[4435] = 6'd37;
    tile[4436] = 6'd37;
    tile[4437] = 6'd37;
    tile[4438] = 6'd37;
    tile[4439] = 6'd37;
    tile[4440] = 6'd37;
    tile[4441] = 6'd37;
    tile[4442] = 6'd37;
    tile[4443] = 6'd37;
    tile[4444] = 6'd37;
    tile[4445] = 6'd37;
    tile[4446] = 6'd37;
    tile[4447] = 6'd37;
    tile[4448] = 6'd37;
    tile[4449] = 6'd37;
    tile[4450] = 6'd37;
    tile[4451] = 6'd37;
    tile[4452] = 6'd37;
    tile[4453] = 6'd37;
    tile[4454] = 6'd37;
    tile[4455] = 6'd37;
    tile[4456] = 6'd37;
    tile[4457] = 6'd37;
    tile[4458] = 6'd37;
    tile[4459] = 6'd37;
    tile[4460] = 6'd37;
    tile[4461] = 6'd37;
    tile[4462] = 6'd37;
    tile[4463] = 6'd37;
    tile[4464] = 6'd37;
    tile[4465] = 6'd37;
    tile[4466] = 6'd37;
    tile[4467] = 6'd37;
    tile[4468] = 6'd37;
    tile[4469] = 6'd37;
    tile[4470] = 6'd37;
    tile[4471] = 6'd37;
    tile[4472] = 6'd37;
    tile[4473] = 6'd37;
    tile[4474] = 6'd37;
    tile[4475] = 6'd37;
    tile[4476] = 6'd37;
    tile[4477] = 6'd37;
    tile[4478] = 6'd37;
    tile[4479] = 6'd37;
    tile[4480] = 6'd37;
    tile[4481] = 6'd37;
    tile[4482] = 6'd37;
    tile[4483] = 6'd37;
    tile[4484] = 6'd37;
    tile[4485] = 6'd37;
    tile[4486] = 6'd37;
    tile[4487] = 6'd37;
    tile[4488] = 6'd37;
    tile[4489] = 6'd37;
    tile[4490] = 6'd37;
    tile[4491] = 6'd37;
    tile[4492] = 6'd37;
    tile[4493] = 6'd37;
    tile[4494] = 6'd37;
    tile[4495] = 6'd37;
    tile[4496] = 6'd37;
    tile[4497] = 6'd37;
    tile[4498] = 6'd37;
    tile[4499] = 6'd37;
    tile[4500] = 6'd37;
    tile[4501] = 6'd37;
    tile[4502] = 6'd37;
    tile[4503] = 6'd37;
    tile[4504] = 6'd37;
    tile[4505] = 6'd37;
    tile[4506] = 6'd37;
    tile[4507] = 6'd37;
    tile[4508] = 6'd37;
    tile[4509] = 6'd37;
    tile[4510] = 6'd37;
    tile[4511] = 6'd37;
    tile[4512] = 6'd37;
    tile[4513] = 6'd37;
    tile[4514] = 6'd37;
    tile[4515] = 6'd37;
    tile[4516] = 6'd37;
    tile[4517] = 6'd37;
    tile[4518] = 6'd37;
    tile[4519] = 6'd37;
    tile[4520] = 6'd37;
    tile[4521] = 6'd37;
    tile[4522] = 6'd37;
    tile[4523] = 6'd37;
    tile[4524] = 6'd37;
    tile[4525] = 6'd37;
    tile[4526] = 6'd37;
    tile[4527] = 6'd37;
    tile[4528] = 6'd37;
    tile[4529] = 6'd37;
    tile[4530] = 6'd37;
    tile[4531] = 6'd37;
    tile[4532] = 6'd37;
    tile[4533] = 6'd37;
    tile[4534] = 6'd37;
    tile[4535] = 6'd37;
    tile[4536] = 6'd37;
    tile[4537] = 6'd37;
    tile[4538] = 6'd37;
    tile[4539] = 6'd37;
    tile[4540] = 6'd37;
    tile[4541] = 6'd37;
    tile[4542] = 6'd37;
    tile[4543] = 6'd37;
    tile[4544] = 6'd37;
    tile[4545] = 6'd37;
    tile[4546] = 6'd37;
    tile[4547] = 6'd37;
    tile[4548] = 6'd37;
    tile[4549] = 6'd37;
    tile[4550] = 6'd37;
    tile[4551] = 6'd37;
    tile[4552] = 6'd37;
    tile[4553] = 6'd37;
    tile[4554] = 6'd37;
    tile[4555] = 6'd37;
    tile[4556] = 6'd37;
    tile[4557] = 6'd37;
    tile[4558] = 6'd37;
    tile[4559] = 6'd37;
    tile[4560] = 6'd37;
    tile[4561] = 6'd37;
    tile[4562] = 6'd37;
    tile[4563] = 6'd37;
    tile[4564] = 6'd37;
    tile[4565] = 6'd37;
    tile[4566] = 6'd37;
    tile[4567] = 6'd37;
    tile[4568] = 6'd37;
    tile[4569] = 6'd37;
    tile[4570] = 6'd37;
    tile[4571] = 6'd37;
    tile[4572] = 6'd37;
    tile[4573] = 6'd37;
    tile[4574] = 6'd37;
    tile[4575] = 6'd37;
    tile[4576] = 6'd37;
    tile[4577] = 6'd37;
    tile[4578] = 6'd37;
    tile[4579] = 6'd37;
    tile[4580] = 6'd37;
    tile[4581] = 6'd37;
    tile[4582] = 6'd37;
    tile[4583] = 6'd37;
    tile[4584] = 6'd37;
    tile[4585] = 6'd37;
    tile[4586] = 6'd37;
    tile[4587] = 6'd37;
    tile[4588] = 6'd37;
    tile[4589] = 6'd37;
    tile[4590] = 6'd37;
    tile[4591] = 6'd37;
    tile[4592] = 6'd37;
    tile[4593] = 6'd37;
    tile[4594] = 6'd37;
    tile[4595] = 6'd37;
    tile[4596] = 6'd37;
    tile[4597] = 6'd37;
    tile[4598] = 6'd37;
    tile[4599] = 6'd37;
    tile[4600] = 6'd37;
    tile[4601] = 6'd37;
    tile[4602] = 6'd37;
    tile[4603] = 6'd37;
    tile[4604] = 6'd37;
    tile[4605] = 6'd37;
    tile[4606] = 6'd37;
    tile[4607] = 6'd37;
    tile[4608] = 6'd37;
    tile[4609] = 6'd37;
    tile[4610] = 6'd37;
    tile[4611] = 6'd37;
    tile[4612] = 6'd37;
    tile[4613] = 6'd37;
    tile[4614] = 6'd37;
    tile[4615] = 6'd37;
    tile[4616] = 6'd37;
    tile[4617] = 6'd37;
    tile[4618] = 6'd37;
    tile[4619] = 6'd37;
    tile[4620] = 6'd37;
    tile[4621] = 6'd37;
    tile[4622] = 6'd37;
    tile[4623] = 6'd37;
    tile[4624] = 6'd37;
    tile[4625] = 6'd37;
    tile[4626] = 6'd37;
    tile[4627] = 6'd37;
    tile[4628] = 6'd37;
    tile[4629] = 6'd37;
    tile[4630] = 6'd37;
    tile[4631] = 6'd37;
    tile[4632] = 6'd37;
    tile[4633] = 6'd37;
    tile[4634] = 6'd37;
    tile[4635] = 6'd37;
    tile[4636] = 6'd37;
    tile[4637] = 6'd37;
    tile[4638] = 6'd37;
    tile[4639] = 6'd37;
    tile[4640] = 6'd37;
    tile[4641] = 6'd37;
    tile[4642] = 6'd37;
    tile[4643] = 6'd37;
    tile[4644] = 6'd37;
    tile[4645] = 6'd37;
    tile[4646] = 6'd37;
    tile[4647] = 6'd37;
    tile[4648] = 6'd37;
    tile[4649] = 6'd37;
    tile[4650] = 6'd37;
    tile[4651] = 6'd37;
    tile[4652] = 6'd37;
    tile[4653] = 6'd37;
    tile[4654] = 6'd37;
    tile[4655] = 6'd37;
    tile[4656] = 6'd37;
    tile[4657] = 6'd37;
    tile[4658] = 6'd37;
    tile[4659] = 6'd37;
    tile[4660] = 6'd37;
    tile[4661] = 6'd37;
    tile[4662] = 6'd37;
    tile[4663] = 6'd37;
    tile[4664] = 6'd37;
    tile[4665] = 6'd37;
    tile[4666] = 6'd37;
    tile[4667] = 6'd37;
    tile[4668] = 6'd37;
    tile[4669] = 6'd37;
    tile[4670] = 6'd37;
    tile[4671] = 6'd37;
    tile[4672] = 6'd37;
    tile[4673] = 6'd37;
    tile[4674] = 6'd37;
    tile[4675] = 6'd37;
    tile[4676] = 6'd37;
    tile[4677] = 6'd37;
    tile[4678] = 6'd37;
    tile[4679] = 6'd37;
    tile[4680] = 6'd37;
    tile[4681] = 6'd37;
    tile[4682] = 6'd37;
    tile[4683] = 6'd37;
    tile[4684] = 6'd37;
    tile[4685] = 6'd37;
    tile[4686] = 6'd37;
    tile[4687] = 6'd37;
    tile[4688] = 6'd37;
    tile[4689] = 6'd37;
    tile[4690] = 6'd37;
    tile[4691] = 6'd37;
    tile[4692] = 6'd37;
    tile[4693] = 6'd37;
    tile[4694] = 6'd37;
    tile[4695] = 6'd37;
    tile[4696] = 6'd37;
    tile[4697] = 6'd37;
    tile[4698] = 6'd37;
    tile[4699] = 6'd37;
    tile[4700] = 6'd37;
    tile[4701] = 6'd37;
    tile[4702] = 6'd37;
    tile[4703] = 6'd37;
    tile[4704] = 6'd37;
    tile[4705] = 6'd37;
    tile[4706] = 6'd37;
    tile[4707] = 6'd37;
    tile[4708] = 6'd37;
    tile[4709] = 6'd37;
    tile[4710] = 6'd37;
    tile[4711] = 6'd37;
    tile[4712] = 6'd37;
    tile[4713] = 6'd37;
    tile[4714] = 6'd37;
    tile[4715] = 6'd37;
    tile[4716] = 6'd37;
    tile[4717] = 6'd37;
    tile[4718] = 6'd37;
    tile[4719] = 6'd37;
    tile[4720] = 6'd37;
    tile[4721] = 6'd37;
    tile[4722] = 6'd37;
    tile[4723] = 6'd37;
    tile[4724] = 6'd37;
    tile[4725] = 6'd37;
    tile[4726] = 6'd37;
    tile[4727] = 6'd37;
    tile[4728] = 6'd37;
    tile[4729] = 6'd37;
    tile[4730] = 6'd37;
    tile[4731] = 6'd37;
    tile[4732] = 6'd37;
    tile[4733] = 6'd37;
    tile[4734] = 6'd37;
    tile[4735] = 6'd37;
    tile[4736] = 6'd37;
    tile[4737] = 6'd37;
    tile[4738] = 6'd37;
    tile[4739] = 6'd37;
    tile[4740] = 6'd37;
    tile[4741] = 6'd37;
    tile[4742] = 6'd37;
    tile[4743] = 6'd37;
    tile[4744] = 6'd37;
    tile[4745] = 6'd37;
    tile[4746] = 6'd37;
    tile[4747] = 6'd37;
    tile[4748] = 6'd37;
    tile[4749] = 6'd37;
    tile[4750] = 6'd37;
    tile[4751] = 6'd37;
    tile[4752] = 6'd37;
    tile[4753] = 6'd37;
    tile[4754] = 6'd37;
    tile[4755] = 6'd37;
    tile[4756] = 6'd37;
    tile[4757] = 6'd37;
    tile[4758] = 6'd37;
    tile[4759] = 6'd37;
    tile[4760] = 6'd37;
    tile[4761] = 6'd37;
    tile[4762] = 6'd37;
    tile[4763] = 6'd37;
    tile[4764] = 6'd37;
    tile[4765] = 6'd37;
    tile[4766] = 6'd37;
    tile[4767] = 6'd37;
    tile[4768] = 6'd37;
    tile[4769] = 6'd37;
    tile[4770] = 6'd37;
    tile[4771] = 6'd37;
    tile[4772] = 6'd37;
    tile[4773] = 6'd37;
    tile[4774] = 6'd37;
    tile[4775] = 6'd37;
    tile[4776] = 6'd37;
    tile[4777] = 6'd37;
    tile[4778] = 6'd37;
    tile[4779] = 6'd37;
    tile[4780] = 6'd37;
    tile[4781] = 6'd37;
    tile[4782] = 6'd37;
    tile[4783] = 6'd37;
    tile[4784] = 6'd37;
    tile[4785] = 6'd37;
    tile[4786] = 6'd37;
    tile[4787] = 6'd37;
    tile[4788] = 6'd37;
    tile[4789] = 6'd37;
    tile[4790] = 6'd37;
    tile[4791] = 6'd37;
    tile[4792] = 6'd37;
    tile[4793] = 6'd37;
    tile[4794] = 6'd37;
    tile[4795] = 6'd37;
    tile[4796] = 6'd37;
    tile[4797] = 6'd37;
    tile[4798] = 6'd37;
    tile[4799] = 6'd37;