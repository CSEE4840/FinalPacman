localparam logic [1:0] GHOST_LEFT [0:15][0:15] = '{
    '{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd1,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd2,2'd1,2'd1,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd1,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd1,2'd0,2'd1,2'd1,2'd0,2'd0,2'd1,2'd1,2'd0,2'd1,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0,2'd1,2'd0,2'd0,2'd0,2'd1,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0},
    '{2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0,2'd0}
};
