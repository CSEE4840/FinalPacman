0000
0000
0000
03e0
0ff8
1ffc
1ffc
3ffe
3ffe
3f7e
3e3e
1e3c
1c1c
0c30
0000
0000
