05FF
0A18
0D97
0FD9
105F
0FC7
0F31
0ED3
0E1F
0D32
0D19
0E32
0F54
0F3F
0E4B
0DC1
0DE8
0DDC
0D5D
0D77
0E93
0EDC
0C03
068B
01DB
0080
0183
0245
0206
022B
0378
04AE
0470
033C
028C
02AC
02B4
0271
02D2
03CC
0340
FF50
F952
F501
F499
F6AD
F846
F83D
F7B2
F7C7
F81E
F7D3
F711
F6DC
F79A
F899
F900
F8B4
F831
F7EE
F818
F8A3
F952
F9BD
F986
F8A5
F78E
F6E4
F6E5
F725
F6F8
F63B
F5A0
F5EC
F6D5
F70D
F5D3
F449
F454
F623
F7B2
F73E
F5A1
F570
F804
FC60
0107
05C5
0AD5
0F18
10BF
0FCF
0E9F
0F09
103A
103A
0EE7
0E06
0E97
0F76
0F38
0E3E
0DE2
0E38
0E1E
0D68
0D5D
0E52
0E30
0AC9
051E
00C1
FFE7
0144
022E
01D1
0158
01AB
0259
02CC
033C
03CD
03D7
02FA
023B
02BE
0398
0245
FDB6
F828
F512
F596
F7AE
F8C4
F84F
F78C
F77A
F7E4
F81E
F7F1
F7A7
F794
F7BD
F7D3
F793
F739
F753
F80D
F8D2
F901
F8CB
F8EF
F97F
F978
F82A
F68D
F642
F753
F800
F72B
F5E1
F5B3
F668
F67B
F5A2
F54A
F649
F748
F6BA
F59D
F69A
FA6F
FEE7
0215
04F3
0965
0E9B
1171
107B
0E04
0D33
0E6D
0FAD
0FBE
0F6D
0F85
0F70
0E9E
0DEF
0E58
0F12
0EA7
0D75
0D6B
0ED5
0EFF
0B47
04D7
FFCE
FEB8
0039
018F
01E7
022A
02A1
028D
01CE
0174
022C
0334
038F
036D
036B
02D4
000D
FB1B
F695
F516
F664
F80C
F871
F831
F87B
F924
F913
F804
F711
F74E
F87A
F951
F8EE
F7A3
F68C
F695
F7C0
F91F
F9A0
F90F
F82E
F7B9
F7A6
F782
F72C
F6E0
F6C2
F6C6
F6F5
F74D
F75A
F671
F4DB
F429
F57A
F798
F801
F633
F4D3
F6B7
FB7C
0036
0332
05AD
0966
0DBB
106A
1095
0FAC
0F2D
0EFC
0E92
0E7A
0F6E
10A7
1090
0F1C
0E13
0E95
0F77
0F0B
0DC2
0D8A
0E9C
0E7D
0B13
0599
015F
0018
0098
0101
00E9
00F8
0167
01CC
01FA
0225
0241
0202
01C0
024E
0367
031C
FFD2
FA97
F67B
F584
F6E9
F87E
F910
F8ED
F8A3
F833
F794
F72F
F75A
F7C4
F7F0
F7EC
F813
F84D
F82E
F7B0
F765
F7B4
F856
F8B3
F892
F826
F79A
F6F1
F64F
F602
F624
F692
F734
F7FA
F864
F7C2
F64A
F552
F5CB
F6E3
F6F8
F603
F610
F8BA
FCEC
003C
022E
04BE
0933
0DDB
0FF8
0F4E
0E46
0EAF
0FC0
0FCF
0EEF
0E9A
0F4F
0FE6
0F88
0EFA
0F3F
0FD1
0F83
0E88
0E54
0F28
0EFF
0BD5
066B
01E0
0078
018A
02D2
02F3
023C
017E
011B
011A
016D
01D1
01ED
01B1
0159
00CE
FF63
FC98
F920
F694
F5F7
F6C6
F7C4
F855
F8B1
F900
F8E1
F80D
F6FD
F69F
F75F
F8A2
F94F
F8E2
F7DC
F748
F7BB
F8CD
F97F
F935
F84B
F79D
F78C
F7B9
F7A5
F741
F6C5
F64F
F5F6
F601
F699
F74A
F748
F674
F5B6
F5E7
F6A5
F6E8
F6C1
F7B0
FAC6
FEFD
0244
03FF
05AF
08C7
0C98
0F11
0F4C
0E77
0E2F
0EA9
0F06
0EDC
0EAE
0EE2
0F21
0F03
0ECD
0F08
0F94
0FBE
0F42
0EB2
0E75
0DCC
0B73
074F
02FD
0080
0070
01A8
0299
02B1
0270
0268
027C
023B
01B8
01A5
0268
033A
0281
FF54
FAA0
F696
F4D9
F542
F671
F74E
F7CA
F847
F8BD
F8B2
F7FC
F727
F6F1
F776
F81A
F847
F812
F7FE
F831
F830
F791
F6C7
F6D6
F807
F942
F923
F7B6
F686
F6C5
F7CD
F80C
F722
F661
F6E1
F7DE
F7D6
F6CF
F667
F75F
F837
F74D
F5C3
F6C4
FB91
016C
048E
04A0
04F2
081F
0CD5
0FC3
0FC7
0ED8
0EF5
0FB3
0F89
0E68
0DC9
0E68
0F36
0F14
0E75
0E80
0F2F
0F64
0ED0
0E8F
0F5D
1005
0E88
0A9D
062A
0323
01BE
0127
010D
01AD
02AD
030F
027C
01D7
0200
029D
02C8
0291
02BF
0301
0186
FD3E
F7E4
F4AE
F4F0
F6EA
F835
F86B
F8C2
F9A9
FA0F
F93C
F82D
F854
F984
FA21
F95D
F845
F846
F945
F9D5
F913
F7A9
F6D0
F6FF
F7BC
F862
F894
F83D
F790
F70A
F702
F73E
F73C
F6F2
F6E8
F766
F7E1
F7B5
F717
F6CA
F6E5
F6BB
F653
F728
FA8E
FF8B
0362
04A2
04E1
06B9
0A74
0DBE
0EA7
0DF0
0DB3
0E88
0F1D
0E72
0D61
0D52
0E47
0EF9
0EC5
0E6E
0ECE
0F83
0F9A
0F16
0EE0
0F2D
0EBE
0C48
083B
0492
02D9
02DC
0349
0335
02B3
0244
0234
0283
02F9
032F
02DE
024E
022C
028A
023D
FFC6
FB2C
F687
F449
F502
F717
F89B
F901
F8F5
F909
F924
F914
F90D
F94B
F996
F980
F90C
F8B3
F8C1
F8F3
F8D8
F864
F7ED
F7C2
F801
F8A0
F94F
F964
F85B
F69F
F572
F5AA
F6BF
F770
F73A
F6BA
F691
F693
F665
F654
F6CC
F745
F6C0
F5BD
F68C
FAB2
0074
0444
04D6
04B6
0708
0B8F
0F14
0F83
0E2B
0D75
0DC1
0DC1
0D21
0D27
0E7D
0FCD
0F97
0E7E
0E61
0F7E
0FF9
0EB2
0D2E
0D7F
0F0C
0EF1
0BAA
0703
03D7
02E1
02BA
026C
028A
0399
04AB
0480
0347
0243
0204
020D
0224
02BF
039B
02E6
FF0E
F935
F4C2
F3FD
F5E9
F7EA
F8CD
F946
F9FF
FA6B
F9E2
F8E6
F87A
F8AB
F89E
F806
F7A5
F813
F8B8
F8A3
F7F0
F79C
F826
F8FA
F96C
F978
F94F
F8A9
F743
F5C4
F550
F60F
F6D7
F6B6
F62F
F653
F71D
F781
F720
F6CF
F719
F72D
F64D
F5CE
F820
FD73
0290
0444
035A
03D0
07E6
0D49
0FF2
0EEB
0CF8
0CC6
0DF6
0E88
0DF3
0D85
0E1E
0F05
0F4F
0F40
0F76
0F6A
0E25
0C40
0BDA
0DCF
0FE4
0EE7
0A68
055C
02DD
031C
03FA
03EF
034D
0306
0335
0363
035A
0320
0286
0195
011B
01DC
02FC
0215
FDC9
F7E4
F413
F444
F6E5
F8F5
F91C
F858
F80A
F86B
F8DB
F8F0
F8B7
F853
F7EC
F7DE
F86A
F92A
F95F
F8E7
F877
F89A
F8EB
F8C5
F859
F85D
F8BF
F86E
F6DA
F512
F4A5
F5B5
F6D8
F70B
F6D0
F70B
F789
F786
F726
F74E
F7F5
F7D6
F693
F63A
F937
FEE4
038D
04A9
03FB
0557
09CF
0E77
102D
0F3A
0E3E
0E8A
0EF8
0E5A
0D68
0D65
0E04
0DE8
0CF5
0CA6
0DBF
0EE5
0E77
0D11
0CDA
0E54
0F2B
0CF8
0867
048A
0354
03C1
03B2
0296
0195
01A9
0279
0319
031C
02A5
0213
01F8
02D4
041E
03EE
0095
FAD3
F5CF
F434
F5AD
F79D
F824
F7AE
F794
F824
F8A2
F8A8
F899
F8D0
F918
F937
F96B
F9E7
FA32
F9A5
F872
F796
F79C
F80D
F847
F856
F878
F849
F737
F5B4
F515
F5F1
F734
F77D
F6E6
F6A4
F71C
F75D
F6CB
F642
F6A9
F739
F68E
F550
F64B
FAF5
00E1
0424
0413
041B
0762
0CBC
1032
0FE1
0DD0
0CF4
0DC0
0E88
0E45
0D9C
0D56
0D34
0CD7
0CC0
0D7A
0E57
0E2B
0D43
0D5F
0F3F
1103
0FE4
0B76
0647
0329
0291
02F0
02ED
0281
0232
022D
0259
029F
02D0
02A1
0241
028D
03F6
052D
03C5
FECC
F858
F3F5
F36C
F585
F7C2
F8C4
F8D4
F8C3
F8F5
F957
F9AD
F9A3
F90E
F869
F89D
F9DA
FAFF
FAAE
F8FB
F77D
F765
F826
F861
F7D4
F782
F7FA
F860
F7A5
F629
F552
F5B9
F689
F6E0
F6ED
F73A
F772
F6D9
F5C3
F576
F642
F6C6
F604
F586
F7F6
FD72
029A
044C
0388
0447
0879
0DA5
100C
0F1C
0D73
0D27
0DA6
0D87
0D00
0D41
0E31
0E4E
0D14
0C09
0CA3
0E11
0E63
0D7D
0D65
0F35
10F5
0F99
0AC0
055D
0280
025D
02F2
02C8
0220
01DE
0231
02AF
02FE
02FF
02B7
0277
02CB
039F
0391
00F0
FBC2
F66D
F3A6
F3FF
F5C7
F720
F7A6
F803
F8A8
F95C
F9CA
F9D8
F987
F8F2
F88E
F8E5
F9D5
FA72
FA12
F924
F897
F894
F87C
F816
F807
F8B8
F953
F8AD
F6F8
F5C4
F5FC
F6C5
F6E1
F67A
F6AE
F792
F7E4
F6FD
F609
F65F
F75A
F731
F5F7
F64F
FA2F
FFD8
0380
03D7
0391
05E3
0A8F
0E73
0F7B
0EA6
0E06
0E17
0DF8
0D61
0D10
0D4C
0D54
0CB6
0C4B
0D09
0E49
0E6D
0D3D
0C87
0DBB
0F9B
0F5A
0BE3
071F
03C3
029C
0276
0217
017D
013C
0185
0225
02E5
0372
034D
0276
01E7
0291
03B9
0311
FF1E
F945
F4CD
F3C9
F566
F756
F834
F83F
F83D
F881
F8FC
F980
F9BA
F954
F886
F82B
F8C2
F991
F967
F841
F781
F820
F955
F9A3
F8E8
F86B
F8E0
F94A
F86F
F6C6
F5EE
F670
F71B
F6E5
F670
F6DC
F7D3
F7EE
F6F9
F670
F747
F832
F782
F627
F734
FBE6
0175
0428
03DD
0420
078D
0C9A
0FB4
0FA4
0E6A
0E1B
0E6E
0E09
0CF7
0C92
0D52
0E20
0E0A
0D99
0DC0
0E33
0DE3
0CE9
0CC5
0E2D
0F84
0E60
0A5B
058E
024B
0115
0100
014F
01EE
02BC
0338
031F
02BE
0267
0202
0196
01B5
029F
0330
017D
FD06
F7C6
F490
F466
F5F6
F775
F859
F902
F989
F998
F92B
F8B9
F87D
F837
F7CD
F7BB
F864
F944
F96D
F8C4
F82E
F84F
F8B7
F8B1
F85B
F84C
F863
F7D5
F684
F580
F5AC
F66A
F674
F5CD
F5C7
F6EF
F7FB
F799
F67E
F678
F7A1
F7FE
F68C
F579
F7D7
FD6F
0281
0445
0448
062B
0AC3
0F1E
106B
0F59
0E9D
0F31
0FA1
0ECC
0DB1
0DB0
0E45
0DE1
0C8A
0C20
0DB2
0FC0
1019
0EBF
0DB6
0E0B
0E33
0C1A
07E5
03DD
01CC
016B
016B
0131
00FE
0111
0154
01CF
02A9
0391
03C1
02FE
020E
01A8
0124
FF0A
FB1E
F732
F572
F625
F798
F827
F7D4
F7AD
F83F
F90E
F96F
F94C
F901
F8DA
F8E4
F90D
F92C
F915
F8CE
F8A2
F8C8
F902
F8DC
F857
F7FA
F807
F807
F76B
F674
F5FB
F64C
F6BA
F6A1
F65D
F6AF
F76F
F78C
F69C
F59C
F5A8
F667
F69D
F63C
F6E0
F9C3
FDD4
00E3
026A
042F
07C4
0C36
0F26
0FB3
0F48
0F79
100B
0FC4
0E82
0D7D
0D80
0DD8
0D8A
0CD9
0CD6
0DBA
0E9D
0EE7
0F32
101A
10B5
0F30
0B09
0610
02AF
0194
0184
012D
007E
002D
0077
00E9
0114
0113
014E
020A
0343
0474
0477
0216
FD52
F80A
F4CB
F4A7
F66B
F81A
F8D9
F928
F989
F9B6
F949
F895
F84F
F8A3
F915
F950
F990
F9FF
FA2B
F988
F857
F795
F7E2
F8D2
F980
F973
F8C2
F7A4
F657
F548
F4E4
F516
F558
F572
F5D6
F6E0
F80B
F868
F7DE
F756
F75C
F736
F620
F50A
F626
FA40
FF40
0233
02A3
0312
05DE
0A6C
0E12
0F55
0F49
0F9B
1046
1001
0E7D
0D0E
0CE9
0D9B
0DDD
0D78
0D6C
0E41
0F1A
0EF7
0E4F
0E82
0FD2
10B5
0F7A
0C1B
0809
049A
0238
00E9
00BE
0173
022C
022A
01A3
015F
01A2
01E8
01E2
020D
02C8
032B
018E
FD72
F86B
F4D8
F3DA
F4B8
F619
F759
F88C
F9A6
FA19
F982
F855
F79D
F800
F917
F9DE
F9BB
F905
F878
F858
F858
F845
F866
F8FD
F9B0
F9CB
F909
F7DF
F6DF
F622
F571
F4D7
F4B2
F529
F5E3
F66B
F6A6
F6B7
F6A3
F65A
F601
F5E5
F613
F650
F6A2
F7A3
FA0E
FDBB
0166
03AE
0470
04FE
06DA
0A33
0DB2
0FBD
0FEA
0F34
0EC2
0EC6
0EA1
0E0C
0D8E
0DC2
0E79
0EF7
0EEC
0EBE
0EC8
0EC7
0E56
0DC0
0DC3
0E59
0E40
0C31
086F
04BD
02B4
0263
029E
0271
01F0
01BB
021C
02B9
0309
02DB
0264
01F4
0195
00D4
FEFA
FBB9
F7D0
F4D0
F3EC
F4E7
F65E
F727
F748
F776
F7F1
F843
F819
F7E4
F83A
F8EA
F920
F88E
F7EA
F801
F8AE
F914
F8C6
F841
F835
F8AA
F90C
F8DF
F824
F72A
F64B
F5CC
F5BE
F5D3
F5AB
F55B
F55F
F5E1
F64D
F612
F585
F58B
F64C
F6D7
F67C
F628
F7C0
FBE5
00CB
03D6
0448
03E9
0510
0845
0C11
0EB3
0FC1
0FFA
1004
0FBC
0EEA
0E15
0E0F
0EDC
0F81
0F3F
0E84
0E4B
0EB2
0ED0
0E10
0D2F
0D60
0E9A
0F5C
0E39
0B26
073A
03A6
0148
00A9
019F
0317
03D3
0395
032E
0336
033A
0292
01A8
018D
022F
01D9
FF0B
FA66
F628
F3EA
F383
F403
F504
F68B
F834
F924
F8F5
F831
F7A0
F76B
F740
F713
F743
F7F1
F89F
F8C2
F875
F85A
F8BF
F92A
F8F5
F838
F7CE
F83B
F8E4
F8B0
F75E
F5DD
F52C
F552
F5A8
F5E2
F63D
F6BA
F6BD
F5F1
F513
F531
F620
F681
F5B6
F554
F7B6
FD20
02E1
05C5
0541
03E6
04BC
0869
0CE7
0FC2
1042
0F83
0EDB
0EA0
0E67
0E0C
0E05
0EAB
0F8E
0FD8
0F5E
0ECE
0EC1
0EF7
0ED1
0E50
0E18
0E73
0E94
0D2B
09BD
055C
01F7
00DA
01C3
033C
03F8
03D1
038A
039A
037C
0290
0161
0156
02BB
03AD
01BE
FCBB
F73D
F437
F43C
F582
F64A
F693
F755
F8A9
F973
F8DA
F778
F6B8
F736
F838
F8A9
F85D
F808
F82B
F86F
F850
F7FA
F811
F8A2
F8FA
F897
F7EA
F7AE
F7D8
F7AD
F6E4
F61F
F601
F63C
F60E
F57B
F546
F5B3
F605
F5A7
F52F
F576
F62B
F627
F575
F600
F98D
FF3C
03DB
050A
03A3
02B5
0463
082D
0C07
0E73
0F5A
0F5F
0EFE
0E66
0DE0
0DDE
0E81
0F49
0F95
0F58
0F1F
0F3C
0F4D
0EC3
0DB5
0CF2
0D1F
0E02
0E8D
0DA5
0ADF
06E5
0346
019B
0235
03A3
040C
0319
0220
022E
02B6
029C
0207
021D
02EB
02A1
FF98
FAB3
F6C7
F5A0
F659
F6F5
F6D4
F6D1
F783
F84B
F852
F7B2
F741
F785
F837
F8C4
F8F3
F8E9
F8C1
F86D
F805
F7F5
F88D
F97F
F9F8
F96B
F848
F7A5
F801
F885
F7FB
F663
F511
F50D
F5E8
F688
F697
F696
F6BD
F69E
F607
F597
F5D1
F61D
F59C
F4F9
F66B
FB1D
012C
0511
0518
0301
021A
0430
0863
0C72
0EBF
0F33
0EB5
0E26
0DDB
0DC4
0DD7
0E29
0EA5
0EDC
0E6C
0DA2
0D4F
0DCA
0E63
0E3B
0D77
0D22
0DCC
0E86
0DA6
0A8B
067B
038D
02BA
0324
034E
02C5
023E
0249
025D
01B0
00B6
00F5
02E4
0481
02F5
FDD8
F81A
F51E
F55F
F686
F680
F5AB
F5B4
F725
F8C9
F94E
F8D4
F863
F878
F896
F848
F7E5
F80F
F8C8
F96D
F98F
F97D
F9C2
FA3D
FA2A
F920
F7CD
F749
F7C3
F854
F81E
F739
F64B
F5B5
F573
F595
F63D
F71E
F77B
F70E
F67F
F681
F6A5
F5EC
F49C
F4B7
F7F3
FD82
0291
04DC
0470
0336
033A
056B
0940
0D18
0F32
0EFA
0D8B
0C9B
0CD0
0D6A
0DA4
0DB4
0E23
0EAE
0E95
0DCF
0D37
0D66
0DE7
0DE3
0D61
0D57
0E4B
0F2E
0E14
0A39
052B
01A6
0123
0296
03A4
031F
01FF
01C3
0268
02C0
0279
029C
037F
035B
0022
FA7E
F5C9
F48A
F5C5
F68A
F59C
F491
F541
F74F
F8E2
F911
F8A2
F89C
F915
F982
F990
F953
F8EE
F877
F826
F854
F91E
FA19
FA93
FA29
F91E
F82B
F7E6
F83C
F87B
F803
F6FD
F639
F636
F6A9
F6FF
F709
F6F3
F6D6
F6B4
F699
F67F
F627
F58A
F576
F73B
FB5A
0081
0459
057B
0485
034C
0369
0574
08F4
0C97
0ED9
0F20
0E4A
0DB3
0DCE
0DF9
0DA2
0D1E
0D13
0D75
0DA5
0D81
0DAD
0E82
0F40
0EEA
0DBF
0D1F
0DBE
0E69
0D26
0970
0507
023A
0194
01AF
013D
00AC
0139
02CF
03D7
0361
028F
02F2
03E5
02AC
FDD0
F788
F3C2
F3F3
F5D3
F67D
F5AD
F53C
F63A
F7C0
F88A
F8A6
F8F2
F99A
F9E1
F949
F861
F818
F8A5
F973
F9E3
F9DC
F9A1
F972
F955
F915
F878
F7A7
F72D
F768
F7F8
F802
F721
F5E8
F565
F60C
F731
F7A5
F6FC
F5FE
F5BA
F63E
F680
F5BD
F4BF
F561
F89E
FD5E
0175
0399
0405
038E
02F1
0327
054D
0961
0D78
0F3D
0E61
0CDD
0CA4
0D91
0E25
0DC9
0D59
0D8C
0DCE
0D60
0CDA
0D81
0F4D
1095
100E
0E7F
0DE5
0EF2
0FE4
0E46
09B6
049B
01CF
01E4
02F6
031B
0254
01F0
0277
0318
031A
0306
0375
0351
0094
FB39
F62B
F463
F5AA
F718
F6A4
F524
F4B0
F5F9
F7D6
F8FF
F94A
F930
F8F7
F8B7
F8AD
F8F3
F92F
F917
F8F4
F937
F9C7
FA17
F9D7
F92B
F851
F780
F713
F766
F846
F8D1
F84C
F706
F60A
F5E1
F617
F615
F5F3
F61A
F684
F6C1
F681
F5CD
F505
F507
F6DF
FAC5
FF64
02B2
03B2
0328
0288
02A5
03AD
05DD
093D
0CAE
0E70
0E20
0D5B
0DC1
0ED8
0EF8
0DCC
0CDF
0D64
0E8D
0EBE
0DDD
0D54
0DE8
0EB7
0EBF
0E82
0F0F
0FEC
0F20
0BB1
0729
0418
0364
03AD
0353
025E
0211
02EA
03DE
03B3
02A5
01F8
0219
01B6
FF31
FABC
F688
F4A8
F50A
F5D9
F5B1
F4F0
F4CF
F5AE
F6CB
F765
F7A0
F819
F8E4
F95F
F902
F826
F7C0
F856
F962
F9D3
F934
F823
F7A5
F817
F8E0
F91D
F892
F7E7
F7ED
F8B9
F979
F942
F800
F688
F5B3
F57F
F541
F4C3
F4AD
F577
F64D
F5F8
F4E5
F550
F8BF
FDF0
020F
03C6
041D
0461
044A
0339
0264
0423
08CD
0DA2
0FC1
0F4A
0E9A
0F19
0FF0
0FCE
0EBB
0DBB
0D6D
0DB4
0E54
0F2B
0FC1
0F66
0E13
0CB9
0C50
0CFB
0E3B
0F48
0F06
0C6F
07F4
03D3
022E
02D3
0399
02F2
017C
00DB
01AC
0325
0431
03FE
01CD
FD72
F876
F577
F579
F6AA
F6A5
F549
F44E
F48D
F516
F501
F4E9
F5C4
F724
F7BD
F779
F7AF
F8FC
FA16
F9A5
F845
F7A3
F81B
F87A
F7E7
F701
F6CF
F766
F819
F88E
F8FD
F981
F9B4
F94A
F880
F7B9
F70E
F67D
F627
F60C
F5ED
F5C0
F5D2
F614
F5DA
F500
F4F9
F7AC
FCF4
0208
0428
0382
02B2
035B
0470
043E
0341
03C5
06FC
0B79
0EC4
0FD5
0F81
0F07
0EDA
0EBD
0E7F
0E37
0E13
0E3B
0EBE
0F64
0FB6
0F74
0EE7
0E79
0E20
0D8A
0CE5
0CEC
0DBB
0E03
0C20
082B
0448
0293
02F7
0394
0306
01BC
010D
018F
02AB
0358
02B0
0022
FBF1
F7AB
F558
F58C
F6BA
F6F2
F5E6
F4CD
F484
F4B7
F4D6
F518
F5F2
F70E
F7A0
F7A0
F7E6
F8C7
F982
F964
F8D2
F881
F84F
F7B2
F6E7
F6D0
F7A4
F886
F8B7
F88E
F8CE
F95C
F96C
F8C8
F805
F765
F67A
F543
F4AC
F54A
F65F
F6E8
F6F8
F725
F726
F664
F5D8
F7E4
FD3F
02FF
053C
0399
01A2
0240
044B
04CF
0376
02FB
058C
0A2C
0E11
0F96
0F47
0EAC
0EA5
0EFB
0EF5
0E37
0D48
0D3E
0E75
0FBA
0F7E
0DEC
0CDB
0D4C
0E14
0DC8
0D0E
0DA2
0F6D
1003
0D82
0900
0544
03AD
0348
02BF
01F2
0156
0106
011D
0213
038E
038F
003C
FA8A
F5F7
F500
F694
F79F
F69F
F4DE
F431
F4B9
F556
F58F
F601
F710
F829
F88E
F851
F82A
F898
F962
F9ED
F9D4
F928
F856
F7D0
F7C5
F807
F846
F865
F892
F8F6
F967
F985
F918
F834
F71C
F630
F5D9
F64F
F746
F802
F7ED
F71A
F60A
F518
F466
F47A
F669
FAC8
005B
047D
055C
03CF
026B
02C1
03F4
0432
0329
0282
040F
07E5
0C30
0EC4
0ED7
0D85
0CD0
0DD2
0FB6
1097
0F9B
0DFE
0D84
0E38
0E85
0D93
0C82
0CB4
0DBA
0E0A
0D6A
0D5A
0EC0
100A
0EB3
0A58
0561
0274
01FA
0274
0275
01B3
00D0
00BC
01D5
0303
0227
FE32
F8CD
F519
F4A1
F600
F6CD
F636
F531
F49A
F451
F442
F4FD
F69E
F80E
F847
F7C6
F7D1
F8A6
F953
F93C
F8EB
F908
F959
F941
F8DE
F8DF
F959
F9A3
F96F
F935
F931
F8F4
F86A
F86A
F95F
FA1B
F928
F6F7
F590
F5EC
F6C6
F6A5
F614
F6A1
F80B
F83F
F6A5
F5E9
F904
FF26
0421
0508
0329
01FD
0315
04D7
0501
0385
028C
0417
0809
0C64
0F10
0F75
0E9C
0DF6
0DFD
0E16
0DC4
0D70
0DCD
0EC4
0F74
0F38
0E56
0D8C
0D3B
0D38
0D46
0D7B
0E09
0EB8
0EBC
0D19
097E
04F4
019F
0126
02FA
0492
03DA
016B
FFE2
00BC
0263
01C1
FDB0
F843
F49D
F3EA
F4CC
F571
F566
F554
F58D
F5A0
F537
F4BF
F4F7
F605
F75B
F84F
F89B
F86E
F83D
F870
F909
F985
F957
F898
F80D
F859
F941
FA02
FA41
FA2B
F9D9
F922
F83A
F7DF
F865
F90F
F8DA
F7C7
F6C4
F664
F64A
F61D
F64C
F734
F807
F7A2
F697
F73B
FAE4
FFE8
033B
03B2
02DB
02C6
03D2
04D5
04C4
03C9
0317
0425
07AD
0CB6
10B3
1183
0FAD
0DD7
0DB8
0E65
0E35
0D4E
0D41
0E89
0FD1
0FE4
0F48
0F26
0F5C
0EBF
0D2B
0C1F
0CC1
0E35
0E85
0CB7
0955
0584
0267
00F6
015E
0270
0294
01A7
0139
025B
039E
023C
FD66
F790
F3EF
F356
F415
F47A
F462
F480
F4FE
F56C
F584
F58D
F5DD
F65C
F6AF
F6BE
F6E1
F776
F868
F92F
F94E
F8D9
F86C
F88B
F903
F934
F8E1
F88B
F8B6
F92F
F95C
F91E
F907
F985
FA2F
FA21
F8FD
F758
F61D
F5BE
F60C
F6A6
F73F
F776
F6E7
F5C2
F53A
F6D8
FB0E
0060
0455
056E
0458
031C
032D
0438
04D0
040C
02A2
027E
052F
0A51
0F70
11F7
1178
0FE7
0F5B
0FEB
101D
0F1E
0DE6
0DCD
0EB0
0F2B
0E96
0DE0
0E21
0F09
0F59
0E8F
0D7F
0D3A
0DB8
0DAC
0B9F
0774
02F4
0088
00EC
024E
0236
0087
FFBD
0191
03FF
030E
FD9F
F725
F3C9
F40E
F53C
F54C
F4CC
F4F1
F57A
F55F
F4C0
F4CC
F5EE
F734
F7CA
F7EC
F7F7
F78B
F689
F5FD
F6F9
F8CC
F9A5
F8E3
F7DA
F7EE
F8C9
F921
F8B0
F862
F8AE
F8EF
F8A6
F86E
F8E3
F972
F929
F822
F743
F6DF
F692
F65D
F6D3
F7C4
F7C5
F627
F4D0
F6B8
FC35
01F8
048C
03E9
02C7
0318
0461
0548
0552
04C8
03F7
0383
04C0
087B
0D52
1081
10CB
0FC5
0F97
1046
1049
0F26
0E39
0E96
0F74
0F64
0E70
0DF3
0E77
0EE8
0E3C
0D06
0CAD
0D91
0E9E
0E6A
0C39
084E
03F7
0114
00B2
01D6
025B
0184
00F1
021F
0388
01D5
FC45
F64C
F3D1
F4D2
F611
F579
F42B
F40C
F4ED
F53A
F49A
F464
F574
F6F5
F7C7
F7FE
F834
F847
F7D4
F74C
F77A
F837
F88E
F82E
F7D7
F827
F8B3
F8D6
F8D0
F93D
F9CB
F98D
F8AD
F87B
F95C
F9F6
F920
F79A
F6C2
F67E
F5DC
F531
F5E5
F7E2
F8D6
F74F
F581
F724
FC9E
0228
045C
03D3
0343
03A4
03F1
03B1
039A
03D1
037A
02BB
03A5
07B0
0D05
1006
0F83
0DE5
0DA9
0E5F
0E4C
0D82
0D9E
0F03
1030
0FDF
0E9B
0DB1
0D8D
0DB4
0DCA
0DD3
0DBF
0D86
0D96
0E11
0DA4
0AA0
05BF
024A
0248
03CA
0393
01AB
0133
0371
0517
0219
FB1C
F51E
F3A9
F552
F695
F64E
F5D2
F5EC
F5DD
F53C
F4EE
F59E
F68F
F6CD
F6CB
F79C
F8F5
F953
F853
F78E
F84F
F995
F983
F818
F725
F7AB
F899
F896
F7EF
F7F4
F8F9
F9FC
FA31
F9DC
F964
F899
F76B
F686
F666
F66F
F5EB
F582
F66E
F843
F8D3
F728
F5A0
F7A2
FD4D
02DC
04D7
03B3
0277
02C7
03A9
03B4
02F3
0250
0247
0302
04FF
0887
0C7D
0EE4
0EF0
0DD8
0D27
0D05
0CBF
0C53
0C70
0D3B
0E05
0E65
0EC9
0F91
1030
0FB5
0E18
0C61
0BA0
0C1A
0D6D
0EA5
0E30
0AEA
05DA
0204
017E
0324
0424
0385
02E3
0370
038B
00AC
FB1C
F63E
F4B8
F59B
F61D
F53E
F463
F4DC
F624
F6DB
F693
F610
F627
F6EC
F7DA
F866
F857
F7EF
F7C3
F830
F8CE
F8E8
F884
F867
F8DD
F924
F890
F7B7
F7BF
F8B7
F989
F98D
F96D
F9F7
FAB5
FA7B
F924
F7C8
F721
F6C4
F655
F66B
F762
F810
F712
F549
F5A4
F9BF
FF95
0381
0429
034F
0302
0354
0370
0377
0409
049A
03E6
023F
0203
04FF
09F5
0DCE
0EE9
0E5A
0DE0
0DD7
0DBA
0D97
0DE8
0E67
0E2B
0D0F
0C1B
0C3F
0D39
0E13
0E5D
0E46
0DF0
0D69
0D2F
0DB8
0E31
0CD0
0915
04EA
029C
024B
025D
0229
02B0
0421
0428
0059
F9E1
F506
F470
F659
F73F
F62A
F4E4
F4C4
F512
F4D2
F483
F51B
F62F
F683
F624
F698
F879
FA2F
F9E4
F802
F69F
F6E0
F7FE
F8CA
F91C
F969
F9B3
F998
F923
F8E2
F919
F970
F993
F9AF
F9FA
FA46
FA5A
FA63
FA6E
F9F5
F883
F6B7
F5DE
F65D
F70F
F6A2
F573
F57B
F840
FD06
0169
0387
037B
02D0
02D5
0380
03D7
034C
027F
0269
02FA
032E
02AA
029D
047B
0823
0BD5
0E0C
0EC9
0EDF
0E9D
0DC8
0CB1
0C44
0CE1
0DCF
0E40
0E40
0E33
0DF8
0D4F
0CAE
0CD4
0D92
0DD0
0D34
0CDA
0D9D
0E32
0C41
0794
02F5
0132
0221
0373
03CA
03A0
0336
014D
FCC7
F6E9
F2B1
F1E3
F37E
F55D
F677
F703
F730
F6BE
F5B9
F4BA
F441
F44B
F4C0
F5CF
F777
F90E
F9C0
F979
F8EE
F8AE
F896
F86E
F88C
F95C
FA94
FB63
FB5E
FAD0
FA26
F980
F906
F921
F9F3
FAD6
FAF6
FA7A
FA60
FAEA
FAD3
F8DA
F5DD
F459
F57F
F781
F7B5
F61F
F5D1
F950
FF4F
03E9
04E5
03BD
0321
038E
0367
020E
0128
0242
043E
047D
0284
0116
0302
07B7
0BF5
0DA2
0D94
0D9B
0E03
0DFB
0D78
0D62
0DFA
0E44
0D8A
0C92
0C98
0D88
0E38
0E29
0E0B
0E47
0E32
0D54
0C97
0D0A
0DEF
0D2D
09EF
05D9
031E
0233
0216
023B
02DC
0367
0214
FE01
F8D3
F53C
F432
F489
F4E8
F525
F57D
F59C
F52B
F4B8
F518
F5FB
F623
F54B
F4DB
F610
F820
F92C
F8A8
F7E7
F837
F956
FA09
F9BB
F8FB
F897
F8DB
F999
FA72
FAE3
FA86
F9AB
F944
F9D5
FAAD
FAC1
F9F8
F925
F8CB
F877
F795
F686
F65E
F776
F89A
F820
F5F3
F446
F5D4
FB24
0196
057F
0582
03AA
02E1
03AA
0424
031B
01D2
0210
0368
03CD
02BA
026E
0533
0A28
0DFB
0EA2
0D5A
0CA3
0D60
0E9F
0F4E
0F35
0E90
0DA1
0CCF
0C81
0CB4
0D0F
0D79
0E21
0EBF
0E7F
0D51
0CB1
0DEB
0FB3
0EF7
0AAC
0587
02D9
02B3
029E
019A
015E
0301
0430
01A2
FBB3
F68F
F541
F653
F65E
F4A1
F341
F3B9
F4F4
F559
F522
F58A
F697
F707
F670
F628
F76C
F984
FA9C
FA02
F8B8
F7F0
F7DC
F80D
F84D
F8B0
F928
F974
F97D
F97D
F9BF
FA46
FACD
FB02
FAB8
F9F4
F8FF
F849
F801
F7EA
F7AB
F736
F6CD
F6B9
F6FE
F73F
F704
F682
F708
F9FF
FF17
03D6
05B0
0492
02DB
02A2
0394
0405
0376
0309
036E
03CD
0357
0303
048F
081B
0BC7
0DD6
0E53
0E61
0E8D
0E84
0E12
0D87
0D1B
0CB4
0C7C
0CE8
0DD2
0E53
0E07
0DB8
0E10
0E49
0D47
0BBB
0BB2
0D96
0EBE
0C5B
073B
031B
0220
02A4
0240
015F
020B
03E4
038F
FEDA
F800
F385
F35E
F560
F666
F5B6
F4C5
F4AC
F510
F545
F55F
F5D1
F6B5
F7B9
F880
F8C8
F87C
F7D4
F75E
F79E
F890
F993
F9F8
F9B5
F963
F98F
FA14
FA30
F951
F7DF
F725
F815
FA14
FB6E
FB14
F9A4
F87C
F837
F84E
F7FD
F723
F64D
F627
F6C9
F777
F71A
F59C
F4C4
F710
FCD3
02F3
05B0
04AD
030C
033F
043C
03C7
023F
0234
0457
05F7
04AC
022C
0289
06EE
0C22
0EB3
0EBF
0E85
0EC8
0E7C
0D58
0CA0
0D10
0DAB
0D6D
0D15
0DF2
0F87
0FFE
0EE2
0DCA
0DC8
0DC9
0CA5
0B77
0C0C
0DAE
0D71
0A0C
05B6
0360
032B
0311
024F
0234
032D
0300
FF71
F9A4
F537
F42B
F524
F5C2
F566
F508
F54D
F5D5
F62A
F66C
F6B1
F68C
F5C5
F512
F57B
F71C
F902
FA28
FA33
F973
F8AE
F8B4
F9AC
FAB1
FA91
F917
F773
F70A
F807
F94B
F9CB
F994
F94D
F93A
F91C
F8D5
F8AE
F8D5
F8E8
F824
F63E
F424
F389
F517
F738
F78C
F602
F5B1
F992
007D
05B0
05EC
0320
01C3
033A
04B4
03C3
01F2
0247
04A0
05DB
0484
033D
055A
0A63
0E94
0F6D
0E0D
0CE3
0CB5
0CE6
0D4E
0E39
0F2F
0F45
0E93
0E4A
0EEA
0F82
0F20
0E41
0DDA
0DAC
0CE1
0C13
0CF9
0F5D
101E
0CB4
06D7
02E5
02C8
0424
0403
02AB
0256
0314
021B
FDA8
F7D3
F456
F447
F585
F5D9
F542
F4EB
F52F
F585
F5A2
F5BB
F5C8
F57D
F522
F5AB
F765
F929
F999
F8EC
F89F
F966
FA36
F9C3
F84E
F753
F7A6
F880
F8AE
F81C
F7CB
F869
F98D
FA5B
FA70
F9F3
F928
F843
F799
F769
F773
F70C
F5F3
F4F1
F514
F63C
F6F8
F65F
F5BC
F78B
FC81
0235
0553
04F9
034B
02B4
0362
03F2
03CD
03BE
042E
0428
02E9
01AE
02D4
06FE
0C0A
0F2A
0F91
0E99
0DC4
0D74
0D6B
0D9D
0E05
0E52
0E56
0E61
0EB8
0EEF
0E75
0D8D
0D1F
0D6D
0DBD
0DA1
0DD4
0EEA
0F9D
0DBD
092B
049F
02A4
02CE
02FB
029E
031D
04AE
04AC
007D
F97C
F43B
F393
F5B6
F6EA
F5E7
F470
F43A
F4F4
F574
F58F
F5EA
F6A5
F72E
F74E
F787
F82F
F8CE
F8D8
F88B
F883
F8C0
F8C4
F881
F88D
F940
FA1E
FA59
F9C1
F8F4
F8AB
F8FD
F95E
F944
F8B5
F843
F879
F948
F9EA
F990
F83C
F6D2
F630
F662
F6C0
F68C
F5AA
F50D
F65C
FA81
0027
0452
0516
0396
02A6
038D
04D4
04BC
03C9
03BD
0499
0472
02B2
01BF
0422
08FE
0CEF
0E12
0DB6
0DE1
0EA2
0ED5
0E74
0E83
0EFC
0E91
0D00
0C05
0CEF
0E91
0EE2
0DDD
0D39
0DB5
0E3D
0DFD
0DA8
0DCD
0D17
09F3
057E
02D5
0319
03FA
032E
01A8
0195
0264
011A
FCA0
F7A5
F554
F581
F591
F465
F38E
F479
F621
F6A0
F5D2
F51B
F535
F5A6
F60D
F6B6
F7BD
F895
F8E0
F904
F966
F997
F8EE
F7D2
F78B
F893
F9D4
FA13
F977
F907
F92B
F970
F97B
F97B
F99E
F9C1
F9B5
F980
F938
F8D3
F842
F7A1
F729
F6EC
F6CF
F6B8
F69C
F695
F73B
F997
FDEB
027E
04C2
0422
02B8
02AA
0397
03A5
027D
01C1
026D
0335
0298
01AE
0335
07C7
0C9B
0EB9
0E38
0D54
0D5F
0DE7
0E46
0E88
0EC1
0EA6
0E3F
0E35
0EC9
0F20
0E6B
0D62
0D65
0E55
0E9B
0DC1
0D59
0E63
0F19
0CF9
0865
0476
0327
033F
02B4
01C7
0228
038E
032B
FF1F
F91E
F490
F309
F3A0
F4F6
F65F
F754
F72A
F5F3
F4C5
F48B
F4FF
F55D
F5BB
F6C3
F837
F8D0
F80B
F730
F7B0
F923
F9D8
F92C
F847
F879
F99D
FA8B
FA96
FA0C
F97A
F908
F8B9
F8BD
F921
F986
F995
F983
F9B8
FA05
F9B1
F86B
F6D8
F605
F656
F719
F745
F6A3
F64A
F7B6
FB42
FF91
029D
0372
02E1
026D
02C0
034C
035D
030B
02E5
02FF
02D4
0227
01AF
029C
0573
0963
0CD9
0EBD
0F2D
0EF7
0EA1
0E26
0D88
0D25
0D4F
0DE4
0E88
0F18
0F9E
0FD2
0F38
0E00
0D47
0DD4
0EE6
0F04
0E10
0D71
0DCD
0DA5
0B24
06D1
0344
022D
02AC
02F5
02A3
0251
0198
FF20
FAE8
F70C
F55B
F538
F4EE
F449
F480
F5CB
F6AC
F617
F515
F546
F662
F69F
F586
F4E2
F636
F879
F976
F8B6
F7CF
F80F
F90C
F9B6
F9CC
F9C6
F9CC
F997
F925
F8E3
F8F7
F8EC
F86F
F7E7
F7F1
F88E
F945
F9BF
F9E0
F97C
F893
F79A
F728
F740
F758
F714
F6A1
F641
F5D9
F575
F600
F8B1
FD71
0240
04D4
04BC
0383
02EF
0367
040B
03FC
035A
0300
0355
03B8
0363
02E3
03ED
076B
0C08
0F34
0FB9
0ECD
0E5D
0EDB
0F52
0F33
0EFA
0EF0
0E92
0DAF
0D36
0DF6
0F43
0FBB
0F23
0E77
0E44
0E02
0D75
0D86
0E9B
0EE3
0C0A
06C4
02B9
0233
036A
036D
023C
0212
031B
0268
FDFA
F80C
F4B1
F4E2
F5E4
F57D
F4A9
F537
F68E
F6A7
F545
F440
F4BD
F5C8
F620
F623
F6ED
F85A
F91D
F8A8
F7F4
F7FB
F86E
F88B
F86E
F8AF
F930
F947
F8DB
F889
F899
F89B
F839
F7D7
F80E
F8CC
F968
F98D
F997
F9E5
FA2C
F9C6
F87E
F6C9
F578
F536
F5FB
F6C1
F669
F54D
F579
F8AB
FE21
02FC
04EE
0435
02E1
028E
0329
03B7
03B2
0366
035B
03B0
03F5
0397
02DB
0341
0639
0B1D
0F39
1073
0F68
0E52
0E4B
0E7D
0DF6
0D3D
0D60
0E43
0ED6
0EC4
0EC1
0F07
0EDA
0DFB
0D70
0DF0
0E8A
0E11
0D31
0D8B
0EC2
0E23
0A12
04B9
01C5
0208
030D
02FE
02CD
0382
035D
FFC5
F971
F458
F337
F4B2
F5B6
F55F
F52A
F5F1
F68E
F5E9
F4CC
F49A
F536
F579
F53B
F581
F6B6
F7E3
F80B
F78A
F778
F81D
F8BB
F8C1
F883
F897
F8F9
F943
F95F
F971
F966
F8FF
F857
F7D9
F7C9
F817
F898
F92B
F9A5
F9D4
F999
F8EF
F7E9
F6D2
F631
F668
F709
F6FE
F5D9
F4FC
F6A1
FB57
00E9
0465
04ED
0416
03C0
0426
044C
03B3
0320
0393
04D4
056D
044C
0251
01EB
04DC
0A3E
0EFE
10B3
0FD8
0ECD
0EE8
0F5C
0F0C
0E50
0E3B
0ED1
0F16
0EB3
0E7B
0F04
0F98
0F49
0E78
0E41
0E99
0E6F
0DB1
0DC0
0EFC
0F41
0C4E
0726
0353
02B3
0383
0341
0226
0212
02BC
0140
FC2B
F62A
F32E
F3D1
F53D
F537
F47E
F4C6
F5ED
F667
F5B2
F4EA
F4EF
F52E
F4E7
F4A1
F562
F6F3
F809
F800
F793
F7A6
F818
F83F
F807
F803
F87E
F903
F90A
F8B1
F876
F874
F856
F7F5
F7A3
F7BD
F83A
F8C8
F929
F955
F948
F8C5
F789
F5CE
F479
F46B
F582
F695
F6B3
F65E
F73B
FA5B
FEDD
028D
03DA
0331
0257
0295
03B4
0487
0458
03A6
037A
03FF
0428
0336
0251
03BE
082F
0D71
1074
106C
0F39
0ECF
0F13
0ED8
0E18
0DFA
0ED3
0F87
0F4D
0EE3
0F3D
0FDF
0FA8
0EBC
0E5D
0ED8
0EF9
0E19
0D7D
0E6B
0F80
0DD5
08F6
0408
020B
0274
02CD
0278
02D3
03D8
02EF
FE43
F7E3
F3EA
F3D2
F546
F5B7
F54F
F585
F647
F63A
F536
F4A1
F54E
F64E
F682
F64A
F6CB
F80C
F8D8
F887
F7E5
F7E9
F85B
F870
F825
F821
F89D
F91D
F94B
F953
F95B
F927
F888
F7D2
F78F
F7E0
F864
F8BF
F8EF
F910
F918
F8EB
F873
F795
F65D
F55D
F54E
F600
F64E
F5AF
F57E
F7D4
FCEB
0246
04DF
041C
0235
01B2
02EE
044A
0464
038F
0327
03C2
0469
03C8
022F
01ED
0508
0A9E
0F63
10FD
1030
0F54
0F5D
0F58
0E87
0DB1
0DE5
0EC7
0F37
0F1E
0F57
0FE0
0F96
0E45
0D76
0E3E
0F56
0EE1
0D56
0CF9
0E37
0E58
0AED
0564
019D
0141
0256
02AA
0290
030F
02FD
001D
FA9E
F593
F38C
F401
F4C4
F4D5
F4D5
F538
F573
F532
F50A
F570
F5D2
F5A0
F566
F605
F745
F827
F85E
F87D
F8C5
F8BF
F832
F7C7
F826
F8D6
F8D1
F80D
F7A8
F84C
F942
F990
F93D
F8E7
F8B1
F870
F85D
F8D3
F97F
F9A4
F917
F859
F7A3
F693
F534
F49E
F5A9
F740
F75A
F5FE
F602
F9CD
0011
04E5
05E6
044B
02E6
0312
03F9
0448
03DB
0393
03FE
048D
044B
0338
02D6
04FB
09BB
0EB0
1110
107C
0F15
0EB4
0F1E
0F4C
0F40
0F96
1011
0FDA
0F19
0EFE
0FD3
102B
0EE6
0D38
0D2F
0E90
0F0D
0DE5
0D3C
0E94
0FBB
0D52
079A
0298
012D
020B
0264
01F1
025A
034D
01E8
FCC9
F6B0
F374
F38E
F45B
F41D
F3C5
F4A7
F62D
F6C0
F5FB
F4FE
F4BA
F4FB
F537
F57B
F618
F6F6
F7CC
F886
F8F7
F8B6
F7D6
F73D
F79C
F86D
F8A5
F82E
F7E1
F829
F866
F7FE
F773
F7B4
F8A9
F941
F8FA
F885
F88E
F8B1
F84B
F79A
F739
F709
F672
F592
F530
F588
F5DF
F5CA
F64C
F8E8
FD8A
0214
045B
043C
0356
031E
03AD
042F
0405
0373
035B
0419
04D3
0478
0390
0436
07AD
0C82
0FD2
1066
0FBB
0FB2
102E
0FDA
0E9B
0DE5
0E7F
0F7B
0FDA
0FFB
1076
10B6
0FF1
0ECF
0E9E
0F16
0E90
0CDB
0C3E
0E37
1052
0E86
08A6
033A
01F2
0355
03A6
025B
0215
0396
03B6
FF9D
F923
F4E7
F4B2
F5E5
F5AE
F4A0
F4DC
F657
F700
F614
F52A
F5A5
F6B2
F6AF
F5A5
F544
F693
F894
F98A
F8F2
F7C1
F716
F748
F7FC
F896
F8A1
F82C
F7CC
F7F0
F84B
F83D
F7B1
F742
F77E
F843
F8ED
F90B
F8BE
F878
F870
F864
F7DF
F6B5
F55A
F4B1
F528
F616
F64F
F5A5
F57E
F77D
FBB3
0062
0381
045A
03D5
0354
036B
0389
02FB
020F
01EC
031A
0472
043F
02A4
0237
0550
0AF7
0F86
10A5
0F97
0F0B
0FA4
0FD8
0EBD
0D88
0DB6
0EDF
0F63
0EC3
0E20
0E5C
0EEE
0EFC
0EB1
0E9A
0E90
0E32
0DFE
0EB5
0FA1
0EB4
0AF0
0606
02A2
0195
018F
0191
0224
038D
0418
0199
FC56
F73C
F4DC
F514
F5F8
F64C
F642
F649
F62A
F5A3
F515
F4FC
F51D
F4F4
F4BB
F55C
F71E
F906
F9D2
F960
F8B3
F8AE
F921
F940
F8BC
F819
F7EF
F840
F896
F8A7
F895
F8A1
F8D7
F91B
F960
F99F
F9A8
F93A
F876
F7FA
F83A
F8BD
F880
F73C
F5FC
F5F1
F6E4
F745
F629
F4CD
F59E
F99E
FF0F
0302
040F
034D
02C1
0337
03D2
0386
0291
0234
0317
044B
045D
0347
02DF
04F6
092C
0D20
0EDC
0EB1
0E65
0EE2
0F62
0EEF
0DF0
0D95
0E32
0EE1
0EDD
0E85
0E9B
0EFE
0EE0
0E23
0DAA
0E0F
0EA8
0E86
0DF8
0E29
0F12
0EC3
0B8D
0677
029B
01D7
02F2
0378
02C1
0232
02A7
02CA
00AB
FC5F
F822
F5DE
F560
F538
F4B6
F451
F48A
F52B
F5C1
F630
F674
F641
F572
F49D
F4BA
F5F8
F778
F854
F898
F8CB
F8FB
F8C8
F846
F82C
F8D2
F982
F951
F86F
F80B
F8CF
F9F7
FA48
F991
F8B6
F865
F865
F83E
F81C
F88A
F972
F9F2
F94C
F7C0
F63E
F579
F57F
F60A
F6C0
F714
F683
F569
F55A
F7F2
FCF3
01F5
0477
0431
0312
02EB
039B
03CE
031F
02A7
0350
0461
0451
02F6
0229
03EB
082C
0CBC
0F54
0F91
0ED0
0E8F
0F21
0FD8
100D
0FB6
0F2C
0EA3
0E1E
0DBF
0DD8
0E6A
0EE1
0EB3
0E2D
0E1C
0E97
0EB6
0DEA
0D21
0DB0
0F09
0E8F
0A8F
04E0
0154
0182
0333
0387
0275
020C
02C6
0254
FEAE
F91C
F50E
F43E
F537
F5BA
F566
F53C
F598
F5CD
F589
F564
F5C8
F627
F5E6
F57D
F5F2
F758
F890
F8C3
F862
F850
F88E
F875
F7F9
F7E6
F8B2
F9BA
FA04
F976
F8E2
F8E2
F92F
F929
F8B1
F837
F81F
F86C
F8EF
F96A
F989
F90E
F81E
F748
F6EA
F6CC
F676
F5E5
F598
F5C3
F5DC
F563
F511
F6AA
FB0A
00A8
048B
051A
0399
02A9
036B
04A1
0494
034C
0254
029C
0355
034A
02CA
0391
06AF
0B11
0E61
0F48
0E7D
0DC4
0E1A
0F0E
0F9C
0F51
0E8B
0DF0
0DD2
0E0D
0E45
0E30
0DCC
0D72
0DA5
0E92
0F9E
0FCE
0EE1
0DDC
0DDF
0E6D
0D7D
09D4
04F6
01F8
022A
03AA
03DC
02AF
0252
03AA
0466
019B
FB9E
F618
F41E
F526
F65D
F62B
F566
F55A
F5E4
F60A
F5AC
F58F
F610
F693
F686
F645
F69E
F7B6
F8E7
F992
F9AC
F972
F90A
F89E
F87F
F8C4
F907
F8CE
F842
F80F
F886
F928
F947
F8E1
F895
F8C6
F91C
F90C
F891
F82D
F846
F8B1
F8E4
F86F
F74E
F5FC
F531
F552
F5F2
F615
F55B
F4D4
F64E
FA6F
FFA9
036A
0476
03D7
0372
03F0
046B
03F2
02E8
0272
02E9
0360
02ED
0220
02B9
05C6
0A42
0DD5
0EF3
0E26
0D31
0D2F
0DD4
0E48
0E58
0E75
0ECB
0EEB
0E79
0DD5
0DA8
0DF3
0E18
0DCD
0D8B
0DC3
0E1C
0E03
0DC7
0E4A
0F5F
0F28
0C09
06F8
0301
0216
0312
037C
02B5
0256
0363
0438
022A
FCEC
F74B
F45C
F481
F5A7
F5F2
F572
F53C
F5C0
F66D
F69B
F646
F5D6
F5A0
F5CF
F677
F77A
F86D
F8E6
F8EE
F8F7
F942
F986
F95A
F8C7
F84C
F844
F88E
F8D4
F8FA
F91F
F940
F929
F8D1
F895
F8D8
F978
F9D9
F98D
F8D9
F85D
F85F
F875
F7FB
F6D3
F59D
F539
F5E1
F6C7
F6B7
F561
F425
F534
F981
FF70
03EA
050C
03BD
0288
02EB
0423
047E
038B
0289
02B6
03B2
03F1
02CF
01C6
0321
0776
0CA7
0FB0
0F87
0DF7
0D8A
0ED5
1035
1004
0E8A
0D67
0D8E
0E62
0EBF
0E54
0DB0
0D63
0D91
0E26
0ED2
0EE6
0DEB
0C9A
0C8A
0E1B
0F40
0D56
0861
0393
01EC
02FB
03D0
02EC
01DA
026E
0395
024A
FD7E
F7C4
F499
F4C5
F62B
F6A2
F608
F57F
F594
F5E7
F619
F639
F649
F604
F568
F510
F5A6
F70F
F876
F926
F927
F8FA
F902
F93E
F978
F981
F948
F8ED
F8B1
F8B4
F8CF
F8C8
F8A6
F8A2
F8C8
F8D5
F896
F848
F862
F903
F9CA
FA2F
F9F2
F911
F7AF
F636
F561
F5A6
F67B
F699
F55C
F3E4
F466
F80F
FDA5
0272
048C
043D
0345
0306
0376
03AE
0334
028E
0296
0369
0426
03F4
034A
03DA
06DB
0B6A
0F08
0FF1
0ECC
0DC3
0E17
0F0E
0F54
0EC9
0E5E
0E8A
0EB6
0E57
0DDF
0E07
0E97
0EA9
0E14
0DC2
0E3C
0EB7
0E40
0D6A
0D97
0E83
0DCB
09DA
0484
016D
01E1
0382
0398
027C
0272
03A3
0334
FF00
F8DD
F4D7
F494
F5EB
F61F
F527
F4E3
F60B
F740
F732
F64C
F5C1
F5BA
F585
F50B
F517
F622
F78C
F86E
F89F
F884
F852
F80C
F812
F8DE
FA18
FA9D
F9DC
F8B6
F868
F8FC
F96B
F922
F8A6
F893
F8B0
F87D
F840
F8B1
F9B2
FA2C
F977
F849
F7AC
F7A1
F765
F6D3
F692
F6C5
F686
F552
F482
F657
FB43
00E2
042B
045A
0337
02BE
032E
0382
0329
02BB
02F9
03A8
03BC
02BB
01A6
0253
0599
0A3F
0DD8
0EEF
0E45
0DCD
0E84
0FA0
0FE7
0F4B
0ECA
0EF4
0F36
0ECB
0DE2
0D5C
0DA3
0E44
0EB8
0EFD
0F26
0EE1
0DFC
0D3C
0DB7
0F0F
0F0F
0BEB
06BD
02C4
01F4
02E9
0300
01D0
015E
02B1
0391
00EB
FAFA
F596
F402
F57B
F6BA
F61D
F4FC
F50D
F5E6
F601
F534
F4D6
F58F
F657
F632
F5CE
F682
F834
F95F
F929
F864
F83F
F8A9
F8C2
F857
F81B
F860
F897
F854
F81B
F88B
F941
F958
F8BE
F84E
F88F
F90D
F932
F926
F95D
F9A1
F946
F842
F75D
F710
F6DE
F64C
F5DB
F642
F712
F712
F63D
F681
F9C5
FF64
044C
05EE
04AF
0322
0321
0421
0461
033D
01E7
01DA
02FE
03C1
0334
029B
042E
0855
0CCC
0EFA
0EAF
0DEC
0E36
0F01
0F06
0E59
0E33
0EF6
0F82
0EE7
0DD6
0D99
0E3B
0EA0
0E52
0E1A
0E97
0F16
0E9D
0DA3
0DA7
0ED7
0F28
0C97
07D8
03D7
027A
02CF
02C7
0207
01FB
033D
03ED
0187
FC0E
F68B
F3FD
F467
F56B
F55F
F4DD
F532
F646
F6DA
F66F
F5F3
F63F
F6D1
F6A1
F5DF
F5CD
F6F0
F840
F89D
F84F
F861
F907
F96A
F90F
F893
F8AA
F917
F91C
F8B8
F8A4
F91B
F966
F8EB
F816
F7BD
F809
F87E
F8D2
F919
F945
F90B
F86B
F7D2
F779
F70B
F647
F5AB
F5D8
F66D
F64F
F578
F5B6
F8D0
FE29
02FE
0509
047A
034C
0313
03C0
043A
03D6
0305
02B7
0333
03AF
033C
024F
02E8
0681
0BD8
0FAA
100E
0E79
0DC8
0ED2
0FDA
0F43
0DB7
0D04
0DA5
0E6D
0E72
0E33
0E71
0EDD
0EB5
0E21
0DF8
0E56
0E6B
0DE4
0DA6
0E6D
0F25
0DA7
095A
0462
019F
01C4
0301
036C
0307
02ED
032A
0236
FEC3
F9AA
F575
F3F6
F4AC
F5AD
F5D2
F582
F58E
F600
F649
F61C
F5A5
F520
F4BB
F4D5
F5DE
F797
F8E9
F8FA
F84D
F829
F8E4
F976
F901
F816
F7E1
F882
F8FC
F8B6
F834
F832
F887
F889
F832
F82A
F8B7
F949
F961
F93F
F94A
F949
F8C0
F7C6
F6E6
F665
F624
F632
F6C0
F768
F72A
F5D1
F504
F6FB
FBE2
013C
0458
04DD
0470
045B
046F
0402
0330
02BD
030B
03B1
03FA
03A3
032D
03A4
05E9
09CE
0DCA
1008
1012
0F22
0EAB
0EE3
0F11
0ECA
0E58
0E0D
0DDF
0DC2
0DEC
0E6F
0ED7
0EAF
0E48
0E6E
0F31
0F89
0E9E
0D18
0C84
0D79
0EB5
0E42
0B57
071D
03B2
024E
0259
0255
01A9
0146
0244
03FD
0421
010B
FBD0
F75D
F591
F5AE
F5DE
F56A
F4F9
F514
F568
F573
F558
F57D
F5D3
F5E8
F5A7
F596
F62F
F744
F847
F8E7
F928
F920
F8E5
F898
F850
F80C
F7DB
F7EE
F847
F885
F848
F7BE
F783
F7EF
F8A2
F903
F8FB
F8E9
F904
F918
F8F9
F8C0
F87B
F7F3
F721
F668
F620
F621
F61F
F63B
F6AD
F703
F670
F53B
F545
F84D
FDAA
0281
049A
0462
03D6
03FE
043F
03D0
02FE
02B5
0346
0403
040E
035A
02E8
040B
073B
0B61
0E76
0F34
0E55
0DBD
0E5D
0F64
0FA8
0F2E
0ED7
0EED
0EDA
0E41
0DA6
0DAB
0E1B
0E42
0E00
0DF2
0E6B
0EE5
0EBE
0E32
0E02
0E64
0E99
0D88
0AB3
06B1
030E
0148
0182
0256
0247
017E
0177
02BD
0389
016F
FC71
F76F
F52C
F585
F636
F5D4
F504
F4F9
F5AC
F622
F5EB
F59B
F5CB
F64E
F697
F6A6
F701
F7EB
F8F8
F983
F957
F8D6
F88F
F8B7
F8FB
F8DC
F84A
F7AE
F772
F799
F7F7
F87F
F924
F9A2
F99E
F922
F8A9
F893
F8B4
F8AC
F87E
F86E
F85A
F7CD
F6D1
F619
F616
F659
F655
F64A
F6C0
F748
F6C7
F561
F553
F8C3
FED0
03DF
053C
03CF
029C
032E
045B
0462
032E
0235
0285
039B
0427
03AA
032A
0455
07D9
0C7C
0FE3
1099
0F67
0E62
0EA5
0F5D
0F3E
0E41
0D73
0D65
0D99
0D71
0D18
0D21
0D9E
0E15
0E43
0E67
0EA9
0EB3
0E3A
0DA4
0DA9
0E48
0E75
0CE1
0934
049B
012B
0039
0128
0208
01B6
011E
01E5
03E0
0488
01A0
FBFD
F6F2
F4E0
F51E
F581
F520
F4CA
F53D
F602
F63D
F5D9
F56B
F554
F581
F5F7
F6F1
F84D
F950
F968
F8E9
F8A1
F8DC
F927
F90E
F8A8
F85F
F872
F8C4
F90B
F915
F8F2
F8DA
F8F7
F934
F955
F92A
F8BE
F849
F803
F80D
F870
F8F0
F908
F862
F764
F6D2
F6D5
F6CB
F655
F612
F6A9
F77D
F721
F587
F4EF
F7C6
FDA5
0337
057E
04AB
0346
031D
03C7
0403
039A
0377
0435
0525
0514
03D8
02E9
0427
07EF
0C7F
0F64
0FB3
0EB3
0E43
0EC8
0F33
0EC9
0E2B
0E3C
0EB9
0EA1
0DBE
0D03
0D38
0DFC
0E68
0E5D
0E7A
0EEA
0EF1
0DF9
0CAA
0C44
0D07
0DA3
0C68
08ED
04A4
01BF
0159
026F
02FB
0230
015F
022D
0409
0426
0083
FA89
F5E3
F4AE
F5A1
F625
F563
F484
F48C
F51D
F572
F58F
F5E3
F649
F636
F5D7
F62E
F7AF
F951
F9A0
F888
F77F
F7C6
F90D
FA01
F9E2
F928
F8C1
F8F7
F94A
F93B
F8E0
F89F
F89C
F8A9
F8AC
F8C5
F8F7
F904
F8CD
F8B4
F92B
F9E1
F9BD
F82E
F632
F56A
F622
F6F7
F6B5
F5DA
F5A8
F628
F62B
F56B
F5B0
F8EB
FE7D
0351
04FA
0414
031C
037B
0473
04B3
041B
03A4
03F4
0485
0452
0346
02BE
046D
088D
0D39
0FE0
0FA2
0E0F
0D63
0E29
0F0B
0EE2
0E29
0E02
0E7D
0EA9
0E22
0DAB
0E04
0EBA
0EC5
0DFE
0D52
0D65
0DAD
0D57
0CAA
0CC0
0DD4
0E74
0CC9
08AA
0423
01C5
023C
03BC
03ED
0273
0125
01A8
031A
02B4
FEE1
F938
F502
F3F2
F4DA
F58F
F54D
F4DB
F4FD
F58C
F60D
F660
F696
F68D
F62F
F5E2
F64A
F771
F897
F900
F8CF
F8B0
F8EA
F921
F8FF
F8BD
F8D4
F94F
F9AC
F981
F910
F907
F9A3
FA52
FA55
F9A9
F900
F8CD
F8B8
F845
F7BE
F7FB
F91D
F9FB
F95D
F784
F5ED
F587
F5D2
F5F9
F60C
F684
F709
F6C2
F60A
F6DC
FAB5
004D
045F
04EF
0341
0225
02D8
042A
047D
03BF
0333
03AF
049A
04BB
03D8
0352
04E6
08D3
0D3D
0FB9
0F84
0E25
0DAB
0E7C
0F40
0ED0
0DA8
0D21
0DA9
0E6C
0E8F
0E2F
0DF3
0E18
0E49
0E45
0E3B
0E57
0E5C
0DFA
0D6F
0D58
0DCB
0DD4
0C25
0878
0437
0189
015F
0292
032C
0290
01F5
0276
032A
01D2
FD82
F812
F472
F3CA
F4C7
F582
F570
F535
F541
F55E
F555
F553
F570
F571
F540
F566
F67A
F83B
F98D
F9A5
F8E4
F84D
F852
F88C
F888
F875
F8C4
F965
F9C1
F974
F8E0
F8BB
F926
F97F
F93B
F8AE
F895
F906
F944
F8D5
F84B
F87C
F92D
F91B
F7A6
F5DB
F547
F606
F6C2
F6A6
F667
F6DE
F770
F6EE
F5DC
F6A0
FAC1
008C
0473
04C5
0341
02BD
03E9
051B
04D0
0389
02E0
0374
044C
042D
0349
0348
05A2
09F7
0E1D
0FF9
0F51
0DDC
0D70
0E4A
0F2A
0F02
0E23
0DA7
0E14
0EE8
0F51
0EFA
0E28
0D64
0D24
0D97
0E82
0F56
0F90
0F31
0EC7
0EC8
0EE6
0E11
0B6B
0752
037D
01BE
0253
0395
039E
0264
019B
0258
0345
01D0
FD34
F7AA
F44E
F41A
F55F
F5FD
F57E
F4DD
F4DE
F54D
F597
F58D
F563
F553
F580
F606
F6DD
F7C3
F856
F871
F84C
F83A
F85E
F89E
F8DF
F914
F931
F927
F904
F8FB
F937
F9A8
F9F4
F9B9
F906
F86D
F869
F8B6
F8A6
F81F
F7F0
F8C4
F9FB
FA1B
F897
F6A5
F5E4
F673
F70D
F6E6
F68D
F6A8
F6B4
F5F7
F550
F6E5
FB81
0101
0437
0439
0314
0311
041F
0479
035A
0217
0253
03DA
04D6
040F
0291
02C2
05EE
0AD1
0EA9
0FB1
0E87
0D47
0D6A
0E9F
0F8A
0F4E
0E48
0D71
0D58
0DD2
0E50
0E5D
0DE8
0D5A
0D50
0E01
0EF8
0F6D
0F03
0E28
0DB9
0E29
0EDD
0E6B
0BB2
0728
02EA
0125
01FD
034D
02FE
0172
00E6
0250
039B
01CD
FC9B
F70A
F44E
F4B7
F60C
F661
F5C6
F54F
F56A
F5B1
F5C3
F59C
F53E
F4B1
F45D
F4E0
F64F
F7E1
F8B6
F8BF
F8A6
F8DE
F928
F91D
F8DA
F8CF
F914
F946
F91C
F8D4
F8E3
F95A
F9CA
F9BD
F944
F8E1
F8E3
F90B
F8F3
F8BF
F8FD
F9C7
FA56
F9C8
F847
F6F4
F69B
F6C6
F692
F603
F5E8
F673
F6BE
F648
F649
F89B
FD3D
01D1
03EC
0398
02F0
0375
0480
0490
0375
0281
02C3
03B5
03FA
0316
0224
02DA
05ED
0A5D
0E32
0FF7
0FA9
0E7B
0DCE
0E31
0F19
0F7A
0EC2
0D6C
0C91
0CDE
0DDD
0E6E
0E07
0D53
0D64
0E5A
0F39
0F1F
0E3C
0D78
0D72
0E0F
0E94
0DEE
0B36
06AE
024F
0090
01E9
03FF
0418
0243
0112
01F3
02E7
00D9
FB9E
F666
F41D
F47A
F522
F4DE
F484
F501
F5CE
F5E9
F573
F55A
F5C8
F5E7
F54B
F4CB
F575
F720
F890
F8EC
F894
F873
F8DC
F95F
F98C
F96B
F93F
F91D
F8FF
F905
F959
F9D8
FA0B
F9A1
F8F2
F8CE
F989
FA6B
FA6E
F984
F8B3
F8C0
F911
F872
F6BD
F547
F557
F693
F76A
F6F0
F5D9
F58D
F6E0
F9C7
FDBD
01D4
04B8
0584
04B7
03E1
0400
048A
0456
034D
0288
02BA
0334
0304
02B1
0402
07D4
0CA7
0FCB
0FF3
0E52
0D2D
0D8B
0E94
0F05
0EB7
0E67
0E6C
0E44
0D8F
0CDD
0D0B
0E02
0EAB
0E3F
0D3E
0CAB
0CD7
0D5B
0E07
0EDB
0F0C
0D25
08E3
0458
0219
0276
0359
0326
0297
02FE
0383
01A9
FCCA
F79E
F54F
F5EA
F6C7
F619
F4B5
F43B
F4B9
F504
F4B5
F49E
F53C
F5CE
F590
F51B
F5B1
F775
F921
F996
F90F
F88C
F88F
F8C7
F8C1
F878
F83A
F83F
F891
F91E
F9AE
F9EB
F9A4
F918
F8CA
F90A
F9BA
FA6F
FAC1
FA8E
FA17
F9BA
F974
F8CE
F776
F5E0
F510
F589
F698
F6EE
F616
F521
F5D2
F8FB
FDB7
0207
044A
045F
038A
0332
0394
03CD
033A
0276
0298
03A1
0432
034B
01F3
028C
0633
0B3A
0EB0
0F39
0E19
0D68
0DDC
0E90
0E94
0E1F
0E03
0E71
0EC5
0E83
0DF9
0DAB
0D88
0D37
0CF5
0D69
0E76
0EEC
0E01
0CB8
0CCC
0E10
0DEA
0A60
0512
01DC
0257
040F
03E9
0228
0192
0305
03A2
0054
FA05
F4DD
F394
F4E4
F5FA
F5EF
F5D8
F64F
F689
F5DB
F4EC
F4B3
F51E
F576
F5B9
F69F
F839
F968
F93B
F843
F7DD
F87F
F952
F977
F8FC
F87F
F853
F861
F888
F8BB
F8CD
F89A
F868
F8C5
F9C7
FAB8
FACE
FA20
F978
F957
F965
F906
F817
F706
F651
F628
F673
F6E2
F6FC
F665
F57B
F586
F7D6
FC61
0168
04B4
0562
0475
03A2
03AF
0403
03CB
0326
02EC
036C
03D9
034F
023A
0252
04DE
092D
0D0D
0ECE
0E9D
0DEE
0DCB
0E1E
0E56
0E4D
0E36
0E0F
0DA8
0D32
0D48
0E1B
0EE8
0EB6
0DA8
0CF4
0D51
0DF2
0DC1
0D32
0DC9
0F8F
0FF9
0C91
065C
016D
0093
026D
0396
02FE
028F
037B
03C2
00A4
FAAC
F59A
F421
F523
F5C3
F522
F4B1
F558
F5FD
F56E
F45F
F465
F58A
F64A
F5E8
F58C
F695
F895
F9DB
F9A9
F8F2
F8DB
F94D
F975
F917
F8B3
F8A6
F8C9
F8ED
F918
F934
F901
F888
F855
F8D3
F9A2
F9F2
F98B
F915
F929
F978
F942
F84C
F71D
F64C
F60B
F64B
F6D9
F740
F6DD
F5AC
F4E3
F64C
FA8B
001B
0454
05AD
04E4
03F0
03F7
0473
0446
0357
02BD
0344
0439
042A
02E8
0245
044A
08CD
0D4E
0F54
0EBA
0D67
0D0D
0DA7
0E34
0E3F
0E36
0E71
0E9C
0E4D
0DBC
0D87
0DD6
0E31
0E41
0E4D
0EA6
0EF6
0E9B
0DD3
0DC0
0EBD
0F2F
0CE5
07E9
0314
013D
0235
0361
0321
0288
0316
03CB
01EF
FCCE
F736
F47D
F4DC
F5D1
F589
F4A8
F481
F4F2
F4F9
F4A2
F4F8
F615
F699
F5B8
F4B6
F556
F75B
F8CE
F8A2
F7F6
F853
F993
FA4E
F9ED
F945
F922
F933
F8DE
F85D
F847
F885
F886
F847
F861
F8FA
F95B
F8EE
F825
F7EA
F864
F8D5
F8B6
F849
F7F4
F798
F6F9
F65A
F607
F5A2
F4B3
F3E1
F4E9
F8D3
FE6E
0309
04CD
0439
033E
0337
03EE
0458
03F4
0353
0359
040E
0469
03A1
02A2
0387
073B
0BFE
0EF0
0F04
0DE1
0DAC
0EA3
0F5B
0F01
0E52
0E36
0E67
0E20
0D93
0DC1
0EDB
0FC2
0F77
0E7C
0E0F
0E71
0EB2
0E4F
0E1B
0EDB
0F74
0DA6
08E2
039E
0104
0199
02FB
030A
0251
02A2
03D2
0337
FEF5
F8D8
F4CB
F48B
F614
F67D
F564
F4A1
F545
F637
F60F
F51A
F4B9
F555
F5FF
F623
F66C
F78D
F8FF
F9B5
F99D
F986
F9CA
F9D1
F931
F876
F865
F8E6
F93B
F91A
F8EA
F8E2
F8AA
F825
F7E3
F84D
F8DA
F8C8
F84F
F84C
F8E3
F92C
F87C
F762
F6D5
F6CB
F67A
F5BC
F55E
F5AF
F5CA
F519
F4EE
F76D
FCCA
026F
055C
04FE
0351
0285
02FE
03B1
03CD
038E
039D
041A
0467
03EB
0313
0367
062B
0AB3
0E8C
0FBE
0EB7
0D9B
0DC8
0E9E
0ECE
0E2F
0DAC
0DB8
0DC9
0D7B
0D63
0E1E
0F25
0F55
0E89
0DD1
0DEA
0E3C
0DF4
0D7E
0DF2
0F06
0E9A
0B12
05AF
01A0
00BA
01D1
029E
0282
028E
0327
02C4
FFBE
FAB5
F658
F4A7
F51A
F5C7
F5BC
F589
F5CE
F62E
F60A
F585
F53F
F552
F54C
F52E
F5B5
F751
F93D
FA30
F9D5
F914
F8D0
F8FF
F920
F91A
F918
F8F8
F880
F7FF
F826
F906
F9BA
F96A
F869
F7D0
F817
F8A6
F8D8
F8D5
F912
F962
F929
F83C
F71A
F644
F5D2
F5C5
F632
F6D4
F6E0
F5FE
F560
F71E
FBDF
0195
0518
052C
037C
0295
034D
0460
045E
036F
02F9
03B7
04B8
0483
0323
028A
04A7
0926
0D80
0F66
0EF1
0E1E
0E5B
0F2F
0F58
0E9B
0DE3
0DD6
0E1A
0E17
0DF2
0E34
0EC9
0EFC
0E85
0E08
0E2B
0E96
0E7E
0DF7
0DF6
0EAD
0E99
0BFE
0748
031D
01AC
026C
0316
0295
01FD
0266
02B2
0095
FBB0
F68B
F407
F468
F596
F5D1
F551
F521
F55F
F554
F4D3
F48C
F4F7
F5A4
F607
F654
F710
F814
F8AD
F89B
F861
F87D
F8C3
F8C7
F893
F887
F8A7
F89C
F860
F868
F8E7
F95D
F946
F8E0
F8CA
F917
F93E
F8F0
F888
F874
F898
F894
F855
F809
F79B
F6D4
F602
F5E3
F684
F6D0
F5EC
F4D4
F5CC
F9E2
FF6F
0379
047B
038B
02D7
0355
0435
0446
037B
02EB
0368
045E
045E
02F3
01C2
032C
07A9
0CE6
0FEA
0FFD
0EFA
0EE4
0FC8
104D
0FB6
0EB3
0E35
0E45
0E5D
0E53
0E55
0E50
0E08
0DC1
0E21
0F1B
0F93
0EAB
0D3C
0D20
0EB1
0FBB
0DA7
08A3
03CC
01E8
028C
031F
0244
0140
01AE
02C4
01E6
FDE3
F8B3
F564
F4DC
F56C
F55E
F4D8
F4ED
F5B5
F636
F5EB
F571
F56B
F588
F528
F49F
F503
F69C
F84A
F8CA
F833
F7A7
F7E8
F8A8
F938
F951
F91D
F8D6
F8A4
F8A1
F8C6
F8DF
F8CA
F8BC
F8F8
F94F
F941
F8C3
F874
F8D3
F985
F9C4
F950
F887
F7B1
F6B8
F5CA
F590
F65C
F747
F6FD
F59D
F53C
F7D3
FCEE
01DE
044F
0449
038B
0367
03A6
0372
02B8
0251
02E2
03EF
0452
0391
02A8
034F
0655
0A9E
0DFE
0F21
0EA2
0E29
0EA1
0F7C
0FB5
0F1A
0E60
0E21
0E42
0E58
0E4A
0E49
0E57
0E42
0E1E
0E45
0EB2
0ECB
0E40
0DCC
0E52
0F2A
0E35
0A48
051E
01E2
01CC
02F8
0311
023B
0242
033F
02B4
FEB1
F8CA
F4A7
F3FE
F517
F57B
F4E2
F4BC
F591
F63D
F5C7
F4D7
F4A1
F52B
F57F
F549
F554
F64D
F7C6
F8C8
F8F7
F8C4
F8B5
F8CF
F8D1
F89E
F848
F7F9
F7F6
F873
F941
F9CD
F9BD
F95E
F930
F947
F951
F92A
F90A
F925
F962
F970
F914
F840
F71E
F629
F5F0
F66F
F6CF
F657
F5CA
F720
FB52
00CD
04A6
0570
045B
0388
03B9
0407
038D
02C1
02C4
03BD
047B
03E8
02A2
02B4
0589
0A44
0E4B
0FB9
0F0D
0E39
0E4E
0EB4
0E92
0E1E
0E13
0E74
0E97
0E3E
0DF2
0E19
0E5B
0E41
0E07
0E1D
0E34
0DB2
0D07
0D5C
0E8B
0E76
0B6F
06A1
02FA
01F0
0256
0286
0278
02D3
02D1
00A1
FC04
F74B
F4E8
F4ED
F59D
F5C2
F580
F53D
F4F6
F4B7
F4D2
F546
F56F
F4E5
F44C
F4A1
F5E2
F709
F780
F7C9
F861
F8E3
F8C7
F86B
F883
F8EC
F8E0
F844
F7E5
F844
F8CF
F8B9
F839
F835
F8E8
F988
F974
F91B
F935
F9B4
F9EF
F986
F897
F769
F669
F62E
F6CC
F75A
F6DB
F5D2
F658
F9F1
FF85
0412
0594
04B6
0389
0339
037B
03A8
0399
0392
03CA
0417
03FB
0345
02D2
043E
0835
0D27
1056
1074
0EDF
0DE9
0E3D
0EB0
0E59
0DC3
0DC2
0E30
0E7E
0EB9
0F27
0F6E
0F03
0E3C
0E02
0E6C
0E89
0DF7
0DBA
0E92
0F0D
0CCF
07E2
0342
0174
01CF
0235
0239
02DF
03BE
0271
FDB2
F7AF
F3F9
F3A6
F4AB
F4FC
F4C4
F514
F5BC
F5C9
F545
F529
F5B4
F60C
F5AD
F54C
F5CD
F701
F7EC
F817
F7F2
F7F7
F80A
F7FD
F80C
F877
F8F2
F913
F8E8
F8B9
F884
F833
F810
F881
F950
F9BB
F954
F889
F81C
F853
F8D8
F92B
F8FF
F82D
F6E9
F5EE
F5E8
F67D
F691
F5FB
F64C
F92E
FE2E
02DB
0512
04D1
03B1
031F
034F
03AA
03BC
0397
038E
03C6
03DF
0352
027B
030D
0682
0BE0
1010
10F7
0FA6
0EB0
0EF6
0F2B
0E47
0D31
0D50
0E61
0EE1
0E5A
0DF0
0E72
0F1F
0F06
0E77
0E3F
0E3F
0DF6
0DCC
0E82
0F4D
0DF5
099A
046F
0190
018D
0257
0278
029F
0364
0320
FFC4
FA15
F56B
F403
F4E4
F5B5
F597
F54E
F555
F530
F4A4
F473
F528
F606
F609
F577
F57F
F680
F798
F7F1
F7C3
F7C0
F80D
F841
F82E
F82D
F881
F8E3
F8E7
F89E
F87C
F8C0
F93B
F993
F994
F946
F8E3
F8AC
F8A1
F89F
F8AB
F8E4
F909
F87E
F71E
F5D1
F5BB
F6C0
F764
F69F
F58C
F69A
FACE
005E
045F
057E
04B6
03CA
038E
03A6
0372
02F4
02D0
036C
0435
0426
033F
031E
058C
0A48
0EC2
1096
0FFC
0F19
0F2D
0F6A
0ECF
0DDE
0DBE
0E62
0EB4
0E4E
0DFA
0E42
0E85
0E10
0D69
0D93
0E64
0EC1
0E86
0EBA
0F66
0E9D
0AE8
05C2
0240
017F
01D5
01B5
01C2
02ED
03BB
0167
FBC6
F647
F422
F4CE
F576
F4DB
F445
F4DB
F5DE
F60D
F58D
F568
F5C3
F5B9
F50A
F4C1
F5C2
F76D
F87D
F899
F85E
F83A
F817
F806
F859
F8FD
F947
F8DA
F840
F842
F8D2
F92D
F8FB
F8CA
F91B
F98F
F97A
F8DD
F859
F855
F89D
F8C5
F886
F7CC
F6D9
F646
F679
F704
F703
F674
F6DC
F9D1
FECF
032C
04C1
041F
038E
043C
052F
0500
03DF
033D
03C3
0464
03C3
023B
01E0
0457
08EE
0D2F
0F39
0F4C
0EFE
0F45
0FA8
0F55
0E78
0DF8
0E30
0E92
0EAC
0EB6
0EE0
0EB9
0DE6
0D05
0D09
0DCF
0E21
0D93
0D65
0E96
0FA8
0DCE
089D
0336
00E6
0188
0273
0240
01FE
0271
01E9
FE42
F855
F3C8
F302
F4A7
F5BE
F54B
F49F
F4D7
F572
F58D
F547
F549
F597
F5B4
F5AC
F626
F753
F86D
F8B5
F86B
F84C
F87A
F88F
F879
F8A5
F931
F989
F926
F85D
F7FE
F851
F8CB
F8D6
F896
F89A
F906
F962
F94F
F8FD
F8DC
F8F1
F8C4
F7F7
F6DF
F645
F67E
F6DF
F67E
F589
F58D
F807
FCB7
0192
0473
04DE
0419
03B4
0423
04B3
04A9
0423
03D5
0409
0425
0367
024B
02AB
05E9
0AFF
0F11
1035
0F36
0E41
0E6A
0F07
0F36
0F17
0F28
0F41
0EE5
0E51
0E35
0E8A
0E88
0E12
0E10
0ED7
0F48
0E70
0D56
0DBD
0F25
0E99
0A4E
0470
00F7
0120
0290
02F4
02A4
02BD
024E
FF5E
FA2F
F5A7
F404
F480
F4F5
F4BB
F4B8
F532
F537
F470
F414
F50D
F651
F642
F525
F4E4
F662
F85C
F925
F8B4
F83D
F869
F8BF
F8C4
F8B8
F8ED
F91A
F8DF
F880
F87C
F8BE
F8D1
F8A6
F8A2
F8E5
F91B
F904
F8D8
F8EC
F93C
F96A
F920
F845
F70C
F5FF
F5C9
F677
F70A
F684
F59B
F68F
FAA3
0030
040E
04C4
03B1
0316
03A6
044F
040A
0327
02BC
0340
0406
041A
0368
0324
04E3
08F1
0D7C
100D
0FFC
0EEB
0E95
0EEC
0ED6
0E21
0DC0
0E40
0EF6
0F0F
0EC7
0ECA
0EF1
0E8F
0DD4
0DC0
0E6E
0EBB
0E2B
0DE3
0EAB
0EF0
0C55
0719
025F
00B0
014D
01FA
022D
02E2
039B
01E8
FCCF
F6FF
F401
F433
F511
F4FB
F4C3
F572
F640
F5E3
F4D6
F4BF
F5D8
F67A
F5B5
F4E7
F5CA
F7E6
F93D
F902
F84F
F846
F8B0
F8D3
F8BA
F8F1
F972
F99F
F937
F8C5
F8C2
F8F6
F8F7
F8DA
F8E1
F8EA
F8B2
F871
F89F
F931
F990
F93C
F83E
F704
F61E
F604
F6A8
F72F
F69B
F529
F4D1
F795
FD16
0272
04F7
04A3
0386
033D
03A1
03C4
0369
032B
037F
0401
03D0
02C1
0201
034C
0737
0C38
0FAC
1025
0EB6
0D98
0DCC
0E8A
0ED7
0EC7
0ED4
0EDE
0E8A
0E1C
0E29
0E98
0EB7
0E4A
0DE7
0DEF
0DEF
0D92
0D9A
0EB3
0F98
0DDD
0926
0440
020E
024E
02AA
023A
023F
0333
02FB
FF5E
F981
F525
F45F
F57A
F5BC
F4D1
F453
F4EA
F588
F55E
F50B
F564
F60F
F62B
F5D1
F60B
F745
F89C
F90D
F8BD
F88D
F8DE
F94B
F971
F951
F90A
F8A8
F852
F83D
F869
F8A7
F8E0
F936
F9AD
F9F8
F9C2
F92B
F8B2
F8A3
F8C4
F8A5
F817
F736
F65A
F5FE
F65B
F6DB
F67A
F522
F465
F63E
FAE6
004D
03E5
04DE
0467
040A
042B
0437
03CE
0349
0333
0393
03DA
0389
02FE
0382
060F
0A07
0D77
0EF5
0EDA
0E7C
0E8D
0EBC
0EAC
0E9A
0EC9
0EE2
0E79
0DF1
0E02
0E7C
0E6D
0DAB
0D3E
0DC1
0E44
0DC4
0D02
0D96
0F2A
0F0E
0B63
05DE
0216
0175
0232
0260
024E
02DC
02EE
0063
FB53
F6A5
F4D5
F54A
F5A2
F4EC
F455
F4E2
F5E6
F63B
F5F3
F5E0
F617
F5FA
F592
F5CA
F712
F898
F94A
F91E
F8E3
F906
F921
F8D6
F868
F83E
F847
F843
F850
F8A8
F915
F930
F90A
F922
F994
F9D4
F970
F8C5
F883
F8B7
F8B8
F821
F74C
F6B4
F65A
F611
F5F0
F605
F600
F5DC
F6B5
FA03
FF77
0452
05DF
045F
02B3
02DE
03F5
03F6
02C9
0228
02D8
037C
02D4
0222
03F5
08BC
0DC4
101A
0F91
0E43
0DE0
0E57
0EDF
0F2A
0F47
0F15
0E7D
0DE1
0DB4
0DD5
0DCF
0DB2
0DE9
0E40
0E02
0D54
0D7A
0ED9
0F84
0D0A
07BA
02DC
0124
01E5
029B
026F
0298
0355
0282
FE57
F873
F480
F41D
F578
F607
F56F
F509
F57B
F604
F5F0
F593
F586
F5BA
F5F6
F687
F7B5
F8FA
F980
F93A
F8D0
F896
F850
F7F3
F7FB
F899
F91C
F8C6
F7F8
F7CE
F889
F926
F8EC
F87C
F8C6
F983
F9A5
F909
F8AC
F913
F953
F83F
F62A
F4C3
F50C
F61D
F655
F589
F57C
F7FF
FCEA
01FA
04C0
04BE
039E
033F
03C0
03ED
034F
02E4
0378
042B
03A7
026A
02D2
0654
0B68
0F06
0FDA
0F25
0E97
0E7F
0E70
0E88
0F09
0F7C
0F36
0E74
0E15
0E42
0E4A
0DEA
0DE4
0EAB
0F50
0EC5
0DBA
0DD6
0EDE
0E50
0AA1
05B2
02AB
0241
0293
0263
0287
0391
03B0
0080
FA9C
F592
F3F1
F4B4
F558
F51E
F50F
F597
F5D4
F538
F488
F4A9
F563
F5F3
F64B
F6FC
F808
F8B4
F8AD
F894
F8ED
F940
F8E9
F83D
F80D
F867
F89D
F878
F88B
F935
F9DE
F9BD
F8FF
F891
F8E4
F964
F968
F915
F8DF
F89B
F7C0
F666
F572
F590
F654
F695
F5CA
F4FF
F631
FA50
FFCE
03BB
048C
0390
0335
0420
04B8
03B9
0246
025F
03DB
0469
0308
01F8
041A
0918
0D9F
0F33
0E9D
0E30
0EC1
0F51
0F1C
0EA2
0E8C
0EA0
0E6D
0E2D
0E40
0E6A
0E44
0E10
0E3D
0E80
0E40
0DDA
0E6C
0FE0
101D
0D32
080A
03CA
0259
029C
02AC
0271
02E3
036A
01CC
FD1A
F778
F41B
F3FA
F538
F5BC
F558
F52C
F5B1
F637
F609
F551
F4BA
F4B2
F536
F609
F6EE
F7C5
F879
F8D8
F8B8
F840
F7F5
F836
F8C2
F8F9
F8AE
F872
F8D6
F982
F994
F8DD
F83D
F877
F92A
F968
F8F8
F884
F88A
F8AD
F83D
F72C
F636
F608
F684
F6DB
F668
F58A
F5C3
F89B
FDDD
030E
0567
0498
02FF
02CD
03AA
03D5
02F6
029B
03B5
04E0
044A
02B0
02F9
069F
0BA0
0ED1
0F5A
0EEA
0F08
0F72
0F37
0E5D
0DB7
0DB7
0E17
0E7E
0EC8
0EBC
0E2F
0D9D
0DD2
0EA3
0EE3
0E15
0D78
0E4D
0F84
0E7A
0A44
053A
0261
0216
0268
0240
0282
0391
0374
FFF7
FA05
F53F
F407
F52A
F5EE
F564
F4C6
F519
F5C4
F5CA
F546
F4FB
F526
F57F
F60F
F719
F84B
F8D9
F882
F7FA
F7F8
F851
F864
F824
F819
F877
F8BD
F892
F861
F8BC
F972
F9D5
F9AF
F967
F94B
F935
F8F1
F8A4
F874
F821
F74B
F624
F57B
F5D3
F6A2
F6C9
F5F2
F54A
F6AF
FAED
0090
04BB
05A4
0442
031D
0373
042F
03E4
02F4
02D8
03B7
0403
02ED
023D
047B
097D
0E1B
0FAF
0ECE
0DE9
0E21
0EA2
0E86
0E21
0E2D
0E9C
0ED4
0E9E
0E4A
0E11
0DF0
0E02
0E59
0E84
0E0E
0D8B
0E22
0F8A
0F81
0C5D
0777
03E9
02FA
031C
02A5
0235
031F
044F
02C0
FD6F
F74F
F424
F466
F57F
F572
F4CD
F4EB
F5BB
F620
F5B2
F529
F524
F576
F5D6
F684
F7B2
F8D3
F931
F8DF
F884
F86E
F863
F83D
F82F
F84E
F866
F856
F858
F89C
F8E5
F8D4
F88B
F898
F91F
F997
F98D
F949
F943
F93A
F870
F6C9
F542
F4FE
F605
F712
F6D9
F5AC
F59D
F88B
FDE6
02C2
0494
03C1
02F4
03D9
0534
04E1
0307
01FB
02EF
0432
03BC
0256
02DF
0692
0B5C
0E54
0EDE
0E90
0EAF
0EF5
0ED2
0E8A
0E87
0E8A
0E3F
0E03
0E41
0E8E
0E41
0DB2
0DD4
0E9A
0ECB
0DE2
0D33
0E08
0F38
0E01
099F
04AB
0216
01F4
0250
0248
02A3
0361
0291
FEA8
F919
F53C
F4A6
F5BA
F624
F593
F542
F5B6
F629
F5FE
F59B
F58B
F5AF
F5BA
F5F7
F6F4
F87C
F990
F98C
F8EA
F890
F8B3
F8DA
F8BA
F894
F8B3
F8F6
F908
F8CF
F887
F87D
F8C2
F918
F92F
F8F6
F8AD
F8A9
F8FA
F93E
F8EE
F7E2
F695
F5D1
F5EA
F65B
F638
F54B
F4E4
F708
FC38
022D
058C
052F
0337
0276
034F
03E6
0323
0248
02EB
045B
0477
0300
0290
0581
0AC6
0EFA
101B
0F2D
0E50
0E4E
0E92
0EAB
0EC2
0ED7
0E8E
0DF6
0DB6
0E12
0E6E
0E46
0E03
0E30
0E6A
0DFA
0D47
0D84
0E97
0E66
0B27
0601
0226
0151
0236
02CB
02D0
030B
02E7
008E
FB96
F658
F3B6
F41D
F57E
F5F9
F5A8
F59D
F621
F686
F657
F5D4
F571
F569
F5D7
F6C0
F7DA
F8A4
F8DE
F8BA
F892
F88B
F8A6
F8E9
F944
F96A
F915
F88A
F86C
F8DA
F930
F8E2
F84F
F835
F8A3
F8E8
F898
F81F
F813
F84D
F807
F6F4
F5D8
F5B9
F688
F707
F63D
F4EF
F558
F8FE
FEC8
038D
0507
0401
031D
0397
043B
03B9
02C4
02FE
044D
04C4
037F
0274
044F
08FE
0D94
0FA1
0F7E
0EEC
0EB7
0E96
0E6E
0E83
0E9A
0E31
0D8D
0DAA
0EAF
0F59
0EAB
0D92
0DA2
0EA2
0EC7
0DA0
0D04
0E1F
0EFB
0CBB
07B1
035E
022C
02D2
02CC
020D
026B
03DF
0389
FF5E
F947
F525
F479
F56A
F5C4
F55C
F535
F59D
F5FD
F604
F601
F61B
F616
F601
F677
F7B8
F901
F96D
F914
F8BE
F8BA
F8A6
F84D
F801
F814
F860
F891
F8A2
F8C5
F8F5
F8FA
F8D3
F8BA
F8BC
F8AB
F897
F8DB
F962
F952
F80B
F626
F502
F54D
F652
F6CD
F634
F546
F57A
F7F7
FC8F
0186
049C
04EA
03BD
031F
0398
03FE
0381
02ED
0337
03CB
0365
0260
02EC
0671
0B73
0EF5
0F99
0EA0
0DE8
0DEF
0E30
0E66
0EA0
0EAD
0E4C
0DB7
0D65
0D5B
0D53
0D73
0E1A
0EE7
0EC3
0D7D
0CA1
0D8E
0F06
0E13
09D2
04F8
02B1
0300
037F
030C
02DD
03BE
03E1
00E3
FB37
F629
F43B
F4C0
F583
F5A0
F5B2
F613
F642
F5F6
F5A7
F5BC
F5F1
F5F5
F616
F6CC
F7E5
F8A0
F8AB
F877
F878
F884
F861
F850
F8A5
F92D
F96E
F959
F931
F8FB
F88C
F80C
F7F0
F85A
F8D1
F8E0
F8B9
F8D8
F925
F8E3
F7BB
F655
F5A7
F5F3
F6A2
F6DD
F643
F574
F60F
F96B
FED6
0387
0524
0427
0325
03A3
0483
041A
02E4
02D1
0428
04DA
039F
025C
0405
08BF
0D7F
0F89
0F1B
0E47
0E3C
0E8C
0E97
0E79
0E6A
0E3B
0DE6
0DD9
0E30
0E56
0DFD
0DD0
0E65
0F0C
0EAE
0DAD
0DA2
0EDD
0F3C
0C96
07C6
03F0
02C7
02F2
029E
0239
0310
0430
02AC
FD64
F72A
F3EF
F489
F64A
F693
F585
F4D4
F521
F596
F581
F53A
F53F
F578
F5AB
F620
F738
F8A2
F98B
F98F
F912
F898
F82B
F7B6
F785
F7ED
F8B1
F91F
F8F1
F893
F881
F8AA
F8AC
F873
F85A
F8A0
F916
F94B
F8E5
F7C4
F63C
F529
F54A
F63F
F69F
F5BD
F515
F71B
FC40
01D9
04A8
0441
0318
0342
0447
0495
0402
03BB
0421
0423
032A
02A4
0497
08F4
0D3B
0F20
0EC6
0E05
0E1D
0EBF
0F0A
0EAD
0E17
0DE8
0E53
0EDC
0EC8
0E09
0D7E
0DF6
0EF5
0F19
0DFA
0D04
0D91
0E8C
0D49
08FA
0420
01C0
021C
0323
0379
037C
034A
017A
FCF8
F76C
F41A
F444
F5D6
F632
F530
F47B
F4EA
F5B3
F5F3
F5C3
F59D
F5A3
F5E0
F6A0
F7E9
F900
F917
F876
F831
F89E
F8E8
F877
F7FA
F85A
F93B
F977
F8C7
F818
F838
F8DB
F938
F919
F8E5
F8E7
F8FD
F8ED
F88F
F7AA
F654
F568
F5C6
F6DE
F6F3
F591
F4EC
F7A5
FD5E
02A6
04A7
03F8
0331
037F
03D5
034A
02B5
0338
043F
0443
032B
02CD
04CE
08BD
0CA0
0ED9
0F3D
0EA8
0E17
0E1B
0EA5
0F1D
0EF2
0E4D
0DEC
0E2D
0E9E
0EB9
0E9A
0E8E
0E65
0DCA
0D2D
0D7D
0EAA
0F12
0D1C
0930
0567
034E
029E
026A
0291
032A
0318
0082
FB35
F5AF
F2F7
F3A0
F57D
F649
F5CF
F54C
F571
F5C5
F5BE
F584
F580
F5B9
F605
F682
F755
F82B
F869
F80F
F7E1
F872
F950
F993
F90C
F87A
F88B
F910
F956
F911
F8A0
F886
F8C9
F8FE
F8CC
F859
F81E
F860
F8B5
F84B
F6F0
F5A9
F5A3
F696
F6E7
F5E0
F542
F7A4
FD2F
02CE
0537
0449
02C2
02D0
03F3
0476
03F4
0373
038A
038F
02EA
0265
0398
071E
0BBD
0F58
10A1
0FEE
0EB0
0E33
0EB0
0F5A
0F65
0EF1
0EAD
0EC1
0E99
0DF6
0D7A
0DBF
0E5A
0E63
0DE4
0DE7
0EDD
0F99
0E5C
0AD5
0670
02E7
0113
0112
027F
03F4
0346
FF63
F9CE
F580
F41A
F4B8
F580
F5AE
F5A0
F59A
F56C
F533
F57D
F63E
F68A
F5E0
F536
F5DD
F7A2
F8F4
F8E9
F844
F83E
F8DC
F922
F8A9
F836
F88E
F967
F9E8
F9CA
F976
F93E
F913
F8D8
F89E
F87D
F877
F895
F8C9
F8AD
F7CB
F65C
F571
F5CA
F6AB
F697
F57C
F578
F8A3
FE4A
032E
04BD
038F
0245
0276
035B
037C
02CD
0281
0325
03CB
0366
0289
031E
0656
0B19
0EDC
0FF2
0EF6
0DDE
0DF1
0ECD
0F59
0F3B
0F0E
0F4C
0F7B
0EE4
0DBB
0D17
0D99
0E8E
0EDA
0E6D
0E49
0EF6
0F77
0E38
0AE1
06BF
0383
0200
021B
032C
03F0
02BC
FEB7
F919
F49C
F328
F435
F5AE
F629
F5DD
F592
F57F
F571
F56B
F592
F5C2
F5C5
F5D9
F67B
F795
F862
F858
F7E7
F7ED
F89A
F940
F946
F8DF
F8A4
F8D7
F948
F9B9
F9F3
F9D5
F97D
F943
F943
F933
F8E1
F8A0
F8C3
F8D1
F7EB
F638
F53C
F603
F762
F740
F5B9
F5BC
F995
FFB1
03F9
0449
026D
018B
0280
03A2
0377
0285
0233
02C5
0347
030E
02B9
039D
0679
0A98
0E18
0F5A
0E84
0D6A
0D9B
0EC0
0F50
0EB0
0DEE
0E2E
0F02
0F12
0E28
0D96
0E3F
0F3B
0F1C
0DF7
0D47
0DE6
0EE6
0E8D
0C06
07EE
03C6
012E
011F
030A
049A
0340
FE8F
F8E4
F53F
F491
F56A
F5EC
F586
F4DA
F4AB
F525
F5EC
F676
F65A
F5A4
F4ED
F4F3
F5EB
F75D
F8A9
F983
F9D8
F998
F8DF
F827
F7F8
F859
F8E1
F93F
F979
F99E
F986
F921
F8C7
F8E3
F949
F968
F91A
F8ED
F935
F954
F871
F6D6
F5D2
F605
F66D
F5D1
F4E1
F5FC
FA64
0033
03ED
0403
0237
0162
0261
03B5
03CB
02E5
0278
0325
0401
03DC
02F1
02EF
054F
09AC
0DD8
0FB5
0F14
0DAF
0D4E
0E23
0F0B
0F23
0EBB
0E9E
0EE1
0EF0
0E90
0E44
0E7F
0EE4
0ECE
0E42
0DF2
0E4F
0ED6
0E60
0C0C
0801
03AC
0118
017D
03CB
04FE
0294
FD10
F79E
F4F7
F510
F5EA
F617
F5B9
F573
F54F
F510
F4DD
F512
F583
F5A0
F55C
F569
F64E
F7A3
F896
F8DD
F8CD
F8BF
F8CE
F8F6
F922
F913
F8A6
F82E
F838
F8D1
F954
F939
F8D4
F8DB
F943
F949
F8B5
F84F
F8B2
F932
F8B5
F75F
F677
F698
F6C8
F604
F535
F69A
FB0F
008C
03FB
0437
02DF
0238
02F1
03FB
0424
0375
02EE
033D
03EC
03F9
0334
02E3
04A1
0894
0CE3
0F4D
0F47
0E4C
0E11
0EC4
0F52
0F0B
0E70
0E53
0EAE
0EC2
0E2F
0D72
0D3A
0D90
0DE5
0DE2
0DC6
0DFC
0E76
0E67
0CC1
0921
048D
0137
00D9
02D2
0428
020B
FCAC
F732
F4A0
F50A
F623
F61D
F558
F52F
F5ED
F699
F674
F5E1
F5A2
F5C9
F5E2
F5D5
F610
F6E4
F816
F917
F974
F920
F877
F80F
F844
F8DD
F948
F945
F92E
F968
F9B8
F997
F910
F8C2
F8ED
F914
F8DD
F8AF
F901
F95F
F8E9
F7A7
F6A0
F665
F646
F5A2
F583
F7C8
FC8E
0163
03B6
0378
02A6
02AC
0326
0321
029F
026F
02FA
03C2
03FB
0356
024A
01FE
03C3
07D8
0C91
0F60
0F45
0DDE
0D7C
0E89
0F7F
0F2A
0E21
0DB1
0E1A
0E81
0E63
0E31
0E5A
0E79
0DF7
0D1C
0CDB
0DAC
0EF3
0F5F
0DBE
09CB
04D4
015B
0124
032C
0400
00F8
FB12
F608
F46B
F551
F621
F5BB
F517
F548
F602
F65F
F636
F603
F5EA
F591
F4F7
F4CE
F5A1
F715
F856
F8F2
F8F8
F8A3
F84F
F869
F900
F979
F93B
F890
F86A
F90F
F99D
F93E
F877
F874
F93B
F99D
F91B
F8C2
F970
FA30
F96F
F766
F5FF
F634
F6C7
F661
F618
F85D
FD79
028E
04AB
03EF
02BC
0299
0317
0345
0312
02F9
0324
0366
0393
036B
02B3
01F0
02C2
0668
0BBE
0FA2
101B
0E69
0D4C
0DD8
0ED0
0ED6
0E1F
0DC2
0E2A
0EBC
0EDA
0E89
0E39
0E33
0E71
0EB5
0EB0
0E6C
0E6D
0ECC
0E3D
0B0F
05C7
01A8
0170
03CD
0450
004A
F9D2
F54D
F49B
F5BD
F604
F530
F4BE
F54F
F5F2
F5BD
F4F7
F476
F495
F514
F5A2
F620
F68E
F6FF
F791
F836
F89D
F89A
F88A
F8F2
F997
F99D
F8C6
F80F
F87A
F994
F9EB
F8FC
F7EE
F811
F926
F9CD
F96C
F8E0
F913
F9A7
F990
F88A
F743
F63C
F555
F4B9
F58F
F8E4
FE07
0298
049B
042D
030D
02B6
0344
03E3
03DC
0340
02C4
030B
03D8
0413
02FA
0178
01D1
0567
0AE2
0F1F
1024
0EC8
0D51
0D11
0DBC
0E7B
0EDD
0ECF
0E65
0DEF
0DE0
0E50
0EC5
0ED6
0EBA
0EDB
0F07
0ECB
0E5D
0E3A
0DAE
0B12
0655
0243
01C2
03EC
0466
003D
F975
F4C8
F457
F5E6
F657
F54C
F48D
F505
F5CB
F5DD
F565
F516
F51B
F52F
F546
F5A8
F685
F7AF
F8CA
F986
F9A4
F91E
F864
F81D
F873
F8F0
F929
F930
F937
F92C
F90B
F912
F944
F925
F87C
F7F5
F861
F979
F9F6
F926
F7BB
F6B2
F5FC
F529
F517
F796
FCCD
0215
0473
03BC
025E
025C
0371
0429
03E2
0335
02E8
0319
0363
035D
02FB
02D2
0408
074E
0BA5
0ECA
0F68
0E78
0DED
0E5B
0EB7
0E29
0D4E
0D4F
0E45
0F15
0EDF
0E0F
0DBA
0E35
0EC0
0EA5
0E3B
0E57
0ED6
0E2A
0AE8
05E0
0202
0162
028B
01C1
FD45
F775
F41D
F456
F5E4
F65A
F5A2
F525
F56F
F5B4
F565
F517
F56C
F5FA
F5EE
F56A
F567
F662
F7BB
F892
F8B9
F8A7
F8C7
F915
F952
F96C
F987
F9AF
F9AD
F951
F8D8
F8C6
F94D
F9EA
F9E3
F921
F861
F855
F8BE
F8C8
F825
F746
F683
F5C3
F564
F6A5
FA5A
FF68
034A
0464
0372
0272
028B
0340
038C
0327
0297
0279
02E7
036C
035B
02A1
025C
0429
0846
0CCC
0F4A
0F26
0DF2
0D8A
0E42
0F16
0F31
0EC5
0E78
0E6C
0E40
0DCF
0D7E
0DA4
0DF7
0DDD
0D5A
0D57
0E87
0FE2
0EE8
0A6D
04C3
01CE
0282
036F
00B1
FA99
F530
F374
F45B
F511
F4C3
F4D9
F601
F6EB
F666
F54D
F530
F601
F65C
F5B7
F512
F576
F6B5
F7EE
F8A4
F8E4
F8DA
F8B0
F8B6
F91F
F998
F98C
F906
F8BF
F91A
F992
F98F
F93A
F914
F92E
F95B
F9A0
F9F3
F9EB
F936
F820
F71A
F60D
F4DC
F48E
F6F0
FC46
01F4
04B2
0413
02C2
02F1
03EC
03E5
02D7
024E
02EE
03B8
03BA
032F
02B7
026C
028A
0426
0805
0CD4
0FD5
0FDF
0EB1
0E94
0F8B
0FDF
0EE7
0DE4
0E0E
0EEC
0F26
0E57
0D6E
0D4C
0DA1
0D92
0D22
0D4E
0E7E
0F4E
0DB0
0963
04D2
02CE
033F
02CF
FEA2
F809
F35A
F30A
F51F
F608
F4E1
F3B2
F41D
F566
F5FB
F5BD
F5B7
F636
F65C
F5AF
F519
F5AE
F72A
F859
F8AA
F897
F8A7
F8C6
F8B0
F878
F863
F889
F8BF
F8DE
F8F7
F93E
F9B7
FA0E
F9F6
F994
F961
F996
F9E1
F9B9
F901
F808
F6F9
F5BE
F4CB
F595
F93D
FEA4
02E1
0414
032D
0267
02B4
0359
039B
039D
03A7
0380
0309
02CF
0335
0387
02FC
028D
0475
092F
0E14
1018
0F35
0E06
0E62
0F8D
0FEC
0F55
0EEA
0F45
0FA6
0F2D
0E28
0D9F
0DE6
0E3D
0DED
0D49
0D48
0E2A
0EA6
0CE8
08C5
0490
02BA
02AD
0126
FC50
F66E
F367
F43A
F62A
F669
F53C
F4B6
F569
F5D8
F512
F436
F497
F5B5
F61C
F590
F537
F5D7
F70C
F825
F8F1
F963
F940
F882
F7CB
F7D1
F873
F8D9
F897
F83B
F86F
F90F
F97A
F96D
F92A
F8F7
F8F6
F937
F994
F9AA
F930
F830
F6CA
F54A
F4A9
F65C
FAE1
0083
0453
04CA
0334
020C
024A
02ED
02F3
02A4
02B3
031A
037A
03CB
03EC
0350
0217
01FD
04E3
0A31
0EBE
1006
0ED5
0DF8
0EAB
0F84
0F11
0E20
0E6A
0FDD
1099
0F8E
0DEA
0D7B
0E6F
0F40
0EBF
0D97
0D6C
0E84
0EFD
0CCE
0855
0429
0225
012C
FEA6
F9F7
F5A6
F465
F5C0
F6CC
F5F6
F4AF
F4DC
F613
F675
F57F
F493
F4CF
F599
F5D0
F574
F57B
F64C
F756
F813
F8B2
F958
F994
F914
F85F
F832
F874
F877
F819
F7E8
F839
F8AB
F8C6
F8AF
F8E3
F970
F9CD
F98E
F905
F8CF
F8DF
F855
F6AB
F4DE
F510
F892
FE2D
02C6
0436
0355
02B1
036B
043F
03CA
02A3
0256
0319
03A4
0334
028B
0290
02E3
02C7
02FB
0545
09D1
0E3C
0FFB
0F34
0E2D
0E68
0F41
0F67
0EAE
0DFE
0DFC
0E5E
0E91
0E8B
0EAE
0EFC
0EEB
0E37
0D78
0D92
0E6E
0E9F
0CAD
08CC
04DA
0234
FFFE
FC67
F788
F3E1
F376
F54B
F6A7
F649
F55A
F54C
F5E7
F5F9
F548
F4D1
F53C
F5F5
F621
F5C6
F589
F5CD
F695
F7CF
F926
F9DB
F97A
F88E
F81F
F86D
F8BA
F870
F7FA
F81E
F8C9
F920
F8BF
F855
F89A
F943
F97D
F931
F91E
F99B
F9D3
F8A4
F63B
F48C
F5D4
FA67
0007
03C7
04A0
03F6
039C
03EB
040D
03A0
0343
036E
039B
032B
029C
02E8
03CA
03D3
02B6
0276
0537
0A4A
0E8C
0FBC
0EBA
0E00
0EA2
0F89
0F67
0E74
0DDC
0E10
0E68
0E55
0E30
0E89
0F26
0F30
0E5C
0D84
0DB2
0E9B
0E89
0C2F
0848
04B2
0208
FF03
FAA2
F61B
F3C5
F444
F5BD
F61E
F567
F507
F584
F5DF
F560
F4C9
F526
F626
F691
F5FB
F535
F52A
F5EF
F715
F837
F901
F91D
F88C
F7ED
F7E0
F83E
F853
F7FF
F7F2
F88F
F927
F8F4
F850
F844
F908
F9A9
F959
F887
F840
F8B1
F8CC
F79E
F5CE
F568
F803
FD0F
0210
049B
045D
031F
02CF
0392
0420
03BC
0322
033D
03C3
03B9
02EF
023A
022A
0269
02B9
03ED
06FB
0B2E
0E52
0EFE
0E2A
0DDD
0EC1
0FBB
0FBF
0F1B
0EBE
0ED7
0EDB
0E9A
0E88
0EE5
0F1C
0E97
0DCB
0DD4
0EEE
0FC9
0ED3
0BDA
080A
0469
00D0
FCAF
F866
F55C
F48D
F55F
F632
F5FC
F51D
F499
F4D0
F53A
F532
F4C4
F494
F519
F610
F6B9
F6A4
F632
F62B
F6E5
F7EB
F88E
F8A1
F886
F88B
F88A
F844
F7E3
F7DF
F856
F8D7
F8ED
F8B6
F8AC
F902
F966
F961
F8E7
F867
F854
F878
F806
F6A0
F56C
F67F
FAC9
008B
0483
04F6
0348
022D
02B0
03A2
03C7
036F
0378
03B9
036A
02B2
02A5
0379
03D9
02BF
0177
029A
06ED
0C1A
0F19
0F36
0E2E
0DC5
0E2A
0E97
0EA6
0E8B
0E83
0E88
0E8E
0EB1
0EFB
0F34
0F1D
0EC9
0E90
0EB3
0F12
0F25
0E2F
0BB4
07DA
0344
FE88
F9FF
F63F
F433
F44C
F5A8
F693
F61F
F4FB
F471
F4CB
F525
F4CD
F437
F44A
F51A
F5E2
F60E
F5E9
F617
F6CF
F7B3
F854
F894
F89F
F8A8
F8C6
F8E3
F8D7
F8A4
F891
F8DC
F950
F967
F904
F8C1
F925
F9C4
F9A1
F883
F77A
F797
F86B
F870
F731
F666
F84B
FCF8
01F0
0482
044C
031F
02BE
0340
03AA
0387
034D
0375
03C1
03AD
034D
0337
0396
03C5
032F
0275
033B
0671
0AFD
0E7D
0F77
0E98
0DB0
0DB9
0E32
0E4C
0E1F
0E50
0EED
0F36
0EBB
0E17
0E28
0ECF
0F0F
0E6D
0DAA
0DDC
0EE2
0F2A
0D05
0821
01BA
FBA5
F73C
F4FA
F489
F50E
F58E
F56E
F4C3
F42A
F437
F4E3
F580
F56E
F4DB
F499
F522
F5FD
F64C
F5F0
F5C1
F691
F828
F983
F9FF
F9EB
F9F1
FA33
FA5F
FA58
FA67
FAB9
FAFA
FAB0
F9EE
F974
F9E6
FAED
FB54
FA67
F902
F8D0
FA44
FBA7
FADE
F830
F6AB
F920
FEE3
043A
062D
0539
040A
043E
0530
058F
0526
049F
0454
03F1
034A
02D1
0305
03C1
0465
047C
0411
03AD
0425
0624
096D
0CAF
0E86
0EB3
0E27
0DDD
0DF3
0DF2
0DB0
0D88
0DD1
0E5A
0EB5
0EAE
0E72
0E49
0E58
0E78
0E4E
0DCA
0D80
0E07
0EA8
0D29
07CE
FFA4
F842
F4B6
F4D4
F5E7
F5CF
F4D1
F452
F4B3
F51C
F4FD
F4D8
F55C
F65B
F709
F701
F698
F62E
F5B6
F513
F4A7
F520
F6AE
F8AB
FA21
FA92
FA44
F9E1
F9E3
FA38
FA75
FA4E
F9ED
F9B5
F9CB
F9F8
FA01
F9F3
F9E6
F9B0
F939
F8F9
F9A5
FAFD
FB8A
FA2F
F801
F7BC
FAFF
0043
0440
0535
0441
038A
03D8
0479
04B7
049D
046B
0416
0396
033B
0348
0391
03CC
0411
0485
04C0
044F
03F2
0553
08E8
0CCF
0E9A
0E04
0D04
0D49
0E70
0F01
0E87
0DEA
0DF7
0E6C
0E9D
0E62
0DFD
0DA7
0D8C
0DB9
0DCC
0D47
0C93
0CDB
0E07
0D8E
089C
FFCF
F79C
F422
F4FE
F65D
F5C0
F453
F445
F57A
F624
F59D
F50A
F556
F5E7
F5DB
F577
F5A1
F65C
F6A4
F5EC
F4FE
F50E
F66E
F870
FA24
FAE2
FA8D
F9CB
F9A5
FA53
FAD9
FA41
F902
F87A
F91F
F9F1
F9E6
F959
F95C
FA09
FA6E
FA1A
F9D1
FA25
FA51
F962
F823
F8B4
FC0C
0098
03C3
0477
03CC
0367
03D3
0476
04A3
0451
03F6
0407
0492
051D
050D
0454
03A2
039C
03FB
03E6
0339
0320
04F9
08B6
0C9C
0ECF
0EF5
0E38
0DD9
0E0C
0E33
0DEA
0D8B
0DAD
0E4E
0EAC
0E17
0CDE
0C39
0CF3
0E53
0EB5
0D9C
0C97
0D6C
0F44
0E94
08AB
FF1E
F6DB
F384
F444
F593
F569
F4B1
F4E1
F5AD
F5CE
F52C
F4F0
F5A8
F660
F60D
F509
F490
F513
F5CC
F5F9
F5C2
F5BC
F623
F6F1
F82E
F99A
FA7D
FA60
F9C2
F987
F9E1
FA38
FA1F
F9CF
F98F
F931
F8A6
F894
F981
FAA4
FA9C
F974
F8E3
F9D2
FAC0
F9C9
F7BA
F7B5
FB71
00F1
04A6
0532
042D
03A2
03E7
0441
0468
0499
04C3
04A5
046E
0476
047E
03F9
0320
02FD
03ED
04D3
0475
0381
0437
07BF
0C76
0F7F
0FB3
0E71
0DAE
0DF0
0E4F
0DF9
0D25
0CAE
0D08
0DC1
0E14
0DCE
0D88
0DDA
0E7C
0E79
0D7F
0CA7
0D47
0EBF
0E21
08D3
FFBC
F722
F2F9
F372
F57A
F636
F57A
F4D2
F512
F598
F5A6
F57B
F5A5
F5ED
F5AA
F4F6
F4BB
F553
F5D3
F538
F3FA
F3B1
F537
F7A2
F95B
F9C6
F98A
F976
F9A7
F9D3
F9EC
FA0E
FA20
F9D5
F92F
F89E
F89B
F931
F9DE
FA05
F99E
F95D
F9DA
FA95
FA6A
F935
F8A4
FAA0
FEE6
02D8
042A
0347
026D
02C9
0384
03A5
03A3
0457
054C
054F
044E
038A
03D1
0471
0472
0418
044A
04EE
04F1
043D
0464
06C3
0A93
0DB8
0F08
0EFE
0E99
0E4F
0E25
0E1A
0E17
0DF5
0DC4
0DCA
0DFC
0DCB
0D03
0C73
0CE9
0DB6
0D72
0C6B
0CB1
0EA4
0ED1
0939
FEBB
F561
F260
F4C7
F752
F6C0
F4A9
F40A
F510
F5A5
F4E4
F424
F4AC
F5F0
F68E
F627
F56B
F4ED
F4A1
F474
F48C
F4DC
F51C
F575
F68C
F86E
FA01
FA2F
F957
F8DD
F961
FA21
FA34
F9AD
F93C
F915
F8F4
F8ED
F96D
FA59
FAE1
FA9C
FA27
FA1E
FA1B
F98F
F940
FAE3
FED3
0307
0504
047D
0345
02DE
030D
0305
02ED
036B
045A
04F1
04F0
04D3
04C0
043D
0343
02D8
03D1
0540
055D
0414
03B9
0660
0B1E
0EDB
0F99
0E36
0CFD
0D26
0E16
0E90
0E2A
0D8A
0D73
0DD3
0DE0
0D19
0C26
0C43
0D8F
0E7A
0DB9
0C73
0D01
0F21
0EE4
08D9
FEB1
F631
F353
F49F
F5E5
F557
F486
F500
F5EF
F5D0
F4E7
F49A
F52D
F58A
F518
F48A
F4A5
F521
F53F
F4DE
F470
F441
F465
F528
F6C3
F887
F94B
F8FB
F8E5
F9E2
FB07
FAFB
F9E7
F91B
F924
F94C
F912
F911
F9CD
FA89
FA43
F96B
F95C
FA15
FA12
F8FB
F907
FC44
0159
04AA
0495
0315
02D0
03D2
0443
0384
02F4
0396
048A
049D
0431
0461
050C
0507
0419
0370
03CD
044D
03C7
02D4
036F
0686
0AB5
0DB4
0E95
0E16
0D65
0D1D
0D30
0D3F
0D05
0CD2
0D43
0E56
0EFB
0E45
0CD9
0C73
0DA0
0ED2
0E7B
0D6B
0DB6
0F09
0DCA
0721
FD1A
F533
F2E1
F486
F628
F5E8
F4F5
F4DD
F56A
F588
F50A
F4A5
F4B7
F4F6
F51C
F529
F513
F4C2
F46E
F47A
F4E2
F528
F51F
F55C
F680
F82E
F95D
F9A6
F9AF
FA13
FA8D
FA8E
FA2C
F9DA
F9A5
F94E
F8ED
F8DD
F90B
F8FA
F8B1
F8DF
F9AE
FA05
F90F
F833
FA1F
FF45
0491
068E
0538
0378
0348
03C4
0353
0253
026B
03E0
0513
04D4
03F8
03D7
0444
0424
0373
0362
0462
0530
0475
02CD
0267
04AE
08C2
0C6D
0E37
0E56
0DFE
0E19
0E91
0EA1
0DE7
0D12
0D16
0DC7
0DED
0D17
0C80
0D65
0EE5
0ED2
0CEB
0BED
0E08
10EC
0F3C
06A6
FB50
F3E7
F2EE
F523
F61F
F508
F40B
F49E
F5BD
F5C6
F4BA
F3EB
F429
F50B
F5CB
F60B
F5D9
F56D
F519
F50E
F517
F4DA
F46E
F482
F5AC
F7A9
F97F
FA55
FA10
F933
F872
F85D
F903
F9BF
F9D3
F957
F927
F9A2
FA01
F976
F885
F864
F90E
F912
F7EE
F7C1
FB2A
0181
069C
0735
0488
0289
0324
0496
0486
0328
0278
0336
0416
03EC
034E
036A
0425
046A
03ED
0391
03FC
048F
043B
0313
029E
047A
08AB
0D3D
0FA7
0EEE
0CA3
0B87
0CCB
0EDD
0F66
0E33
0D40
0DC4
0E82
0DCF
0C49
0C13
0D98
0EB9
0DF8
0CF0
0DFF
0FE2
0DF8
05D3
FB08
F3EB
F306
F547
F669
F57E
F478
F4A5
F539
F525
F4C3
F4FD
F5B2
F601
F5A3
F536
F535
F56D
F589
F58E
F586
F542
F4BA
F474
F51A
F6A1
F831
F8FF
F905
F8CF
F8D6
F941
F9E2
FA3E
F9E9
F921
F8B7
F914
F99C
F989
F91E
F949
FA0F
FA2D
F90C
F86E
FAF7
00A5
05ED
0732
04A5
01D2
0199
037F
0511
04F0
03D1
0302
02E2
030D
034A
03B7
043F
047D
0437
03A0
031F
02F3
030A
0336
03AB
051D
0810
0BC8
0E7B
0EFD
0E0D
0D7E
0DFF
0E6B
0DAA
0C87
0CB1
0E2E
0F1C
0E50
0CF1
0CA4
0D1D
0CE2
0C0A
0C71
0E89
0F5A
0B4A
02A1
F9E0
F530
F49F
F562
F587
F538
F51D
F51C
F4F5
F4F2
F563
F5F9
F640
F64A
F65C
F631
F566
F490
F4CF
F5F8
F64B
F4C7
F2E5
F2FF
F55F
F809
F954
F994
F9D1
F9F8
F953
F834
F7DE
F8A2
F961
F94E
F907
F931
F921
F838
F7AA
F927
FBC5
FC37
F958
F718
FAB3
03F3
0C34
0D31
07BA
022B
0120
0359
04CF
03EB
027E
0277
035A
036C
0241
0143
01C9
037A
04D6
04F1
045F
045C
0531
059C
044A
01DA
00E8
0381
08CE
0DAF
0FBA
0F39
0E2B
0DDA
0DFC
0DE4
0DB1
0DD8
0E23
0DEB
0D2F
0CC2
0D2B
0DCC
0D8F
0C62
0B9B
0C7A
0E2E
0DE0
093A
0111
F922
F4DB
F467
F52A
F4FA
F438
F47C
F5EC
F6FB
F6BA
F61F
F670
F743
F71A
F59F
F432
F40A
F4A8
F4D5
F469
F445
F4AD
F4E4
F49D
F4BC
F607
F7EC
F94D
F9F8
FA6B
FA82
F98E
F7E2
F71B
F81D
F995
F99E
F879
F824
F94A
FA42
F9D2
F949
FA4A
FBB4
FB01
F8CC
F985
000C
08EB
0D28
09F7
03A9
004D
0137
0332
039A
0309
0313
03A5
03AA
0322
0315
03CC
0452
03ED
0326
02DE
032C
03A7
042A
048A
0435
032F
02FF
056C
0A09
0E08
0F24
0E1E
0D87
0E72
0F5D
0EB0
0D00
0C1E
0C90
0D37
0D42
0D31
0DA1
0DF6
0D2D
0BAF
0B4F
0CEA
0E80
0C86
0594
FC56
F573
F370
F4D5
F633
F5B4
F461
F42E
F568
F6A0
F6AA
F5D7
F524
F4F4
F504
F51C
F526
F4F2
F477
F441
F4EF
F624
F690
F59F
F491
F517
F713
F8BF
F920
F924
F9C1
FA47
F98B
F801
F754
F808
F8CD
F897
F832
F8D0
F9F8
FA5B
FA2F
FAC9
FBB2
FA91
F74E
F64C
FBDB
05F5
0D18
0C48
066B
023F
0265
03B3
02E9
0119
0132
0358
0507
04DE
0408
03D2
03D7
0344
0289
029C
0350
039B
0352
033E
0377
0322
0274
0375
076A
0C62
0F0D
0EB8
0DE4
0EA9
100B
0FD0
0DF1
0CA7
0D33
0E3C
0E04
0CFA
0CC7
0D93
0DD0
0CCE
0C0B
0D0E
0EB3
0DA9
07F4
FF67
F82B
F4E9
F4CD
F535
F4BC
F416
F45E
F563
F5FC
F5A7
F51A
F50D
F522
F4AA
F408
F45B
F5A9
F67F
F5E3
F4C9
F4C1
F5C0
F646
F5A1
F505
F5E1
F7DC
F95B
F9A6
F96C
F942
F8D5
F80B
F7B1
F855
F943
F997
F99E
FA17
FA94
F9FD
F8B9
F8C4
FAA8
FBDD
FA14
F78B
F988
0192
0A53
0D11
0915
03C0
01D5
02F1
03ED
0384
02ED
02FE
030C
02B2
02CC
03C2
0461
03A5
028C
02BD
03F5
0473
03AD
02FA
0340
0391
031F
0366
0686
0BB0
0F29
0ECA
0CCD
0CCA
0EFF
1074
0F5D
0D6E
0D2F
0E80
0F2B
0E25
0CD4
0CC8
0D8A
0D9C
0CF0
0CF4
0E25
0E93
0B8D
0488
FC0E
F5C1
F370
F3FE
F4EB
F4CD
F41C
F3F2
F48A
F536
F55D
F517
F4CE
F4B1
F4B5
F4E4
F52E
F531
F4AF
F433
F494
F597
F5EC
F4EE
F3D7
F466
F6B3
F907
F9EC
F9A8
F965
F98D
F9A1
F964
F92C
F913
F8C7
F861
F88D
F961
F9E7
F996
F960
FA33
FAF0
F994
F6CB
F6C2
FCAC
0609
0C3A
0B55
060C
0213
01E5
037B
0421
038D
02F7
02D7
02BA
0291
02E8
03BC
0440
040D
03AF
03AB
03A7
0341
02F6
0354
03D6
03A5
0368
050C
0923
0D79
0F3D
0E4A
0D2F
0DDC
0F68
0FCC
0ECA
0DF9
0E41
0EB6
0E46
0D64
0D45
0DF0
0E23
0D4C
0CA5
0D91
0F1A
0E22
0883
FFAD
F7B2
F3BD
F3A7
F4D4
F50D
F434
F387
F3CC
F4A9
F569
F5B1
F57C
F4E5
F446
F427
F4A4
F522
F4F8
F478
F4AB
F5DF
F6EC
F68B
F526
F48A
F5B9
F7BC
F8FE
F928
F909
F929
F93D
F8F8
F8A1
F889
F889
F880
F8D0
F9B1
FA5E
F9F3
F902
F911
FA1B
FA0E
F7EA
F681
FA00
0275
0A6C
0C4D
0855
03CD
02A8
03BB
03C4
0240
0182
02D1
048C
0494
0319
0203
024E
0323
0365
031F
02FB
032A
0362
0371
0343
02CE
0290
03C5
072B
0BA2
0ECB
0F74
0EC5
0EA2
0F4D
0F7B
0E82
0D6D
0D74
0E3A
0E78
0DF7
0DC8
0E66
0EC8
0DEB
0CB5
0D18
0F24
0FD2
0BB7
02DE
F95E
F3B8
F2F1
F46B
F521
F46B
F3A6
F3F4
F4F3
F583
F537
F488
F41B
F43F
F4F4
F5E1
F645
F592
F457
F3EB
F4D6
F5F9
F5EB
F4F5
F4D8
F671
F872
F926
F8BE
F8D3
F9C5
FA25
F911
F7D8
F831
F9B4
FA73
F9BB
F8DB
F8EA
F93E
F8FD
F8FF
FA58
FBAD
FA6B
F74A
F736
FDAC
0759
0CC5
0A76
047C
012E
0228
0408
03FB
02FB
0324
0439
0465
0357
0296
031A
0404
0416
0342
025F
020C
0267
034B
041D
03EB
02AB
0241
04E9
0A30
0EA9
0FA1
0E2F
0D79
0E96
0FA1
0EE0
0D36
0CA6
0D7C
0E32
0DFE
0DE2
0EBB
0F7D
0E9E
0CAE
0C0D
0DC0
0F87
0DCD
0748
FE62
F719
F3B2
F377
F444
F4BC
F4D8
F4E1
F4B0
F41B
F3AA
F421
F55C
F61E
F58E
F46E
F42A
F4DD
F53C
F49C
F3FE
F46E
F559
F567
F49F
F48A
F614
F83D
F97B
F9A7
F9B4
F9F0
F9CE
F956
F96C
FA3D
FAAA
FA0C
F957
F981
F9C5
F8EB
F7CD
F891
FB06
FBE0
F94B
F6E9
FA67
03E1
0C56
0D3D
07CB
02B4
01FD
0396
03D0
0265
01A5
026B
0333
02E6
026D
02D7
0383
0356
02A7
0298
033D
03BA
03D1
03FC
041B
0371
0262
02FC
06A9
0BDC
0F51
0FAE
0EC2
0EC2
0F85
0F6D
0E23
0D00
0D04
0DA4
0DE9
0DC0
0DBA
0DF9
0E00
0D97
0D55
0DD7
0E96
0DC5
09A7
0242
F9FB
F43A
F2C4
F423
F531
F461
F2EB
F2AC
F3CD
F515
F5C6
F61D
F63A
F5B7
F4A2
F403
F497
F58D
F57D
F47C
F406
F4AD
F53C
F4C9
F459
F563
F77E
F8E9
F913
F935
FA25
FAEB
FA44
F8BE
F805
F885
F912
F914
F953
FA2C
FA8D
F9DA
F967
FA6A
FB68
F9F9
F73C
F811
FF4A
08EF
0DA0
0AB0
04BE
01C2
0289
03A2
02F8
01F1
0255
0392
0407
038D
0348
039C
03B9
032F
02AB
02B7
02D7
02A1
02BA
03B8
04B5
0471
03B2
04F4
0936
0E1A
1046
0F2E
0D82
0DB3
0F30
0FBC
0EAB
0D9B
0DF8
0F0C
0F18
0DB1
0C33
0BF6
0CCA
0D9C
0E05
0E64
0E47
0BCF
0597
FD1D
F632
F382
F42E
F531
F4CA
F3C0
F381
F411
F486
F4BE
F564
F651
F64A
F4E2
F39F
F42E
F5FB
F6C2
F585
F3CF
F38D
F486
F4FF
F47B
F480
F651
F8E9
FA2D
F98A
F872
F86D
F979
FA7F
FAA9
F9FD
F8FD
F834
F7F3
F81C
F83E
F844
F8CD
FA34
FB5B
FA84
F809
F752
FBAA
0405
0B09
0C1D
07F0
0355
0208
0390
051F
0537
047F
03D5
031F
0230
01BA
026F
03BF
044B
039F
02B5
0299
032A
039D
03AD
03AD
03C8
03FF
04DB
0739
0AEE
0E2F
0F3D
0E66
0D90
0DD1
0E59
0E24
0DA6
0DF5
0ED6
0EEE
0DE4
0D19
0D94
0E49
0DA0
0C3B
0C7B
0EBC
0F94
0B41
024F
F97F
F4E6
F457
F4D3
F471
F3B1
F39D
F3FD
F40C
F3E6
F44E
F548
F5E0
F577
F49E
F461
F4FE
F59D
F54E
F426
F34A
F3B5
F51E
F646
F663
F5FA
F625
F736
F865
F8DE
F8C7
F8CD
F915
F92D
F8FE
F8FD
F94A
F977
F970
F9C1
FA78
FA92
F976
F86F
F948
FB58
FB87
F885
F5E6
F8D1
017A
09E0
0C1C
0872
03EF
0247
02FD
03FF
04A2
052E
0529
03E5
023E
0201
0359
045D
03D4
02EA
0330
0426
0438
0361
0313
03C0
0411
0330
0288
042E
080D
0BE6
0E07
0EBB
0EE5
0E94
0DC1
0D41
0DC5
0E98
0E8E
0DD5
0D9D
0E36
0E9C
0E2E
0DA6
0DCE
0E06
0D4C
0C39
0C5A
0D2E
0B80
050E
FBFC
F517
F302
F42B
F553
F4F2
F3DA
F36A
F403
F4FE
F595
F581
F513
F4CB
F4C2
F47D
F3B7
F32F
F3E5
F57C
F660
F5DB
F505
F4FC
F54D
F50B
F4B8
F5B9
F808
F9C7
F99F
F889
F840
F8C5
F8C3
F829
F85F
F9AA
FA54
F95E
F844
F8A9
F9AA
F977
F892
F915
FAC6
FA9F
F7C6
F6B1
FC3E
0636
0C61
0A24
0401
0170
03C0
061D
054C
037E
03CE
0563
0548
0361
028F
040E
058F
04E0
032F
02E9
0402
0496
042D
0410
049A
047F
0359
032C
0602
0AD4
0E65
0F16
0E65
0E5E
0EEE
0EC7
0DC8
0D11
0D2D
0D8E
0DB7
0DE0
0E55
0EE5
0F20
0EBA
0DB7
0C98
0C5C
0DA0
0F3A
0E46
08B0
FFEC
F848
F4DF
F4F1
F58A
F502
F3F7
F394
F416
F4EB
F565
F521
F43C
F361
F352
F41F
F504
F54D
F523
F527
F564
F55C
F508
F4EC
F512
F4EE
F4B0
F581
F7A5
F969
F90A
F734
F65D
F7AF
F9BB
FA9B
FA51
FA0F
FA04
F969
F873
F865
F940
F953
F802
F72C
F84B
F9A3
F8B3
F6E7
F907
00DF
097E
0C15
07D6
02A7
01CE
0450
05D1
04BA
0330
0317
03C4
03E1
038C
039F
0406
03FC
037B
034E
03BE
041B
03F4
03C5
03F3
03F8
0377
0368
052A
08A5
0C45
0E94
0F47
0EDE
0DFE
0D3F
0D11
0D6A
0DCA
0DCA
0D92
0D8D
0DD7
0E47
0EDC
0F71
0F40
0DDC
0C9C
0D8F
1035
1095
0B2C
0155
F86E
F47D
F4BE
F5C1
F595
F4D6
F46C
F413
F37D
F354
F416
F4F7
F4F1
F45C
F452
F4FB
F571
F52C
F4A4
F476
F4A6
F4F1
F545
F58B
F570
F4FE
F518
F684
F87E
F967
F908
F8F0
FA05
FB10
FAA7
F963
F8F0
F9A2
FA47
FA28
F9C6
F972
F89B
F761
F779
F9C6
FBE2
FAA4
F770
F817
FFA1
094B
0D42
097D
0369
00FD
0289
0462
0471
03DF
0400
043B
03CD
0377
0418
04E3
049C
039D
032C
0368
0363
02F8
0308
03BA
03EC
0300
024B
03AE
071B
0AA1
0CE3
0E31
0F02
0EE8
0DDF
0D2F
0DC6
0EA2
0E4A
0D17
0CA6
0D66
0E22
0E11
0DEC
0E5C
0E88
0D97
0CBA
0DB4
0F33
0D0E
056B
FBE8
F5DD
F497
F505
F461
F30A
F29F
F341
F3D8
F401
F452
F4E3
F4F7
F463
F412
F48C
F51C
F52A
F54C
F601
F66E
F592
F409
F363
F40B
F517
F602
F760
F962
FACF
FA75
F922
F8C3
F9B2
FA58
F9CC
F920
F94D
F98C
F8E6
F816
F851
F931
F97B
F96C
FA47
FB88
FACB
F7DF
F711
FC9C
0631
0C2F
0A62
04D8
0244
03E4
05A3
04D0
033D
036D
04AB
04B2
037E
0313
0401
0482
038D
028E
02F1
03C4
037C
02AE
02F9
0409
03F4
0289
0244
051B
09BA
0D07
0DC8
0D7F
0DCE
0E7C
0EA4
0E57
0E29
0E10
0DD4
0DD8
0E6B
0EFA
0EDF
0E72
0E4A
0DF5
0CAA
0B38
0B90
0D9F
0DD1
0897
FF35
F72B
F44C
F50A
F589
F498
F3E2
F467
F518
F4EB
F47B
F4BB
F548
F51B
F454
F41B
F4BD
F51F
F48C
F3ED
F460
F58A
F630
F5F6
F580
F558
F59B
F674
F800
F9AC
FA7C
FA25
F973
F941
F974
F96B
F91E
F90C
F943
F959
F95A
F9B9
FA11
F96C
F83C
F876
FA9B
FC0E
FA6B
F7E9
F9F1
023E
0B45
0D9C
0858
01DF
002D
02A4
04A7
0416
02D2
02E2
03CE
0435
0403
03FB
0415
03AC
02E8
02C0
036C
03F1
03AF
035B
03A5
03ED
035A
02AD
03B7
0709
0B20
0DFF
0EF3
0EAC
0E1C
0DAD
0D4B
0CD7
0C6A
0C63
0D1D
0E55
0F13
0EBA
0E09
0E34
0EF8
0ED6
0D8F
0D02
0E46
0EF0
0B16
023A
F8C1
F3A9
F399
F51E
F545
F45E
F427
F4F7
F5CC
F61A
F61D
F5D9
F506
F3F2
F376
F3DF
F485
F4C3
F4BE
F4E7
F51E
F4E7
F459
F421
F485
F523
F5E1
F747
F965
FB19
FB3F
FA17
F8E0
F865
F894
F90E
F986
F99B
F925
F8BC
F93E
FA68
FAB9
F980
F853
F907
FA8F
FA17
F7CA
F834
FEC1
0847
0D7C
0B0B
051A
01F3
02FE
04B3
045C
0335
0368
0484
04AD
03D2
038E
0462
04FA
045F
035A
0311
0358
0351
0307
0341
03F2
03FF
0327
030E
0562
0989
0D12
0E59
0DEA
0D68
0DC9
0EB7
0F47
0F03
0E61
0E21
0E52
0E40
0D8B
0CE8
0D53
0E81
0EED
0DE6
0CE7
0DA5
0EEC
0D11
064D
FD77
F749
F580
F5E6
F5B3
F482
F3A8
F3C7
F42C
F430
F414
F43F
F47E
F47A
F46B
F4AD
F524
F575
F57F
F539
F49F
F419
F45B
F564
F61F
F5BF
F515
F5AD
F79D
F920
F8F7
F82E
F897
F9F1
FA45
F904
F800
F8A0
F9C8
F9C7
F8F3
F8C8
F947
F924
F86C
F8D0
FA8E
FB1D
F8EB
F73C
FB2C
046B
0BFD
0BFA
0672
024C
02BD
04C3
04B2
0318
02B3
03D2
0449
0348
029A
037B
046E
03B0
0228
020D
0383
0492
043B
039C
03BC
03DF
0305
0232
03A4
07E1
0C9C
0F2C
0F39
0E64
0DFD
0DF9
0DD2
0D74
0D32
0D66
0E1A
0ED0
0EDF
0E43
0DB5
0DB2
0DC9
0D6A
0D19
0DE6
0F55
0EA8
096A
00B0
F8B9
F4D2
F475
F4E3
F49E
F440
F49D
F55F
F5BD
F593
F558
F558
F568
F54F
F51E
F50E
F53B
F58D
F5BB
F56D
F4BA
F45C
F4E5
F5BC
F5C9
F534
F581
F75B
F951
F9A0
F8A2
F83A
F913
F9C5
F91A
F809
F851
F9C4
FA89
F9E4
F923
F942
F96D
F8D1
F85B
F91C
FA0A
F982
F8BE
FB71
02B8
0A2B
0C0B
07F4
0337
0250
042C
0502
03DD
0304
03D7
04DB
044C
02C9
023F
032C
0444
0478
0417
03C2
0359
02A8
0232
0262
0299
0217
0193
02D5
0680
0B0F
0E39
0F06
0E3A
0D2D
0C95
0C7F
0CDB
0DAD
0EBE
0F79
0F46
0E2B
0D04
0CEE
0E07
0F08
0EA5
0D75
0D64
0ED7
0F26
0B17
02C3
FA27
F561
F4FA
F62E
F667
F590
F50B
F56B
F5F0
F5C7
F4F9
F41E
F3A4
F388
F37F
F366
F383
F42B
F531
F5FC
F646
F66A
F6B6
F6BF
F602
F504
F528
F6EB
F8E4
F95C
F889
F831
F90F
F9DD
F973
F8A5
F8EC
FA01
FA4C
F96D
F8ED
F9CA
FABB
FA1B
F8A5
F883
F9BE
F9DA
F809
F7D0
FD49
072D
0EEA
0F4C
09C9
044A
02AC
03D8
04C1
0457
03A0
035D
031F
0293
0242
02AE
0379
03E3
03C9
03A9
03D4
0402
03CA
033B
02C4
0299
0274
020B
01B8
027A
051B
0921
0CC6
0E54
0DD5
0D02
0D58
0E82
0F0F
0E77
0DC7
0E25
0F36
0F97
0EC6
0DDB
0DFA
0EAE
0E7F
0D2A
0C44
0D0F
0E22
0C44
05FD
FDBA
F7B5
F5DD
F662
F65A
F512
F410
F473
F573
F5C3
F559
F511
F521
F4D9
F3F5
F348
F39E
F49F
F555
F58D
F5EB
F6A3
F702
F687
F5BD
F570
F593
F5AA
F5E2
F6F2
F8D1
FA50
FA66
F96A
F886
F848
F859
F87A
F8E4
F985
F9BF
F966
F948
F9FD
FAAE
FA1D
F8A6
F811
F8FE
F9B9
F8D1
F833
FBCE
0475
0D5F
1049
0BE2
04F8
0134
01C1
0394
03E3
02EE
0280
0324
03C2
0393
0324
0349
03CD
03E0
0363
0321
0398
0430
0404
031D
026A
0272
02AE
0278
025E
03D7
077A
0BDD
0EB0
0EF2
0DD0
0D3B
0DEB
0EE8
0EF5
0E17
0D70
0DAF
0E31
0DF3
0D18
0CD9
0DC7
0ED5
0EAE
0DB7
0DA9
0EC0
0E45
0931
0040
F813
F4A9
F578
F6C9
F640
F4CA
F44C
F4D3
F50C
F492
F461
F4FD
F589
F539
F4A2
F4BC
F546
F537
F479
F423
F4E7
F60E
F686
F636
F5C5
F56C
F505
F500
F63B
F87A
FA1B
FA07
F928
F923
FA1D
FACA
FA7F
FA02
FA0B
FA0D
F943
F847
F855
F940
F980
F8A7
F833
F913
F9B1
F846
F6A6
F967
023D
0C87
1128
0DBE
06BB
0233
01ED
0349
03A3
030D
02E9
037F
03EF
03C1
0376
03A0
040F
0438
03F3
0389
033B
0317
0325
0366
03A9
0396
0305
0246
0214
034E
065D
0A8B
0E17
0F6D
0EA4
0D69
0D41
0DF3
0E2F
0D81
0CE8
0D4C
0E1D
0E30
0DA0
0DB7
0EDA
0F98
0EA9
0D25
0D5F
0F58
0FA2
0AF3
0247
FA4E
F693
F649
F646
F51F
F40C
F441
F4F7
F4D3
F411
F414
F526
F5E6
F54C
F42D
F416
F51F
F5EE
F5AD
F513
F51D
F596
F59C
F516
F4C9
F514
F56E
F571
F5B6
F70E
F921
FAA2
FAC9
FA17
F976
F926
F8F6
F8F4
F951
F9CA
F9D4
F978
F954
F98D
F96E
F88A
F7B3
F7F1
F8BB
F884
F792
F8F4
FF3A
085F
0E9A
0DFE
088A
03B9
02A5
03BB
041A
0365
034D
0463
0529
046D
0312
02C6
03A3
0443
03DF
0344
0361
03DF
03CE
032C
02D2
030E
0330
02BA
0269
039A
06B6
0A9D
0D8F
0E86
0DD8
0CD3
0CBE
0DC7
0ECF
0EA8
0D87
0CD2
0D48
0E16
0E2C
0DCC
0DF9
0E9E
0E86
0D7B
0D33
0EE5
107C
0DF7
0626
FCC8
F6DA
F590
F612
F5A6
F481
F434
F4D8
F515
F473
F419
F4E8
F60D
F628
F541
F495
F4CD
F551
F563
F51B
F4FD
F52A
F55F
F571
F564
F523
F4B5
F4A1
F597
F770
F90C
F998
F97E
F9A9
FA1A
FA00
F92E
F8A0
F921
FA09
FA07
F902
F84C
F8CA
F9AB
F9AC
F90D
F92C
FA2B
FA5A
F8E8
F84E
FC4B
0501
0D48
0F3F
0A5F
03F6
0169
02FD
04EF
04A8
0342
02F9
03E0
044B
0394
02EA
034B
0405
03DC
02F9
029E
033C
03E0
03C7
0388
03FF
04B8
0477
0336
02B0
048F
0875
0C3A
0E02
0DD3
0D25
0D37
0DF4
0E5E
0DDB
0CEF
0CAF
0D6D
0E4A
0E4E
0DBC
0DA1
0E25
0E3A
0D5F
0CD2
0DDB
0F26
0D3D
066A
FD70
F735
F5D9
F708
F759
F61A
F50B
F536
F5A6
F531
F451
F451
F55A
F630
F5E2
F4F5
F48F
F4F8
F581
F58F
F53B
F4DD
F48D
F446
F433
F489
F532
F5EB
F6A1
F784
F8A0
F994
F9DC
F967
F8BF
F888
F8EE
F997
F9FA
F9CD
F938
F8C0
F8CF
F92B
F924
F882
F825
F91A
FAEC
FB8A
F9CD
F7F4
FA5A
0296
0C6C
110E
0DC4
0696
01CE
01B5
03A0
0455
03AF
036F
040F
045D
03C2
033D
039F
041A
0397
0298
0285
0382
0427
03A9
030C
038D
0493
045D
02A8
018D
032F
073F
0B64
0DBA
0E3D
0E0D
0E08
0E44
0E5C
0E08
0D8B
0D80
0E1F
0EDB
0EF8
0E78
0E0F
0DFE
0D9B
0C88
0BF0
0D3F
0F6C
0EEC
0962
00C3
F9AC
F6B0
F667
F61C
F532
F4EF
F5C6
F660
F599
F434
F3BD
F466
F501
F4CB
F43D
F418
F468
F4D0
F542
F5D7
F649
F625
F581
F50B
F525
F565
F549
F522
F5C4
F763
F932
FA3D
FA46
F9B9
F91C
F8BD
F8BE
F911
F966
F959
F8F4
F8CA
F94F
FA2A
FA88
FA37
F9EE
FA20
FA0D
F8D3
F78E
F960
002F
096A
0F42
0E03
07DF
029A
01A5
0376
049D
0408
0344
0384
0418
0402
03A5
03F2
0499
0465
0338
026A
02D3
038B
0359
02A0
02AF
0392
03DA
02CD
01DB
0322
06E6
0B2D
0DD6
0E69
0DD7
0D33
0D0F
0D8D
0E60
0EE9
0ED3
0E65
0E03
0DA9
0D36
0CF1
0D27
0D78
0D33
0CA1
0D07
0E98
0EFA
0B34
036B
FB80
F73E
F6A9
F6E6
F621
F527
F53F
F5EC
F5C8
F4B8
F40E
F47A
F518
F4EE
F469
F48F
F557
F5CC
F589
F531
F54E
F593
F5A0
F5CA
F678
F715
F6A9
F57A
F526
F69B
F8B0
F987
F8F4
F882
F930
FA24
FA16
F932
F8C8
F95B
FA18
FA3C
FA15
FA2C
FA33
F9AB
F91F
F97B
FA3E
F9BB
F7FD
F851
FE13
07DF
0F7E
0FC4
09DB
03A9
0180
0297
03AE
0379
0332
03BF
043C
03B6
02E0
030E
0420
04AF
0415
033F
032B
0390
0391
0334
033F
03BB
039C
024D
00FE
01A3
04CD
090E
0C70
0E20
0E9C
0EC3
0EF4
0EFC
0E99
0DE9
0D59
0D29
0D1E
0CE7
0CB2
0D12
0DF7
0E42
0D0D
0B59
0B5B
0D88
0F0E
0C4E
04F6
FCC2
F7C6
F69F
F6CB
F62F
F522
F4E1
F55F
F578
F4CD
F441
F480
F4FA
F4CB
F416
F3D2
F468
F535
F581
F564
F561
F58E
F5A6
F5AA
F5E4
F63A
F621
F591
F57C
F6CC
F901
FA80
FA5B
F94B
F8A0
F8B0
F8D7
F8BC
F8D1
F960
F9EA
F9E2
F9A2
F9D7
FA48
FA12
F942
F916
FA18
FAE1
FA1D
F96C
FC7F
0468
0CDA
0FBC
0B93
0513
01E0
02ED
04E3
0502
03EB
0399
0456
04D2
0469
03EF
0430
04B6
04A2
03FE
0378
033A
02D8
0250
0249
030F
03E7
03DF
031E
0303
04CC
0844
0BD7
0DE7
0E11
0D51
0D06
0DAD
0E88
0E90
0DC3
0D14
0D21
0D73
0D56
0D04
0D3B
0DE8
0E04
0D25
0C7A
0D42
0E81
0D3A
07AB
FF9E
F8E5
F5B0
F510
F4EC
F480
F471
F51E
F5C8
F594
F4AF
F403
F416
F4A3
F529
F56C
F563
F518
F4BD
F4A4
F4E5
F52C
F525
F4F6
F508
F565
F59F
F585
F595
F66A
F7DA
F91A
F9AF
F9E6
FA2C
FA54
F9EB
F910
F871
F871
F8C8
F91E
F993
FA44
FABE
FA83
FA01
FA33
FB15
FB37
F9B2
F844
FA4A
010E
09AA
0F56
0FAB
0C3B
0848
05B2
044F
036C
02F7
0335
03F0
047A
0458
03A4
02DF
0287
02D3
0380
040D
042D
040B
03F3
03E5
03B3
036D
0357
0375
0364
02EE
02A8
03A5
065C
09F8
0CFD
0E74
0E7E
0DE5
0D61
0D31
0D41
0D84
0E0B
0EB3
0EE8
0E3C
0D2A
0CCA
0D76
0E1B
0D8A
0C46
0C2F
0DCA
0EA2
0B73
0415
FC31
F798
F69D
F6BA
F618
F541
F55D
F621
F63E
F557
F475
F474
F4DD
F4C0
F42B
F404
F4B6
F59B
F5D4
F54E
F4B6
F4AA
F518
F573
F572
F56E
F5D3
F655
F634
F55A
F4DA
F5CA
F7C7
F92A
F8FA
F82D
F856
F979
FA27
F9B6
F937
F9B6
FA8B
FA63
F959
F8CD
F95C
FA09
F9ED
F997
F9EC
FA64
F9E2
F957
FBC6
029D
0B0D
103C
0FE4
0BDF
0792
04D9
03A5
033E
0320
02EE
0288
024C
02B5
038E
040A
03D8
0383
037B
0367
02FB
02B7
032E
03ED
0408
037A
032D
038A
03CD
0341
02B4
03CD
06FC
0ABC
0D39
0E01
0DDE
0DA3
0DAE
0E0A
0E69
0E54
0DD4
0D90
0DE4
0E47
0E10
0D84
0D65
0D85
0CEB
0BB3
0BAB
0DB1
0F19
0BC5
036B
FAE8
F71A
F79C
F835
F68F
F47F
F47C
F5F4
F676
F554
F445
F47C
F501
F495
F3D0
F411
F528
F598
F4E0
F435
F4C3
F62D
F72B
F717
F65B
F5A2
F527
F4CC
F497
F4C2
F58B
F6FA
F8AB
F9CD
F9DC
F95B
F95B
FA05
FA5F
F9D7
F92C
F941
F9BE
F9AD
F917
F8F9
F9AA
FA43
FA14
F9C4
FA0B
FA11
F8C2
F7CB
FB17
03FA
0E1C
1300
1071
0A33
0576
03FA
0400
03A1
02D5
0276
02BC
0340
03B1
03E2
0394
02DD
0269
02BF
038A
0421
0458
0458
040A
035B
02C5
02E9
038D
03AF
02F7
029B
0431
07A2
0B17
0CFD
0D72
0D6F
0D71
0D75
0D91
0DCC
0DD8
0D8A
0D51
0D98
0E01
0DE7
0D6F
0D5D
0DC6
0DC8
0D27
0D2D
0E8F
0F05
0B01
0273
FA05
F641
F6AC
F73C
F5D7
F44A
F4BB
F642
F665
F4CE
F3A7
F456
F5B8
F63D
F623
F672
F6D2
F612
F46B
F3A0
F49E
F621
F65E
F537
F42D
F467
F579
F640
F64F
F621
F653
F719
F83C
F93A
F9A0
F98E
F9A6
FA30
FAAF
FA96
F9F4
F935
F8A3
F87F
F91B
FA45
FAE5
FA0C
F86A
F7ED
F93B
FA7A
F9E0
F922
FC63
04DF
0E19
11DF
0EA0
0874
0441
0341
0386
036C
031F
0341
0394
0385
032B
02F9
02F0
02D0
02BC
0313
03C8
046B
04A8
046E
03D2
0334
0335
03FB
049E
03F4
0232
0152
033F
079F
0C08
0E60
0E97
0DE6
0D42
0CF3
0D07
0D5E
0D92
0D6D
0D47
0D84
0DEF
0E01
0DA8
0D47
0CFB
0C9E
0C9A
0DD2
0FBD
0F5B
09D4
0082
F8B7
F668
F80A
F8FF
F735
F4D1
F467
F58A
F603
F537
F49D
F521
F5C1
F55F
F497
F4A5
F555
F55C
F477
F3E4
F489
F5AD
F607
F570
F4F2
F545
F5FD
F640
F5F8
F5CF
F653
F773
F8B6
F9A3
F9F7
F9CA
F972
F939
F93F
F99E
FA48
FAC0
FA7C
F9B6
F967
FA0A
FACC
FA8F
F991
F929
F9AD
F9A5
F826
F767
FB2C
0407
0D61
1188
0F2D
09EF
05F5
044C
0398
02E8
02A2
0322
03CC
03E2
0385
034A
0351
0355
0359
03A2
041F
045F
0421
0393
0316
02F7
035D
0411
0472
03F2
02FA
02F3
04FF
0892
0BBB
0D0D
0CF0
0CDD
0D9F
0EAF
0F13
0E75
0D62
0CB5
0CC2
0D18
0D29
0D12
0D62
0E0C
0E2C
0D54
0CA8
0DA7
0F92
0F07
0976
00B9
F9CD
F790
F7F7
F738
F4B0
F313
F443
F694
F719
F561
F3BE
F406
F577
F630
F5B9
F521
F528
F562
F53B
F4E5
F4EE
F562
F5D0
F5F2
F5F8
F61B
F621
F5AE
F4ED
F4B6
F5B5
F78B
F914
F989
F941
F926
F987
F9C5
F963
F8E7
F936
FA26
FA91
F9EA
F903
F8D6
F92F
F948
F92E
F999
FA57
FA22
F8D3
F8F0
FD7E
05FF
0DC1
1019
0CCD
07B1
047D
03D9
0437
043C
03D3
0383
0396
03F0
044A
045D
0417
03C6
03D1
0421
042D
03B1
030A
02A5
026E
023F
0264
0325
03FC
03FC
0333
0327
0569
09AC
0DD0
0FE2
0FD9
0F21
0EBA
0E5C
0D56
0BD6
0B03
0BBC
0D73
0E8F
0E2A
0D1F
0CE2
0D7C
0D98
0CB3
0C46
0DA7
0F3C
0D47
0648
FD97
F85D
F80B
F92D
F805
F4E5
F2F3
F3A1
F519
F518
F3E4
F384
F4D0
F676
F6D9
F607
F547
F562
F5FC
F674
F6AC
F6D0
F6E3
F6C5
F67E
F658
F689
F6C3
F65E
F536
F444
F4CD
F6D6
F8D0
F945
F884
F837
F94A
FAD1
FB4F
FA8D
F983
F8CB
F82E
F7C2
F832
F975
FA2E
F962
F813
F805
F923
F995
F8EE
F9ED
FF92
08B1
0FF8
110D
0CB2
0746
041E
0354
0372
039F
03DD
043D
0495
04CC
04DB
04AE
043D
03D1
03B9
03CE
03A1
033E
032C
0376
0363
0299
01F3
026E
039E
0426
03B5
03CA
0605
0A0C
0DAD
0F16
0E76
0D5E
0CF5
0D2F
0D6F
0D66
0D3E
0D46
0D75
0D71
0D25
0D17
0DB6
0E59
0DD1
0C47
0B9D
0D08
0E99
0C8C
059C
FD28
F7F2
F714
F76F
F620
F3E7
F352
F4CE
F62C
F5C1
F467
F3F3
F4BF
F598
F5A0
F540
F538
F58D
F5DC
F626
F6A5
F728
F73E
F6E1
F68B
F69D
F6FD
F735
F6D7
F5F2
F553
F600
F80E
FA34
FAF5
FA38
F95D
F986
FA3C
FA45
F970
F8CD
F905
F98C
F9AC
F97A
F936
F8A0
F7BE
F795
F8E7
FA81
FA41
F87A
F8F2
FEFF
08CB
101A
106A
0B40
05CF
0374
03AC
0467
04A3
0476
040B
0381
034A
03C3
0484
04AF
0410
0365
0351
03A1
03D8
03DB
03A6
0302
021D
01E5
02EF
0445
044B
02FB
027D
04DD
0992
0DCD
0F64
0EB9
0DB5
0D7C
0DB5
0D93
0CE9
0C39
0C27
0CD9
0DC7
0E38
0E0C
0DB9
0D81
0D28
0CAD
0CC2
0DB2
0DF8
0B01
0427
FC59
F79D
F6EC
F788
F6AB
F4A3
F383
F3E0
F457
F3F3
F396
F46B
F5F6
F6AA
F601
F50E
F4F1
F589
F614
F64C
F656
F625
F5B6
F581
F603
F6ED
F762
F70A
F664
F616
F652
F6FF
F819
F97B
FA8E
FACA
FA6D
FA3D
FA68
FA5C
F9E3
F9B0
FA45
FAF0
FAA2
F964
F84E
F828
F8AD
F932
F95C
F905
F845
F837
FB12
0206
0AC5
1076
1011
0B43
065F
040E
03CF
040D
0433
0474
04A7
045D
03B7
0353
0354
0337
02CE
02AA
032B
03CD
03F2
03CC
03DD
03FC
03B1
032F
0326
0389
0377
02CC
0313
05ED
0AA4
0E55
0EFF
0DA1
0CB9
0D48
0E2A
0E0F
0D21
0C85
0CD8
0D9F
0E01
0DB8
0D30
0CD0
0C80
0BFC
0B9A
0C38
0DF0
0EE6
0C39
050F
FC7A
F71D
F69A
F81C
F7ED
F599
F39D
F3AB
F4BA
F4E9
F418
F39B
F40D
F4A1
F4C0
F502
F60A
F743
F799
F6F2
F615
F57F
F51B
F500
F5A0
F6EE
F808
F81E
F76A
F6B4
F62F
F57B
F4BA
F4D3
F634
F80B
F93C
F9B2
FA0B
FA72
FA7F
FA0E
F981
F91F
F8CB
F88C
F8CE
F9A1
FA2F
F9AE
F8BE
F8CF
F9F8
FA83
F960
F848
FA45
003D
07CF
0DA5
1024
0FB6
0D54
09CB
062A
03CB
035B
0433
0514
0548
04CF
03E2
02D9
0231
0226
026B
0298
02C7
034E
03FD
0425
038B
02DC
02C1
02EA
02A2
0221
026E
03AE
049E
045C
0406
058C
0917
0CA2
0E47
0E3C
0E02
0E49
0E6E
0DF8
0D8E
0DF5
0EB6
0E9D
0D6C
0C55
0C8B
0DC5
0E85
0DCF
0C6D
0C1C
0D2C
0D53
09AD
0234
FAA7
F738
F853
FA6A
FA0B
F77C
F594
F5B3
F65B
F5D0
F4A2
F48A
F5B7
F6AE
F684
F603
F62B
F6A1
F658
F550
F4AB
F508
F5C2
F611
F61A
F659
F6B2
F6C6
F6BB
F6E6
F6F1
F63B
F509
F492
F598
F76D
F8C3
F929
F927
F92B
F922
F920
F98E
FA42
FA5E
F996
F8E7
F93D
FA02
F9FA
F94B
F963
FA91
FB0C
F979
F7C5
F9CE
00D3
097B
0F2D
107A
0F41
0D67
0B03
07CC
04B7
032C
033F
0395
032B
026B
024D
02EC
0383
0376
02E2
0255
024A
02D4
037C
0392
02F0
0239
021C
0289
02F1
031B
0339
0339
02A7
01AA
01BA
0454
08EF
0CFA
0E69
0DBA
0CF0
0D17
0D8C
0D87
0D4B
0D7A
0DEC
0DEA
0D71
0D6B
0E50
0F19
0E57
0C41
0AF9
0C2B
0E92
0E80
095B
00BA
F979
F749
F934
FB16
FA3D
F7DD
F6AB
F746
F7DE
F719
F5D7
F5A0
F655
F685
F5C0
F534
F5BC
F674
F614
F4E6
F45A
F501
F5E7
F5FD
F563
F4EC
F500
F560
F5BF
F5F2
F5B5
F4F9
F479
F53E
F739
F916
F9C9
F9B5
F9B1
F9A8
F90D
F83D
F859
F988
FA75
FA10
F92A
F953
FA8E
FB54
FAE9
FA49
FA45
FA14
F923
F939
FD0B
0480
0BE9
0FB2
0FD6
0ECB
0DBF
0B96
07AE
03DD
0277
0356
043A
03C3
02CF
02B9
0371
03E6
03AB
0358
0378
03C5
03C4
038E
0398
03F1
0428
03DD
0322
0262
0221
0283
02FB
02BC
01DD
01CE
03FE
0802
0B99
0CDC
0C1F
0B44
0B70
0C1A
0C63
0C85
0D37
0E36
0E5F
0D5A
0C5A
0CA3
0DD9
0E6C
0DC6
0D38
0E22
0F72
0DFC
07DF
FF36
F89E
F6E2
F88C
F9F1
F926
F75B
F69A
F720
F79E
F759
F700
F73C
F782
F6EC
F59F
F498
F453
F467
F46D
F494
F506
F540
F4BB
F3F1
F3F2
F4F5
F5FC
F624
F5A6
F51D
F497
F404
F402
F556
F79B
F951
F992
F917
F91A
F9BF
FA38
FA45
FA76
FAEB
FADE
F9F8
F91C
F928
F9A0
F997
F968
FA29
FB7D
FB75
F98B
F8AF
FC8C
04D0
0CD9
109D
1082
0F6B
0E54
0BC7
0752
0347
022B
037F
0488
03D1
029D
02AB
03DA
04C5
04D4
0498
0489
046E
0414
03B7
0386
0345
02CA
0275
02C4
0396
043E
0449
03C5
02F0
022A
025B
0488
0867
0BEF
0D26
0C47
0B5E
0BD0
0CE7
0D3A
0CB0
0C69
0CE4
0D50
0CFA
0C7D
0CCA
0D88
0D8A
0CCD
0CDF
0E82
0FA5
0CED
0592
FCFB
F7D2
F7A1
F9D8
FAF9
F9F8
F832
F6F4
F619
F517
F44C
F481
F593
F659
F621
F587
F588
F617
F64E
F5D1
F544
F54A
F5AA
F5D4
F5C2
F5C0
F5AD
F524
F454
F41B
F4DD
F5D2
F5F7
F581
F59F
F6DB
F86A
F954
F9A0
F9E7
FA51
FA8D
FA80
FA4F
F9E1
F915
F86A
F8C0
FA15
FB22
FAF8
FA72
FAD6
FB7E
FA77
F81F
F83D
FDE9
070E
0DEE
0F55
0DA5
0CEF
0D8A
0C5D
0804
033F
0188
02D4
0451
044A
0396
0372
03A9
0372
02F0
02D1
0308
02F2
028E
02A6
0372
040F
03C5
0307
02A9
02B9
02EE
0371
0453
04A7
0384
01FD
02D5
0743
0CCE
0F91
0E8E
0C79
0C12
0D18
0DA3
0D3D
0D0F
0D93
0DCE
0D26
0C90
0D06
0DC2
0D4F
0C15
0C39
0E4F
0F6D
0BF6
040B
FBF5
F7E6
F822
F9A7
F9D2
F88C
F72F
F66C
F5E1
F54B
F52A
F5E5
F6DE
F6F8
F5F9
F4F3
F50D
F633
F733
F72A
F675
F604
F616
F614
F58D
F4DE
F49F
F4F0
F591
F652
F701
F729
F676
F568
F52E
F67F
F8B8
FA6A
FAC2
FA26
F97F
F957
F9B3
FA45
FA9C
FA78
FA20
FA11
FA2B
F9DC
F940
F95E
FA8C
FB41
F9DF
F7C8
F927
003B
09A7
0F52
0F18
0CC8
0CBC
0E57
0D9D
0927
041F
0210
02C1
036B
02CB
0217
0246
0286
0200
0185
0227
0348
037F
02CB
027C
031A
03AE
0369
02DF
02F2
0373
03AA
03BE
0440
04A0
03B5
0233
02E1
0712
0C3C
0EA2
0DC4
0C83
0CF5
0DF4
0D86
0C1F
0BD8
0D18
0E01
0D70
0CAF
0D21
0DD6
0D30
0BEC
0C67
0EB3
0F46
0ABB
0209
F9E8
F62E
F6B1
F89B
F99F
F93C
F7F3
F671
F56B
F544
F5A1
F5CE
F59F
F588
F5D4
F63C
F651
F60B
F5BD
F59D
F5A3
F5C8
F61C
F68B
F6C2
F68C
F606
F563
F4D2
F4B0
F55A
F682
F720
F68D
F58A
F593
F729
F92D
FA24
F9D3
F954
F9AA
FAA6
FB5A
FB51
FAF7
FAD9
FAE7
FA9A
F9CF
F94B
F9EE
FB2E
FB0E
F8AA
F693
F91F
016C
0B0F
1019
0F57
0D2D
0DC9
0FEC
0EF8
0970
033E
00FB
02C4
050D
054C
040E
02F4
027F
0261
0294
0320
0366
02CD
01F8
022B
036B
0448
03EC
0343
0367
03F1
03E2
0356
0325
0335
02B4
0215
035E
0784
0C71
0EF5
0E7D
0D60
0D74
0DF0
0D74
0C77
0C50
0CD5
0CCD
0C3A
0C7B
0DCE
0E6F
0D44
0C1C
0D66
0FEC
0F10
083A
FE81
F79B
F60C
F7B7
F963
F9D4
F954
F81A
F651
F4DC
F4B1
F574
F5B0
F4CF
F3F1
F451
F5A0
F6A9
F6F9
F6FE
F6E6
F658
F54E
F46A
F425
F43E
F445
F45A
F4E1
F5B6
F635
F61C
F5CE
F58D
F528
F4C0
F535
F716
F96B
FA83
F9DC
F8C1
F8A7
F98C
FA35
F9DB
F906
F8B8
F930
F9DC
FA3D
FA62
FA6B
FA1C
F939
F862
F94F
FD9A
04D1
0BF6
0FBC
0FA2
0E3E
0E23
0EF0
0E22
0A80
05D9
0304
02D8
03DA
047B
04A3
04D9
04FF
049B
03C4
0304
0296
0257
024B
02A1
032D
037D
0387
03D8
04B3
0576
055B
048B
03D0
0351
02A3
023C
039D
0753
0BA3
0E35
0E93
0E21
0DE8
0D88
0C9D
0BFC
0C96
0DCD
0E31
0DA2
0D4B
0D66
0CB9
0B21
0ADF
0D87
1083
0EE8
0740
FDDD
F857
F7CD
F8E8
F8D2
F80D
F80A
F833
F6FE
F4C7
F396
F44C
F58D
F5D3
F545
F4EC
F500
F4E6
F48B
F498
F533
F594
F53A
F4C0
F4D9
F538
F543
F536
F5A7
F649
F62F
F553
F4DB
F56F
F61B
F5AB
F4A4
F4D4
F6C4
F8D2
F954
F8C2
F8CD
F9ED
FAE9
FAB3
F9BF
F93A
F998
FA58
FACD
FAAC
F9FF
F920
F8AF
F908
F9A5
F9BC
F9D2
FBE5
0134
0829
0D76
0F49
0EDB
0E84
0EE2
0E82
0C0E
0831
04F9
03C3
0429
04C4
0491
038C
026D
01F4
0266
0377
0499
0555
0566
04DC
0421
03B5
03B0
03B3
0364
02DC
027E
027D
02C7
033D
03C2
03FB
0394
0314
0400
073E
0B71
0DE4
0D91
0C54
0C91
0E46
0F7E
0F2D
0E65
0E5C
0E90
0DEF
0D06
0D5E
0EC7
0F1B
0D6F
0BEA
0CD8
0EBC
0D54
06BF
FE27
F85D
F6ED
F79E
F815
F829
F86B
F851
F717
F573
F4E4
F589
F601
F577
F4BB
F4D7
F576
F571
F497
F3F6
F45A
F550
F5EC
F5E5
F57F
F501
F4C6
F544
F64B
F6C0
F5D8
F475
F44B
F5A7
F6CB
F627
F48D
F458
F67A
F95A
FAE2
FABD
FA03
F98A
F95C
F95F
F994
F9AC
F942
F893
F866
F8F9
F98F
F996
F99E
FA60
FB22
FA7B
F915
FA3C
0055
0948
0FE6
1120
0EE6
0D6A
0E50
0F6D
0DE6
0989
04B3
01B3
0108
01C9
02EC
03E1
0480
04C7
04B6
045F
03F9
03C3
03B9
0394
0331
02C4
028D
0278
0247
0206
021A
02BC
0399
0430
0457
0420
0380
02C2
0323
05F2
0A99
0E6F
0F41
0DCA
0CC9
0DB2
0F45
0F91
0E7B
0D6C
0D16
0CE3
0C84
0CA3
0D76
0DE6
0D39
0CA1
0D9D
0F01
0D55
06DD
FE40
F813
F631
F6B2
F735
F786
F86A
F95C
F8FA
F741
F5C1
F57C
F5AC
F523
F414
F3B4
F476
F576
F5BE
F56A
F538
F582
F60E
F688
F6A8
F63B
F57D
F528
F59E
F643
F62D
F565
F4EB
F555
F602
F60D
F5AD
F5FA
F752
F8C1
F93B
F8DF
F88B
F8B0
F91D
F997
FA07
FA44
FA35
FA2E
FA92
FB20
FB14
FA46
F9A1
F9D9
FA27
F962
F87E
FA9A
0179
0A8D
10C2
1169
0E95
0C79
0D00
0E77
0E14
0AFF
06CF
03AD
0290
02F8
03D5
0467
0489
0459
03D5
0312
0293
02ED
03EA
0486
0426
0357
0302
0325
0305
026E
0223
02B1
0374
0384
0320
0339
03BB
0392
02D8
039F
0765
0C7A
0F5A
0EA1
0C7F
0BD8
0CF8
0DF0
0D7E
0C43
0B4D
0AE2
0B1E
0C62
0E42
0F1F
0E30
0D18
0DDF
0F6B
0DC9
06DF
FDBB
F7BF
F6E9
F86A
F8DA
F811
F7DC
F881
F87D
F729
F5D9
F5CE
F672
F660
F57A
F4EB
F551
F5E4
F5BD
F512
F4A7
F4AF
F4DB
F521
F59B
F5F3
F5A9
F4F1
F4A9
F540
F61C
F670
F640
F62A
F65F
F65A
F5D9
F57B
F60C
F76D
F8B7
F942
F93F
F953
F9E4
FAC7
FB6E
FB71
FB14
FAFE
FB58
FB6D
FA80
F900
F84B
F8FD
F9F6
F9D9
F96A
FB5F
013A
08EA
0E6B
0FB4
0E6B
0DBC
0EEC
105A
0F88
0BCB
06F2
038B
02B4
036F
03EE
0378
02DC
0318
03E7
0429
0386
02E4
0308
0382
037C
030B
02F8
036F
03BD
0380
0350
03B8
0429
03C8
02FB
0309
0405
0472
0393
0311
0519
094D
0CDF
0DCE
0CF3
0C5E
0CA8
0CD9
0C78
0C53
0CFF
0DE0
0E33
0E2B
0E3F
0E21
0D85
0D41
0E37
0F20
0CDE
0615
FD96
F7FE
F6FA
F81E
F87A
F7EC
F817
F93F
F9DD
F8F6
F76B
F685
F63A
F5B1
F4CF
F45F
F4B2
F50F
F4DA
F482
F4C2
F566
F595
F51D
F4B8
F4F7
F57D
F597
F52C
F4C5
F4C5
F503
F531
F554
F59D
F5FF
F632
F626
F635
F6CA
F7EF
F93F
FA40
FACA
FB0C
FB2E
FB04
FA74
F9F7
FA3C
FB27
FBA1
FAD6
F96D
F8D5
F950
F97A
F869
F7C7
FAAE
01EE
0A5F
0F9C
1032
0E94
0E05
0F4F
1085
0F72
0BC1
0717
039C
0269
02F3
03AC
037A
02AE
0269
02FF
0384
0314
022B
020E
0329
0492
0532
04EA
044F
03C7
0358
032F
0393
0442
046B
03A9
027F
019E
0117
00E4
01C2
049F
0907
0CDF
0E48
0D8B
0C93
0CAA
0D54
0D76
0CEA
0C75
0CA5
0D4B
0DD9
0DE0
0D50
0CB9
0D1A
0EAC
0FB6
0D5F
0693
FDEE
F7E3
F6AC
F88E
FA4A
FA8C
FA35
FA1B
F9B3
F848
F660
F531
F50A
F521
F4F3
F4EE
F57D
F60C
F5B6
F49A
F3CB
F3E1
F45C
F498
F4D6
F5AB
F6BF
F6DB
F572
F3A3
F328
F468
F61D
F6E4
F6AA
F658
F682
F6F1
F75B
F7FC
F91A
FA4A
FAC0
FA59
F9F0
FA46
FB02
FB46
FAF4
FAD2
FB30
FB3E
FA3E
F8F3
F8E2
FA06
FA58
F889
F6B5
F8F6
00BF
0A79
109E
10E8
0DE8
0BC3
0C3B
0E00
0ED1
0D76
0A23
060F
02F2
0204
02E1
03DA
03CE
0361
03D3
0519
05D2
0525
03D3
0313
02FE
02DB
028F
02C6
039D
0411
035C
0230
01D7
0281
032D
0316
027A
01DF
016E
018E
034E
0744
0C14
0F1F
0F28
0D93
0C92
0CBA
0D12
0CF5
0CD6
0D34
0DAC
0D92
0CFA
0CA3
0D13
0E37
0F80
0FBC
0D22
06C6
FE85
F869
F70D
F8FD
FA8A
F9F6
F8BF
F8D0
F9AF
F973
F7A8
F5E9
F576
F5A2
F535
F45D
F425
F49C
F4C7
F460
F466
F586
F6C1
F69C
F52F
F41A
F459
F514
F50C
F475
F489
F59F
F6B1
F6E1
F69A
F6C1
F753
F786
F720
F701
F7FF
F9AB
FAB8
FA89
F9CC
F967
F95D
F929
F8D5
F91A
FA3D
FB61
FB70
FA94
FA19
FA9E
FB1C
FA72
F9A3
FB68
010C
086C
0DB6
0F10
0DE1
0CC7
0CF6
0DD5
0E43
0D70
0AE8
06EE
0312
0162
025D
0448
0525
04CF
047A
0494
0442
030A
01F4
0232
034F
03BD
030B
0273
02E4
03A4
038E
02D5
0293
030D
0369
0311
0264
01DF
017D
0179
02E5
0676
0AE4
0DB8
0DFE
0D3A
0D27
0D91
0D4C
0C68
0C30
0D2A
0E46
0E63
0DBF
0D5E
0DAA
0E59
0F10
0F23
0CEB
070B
FEF5
F8B5
F71D
F8BF
F9F5
F939
F82E
F86B
F90B
F83E
F639
F4F3
F54E
F5F6
F5A0
F4E8
F50F
F5D8
F5FE
F54E
F4EE
F57B
F606
F583
F45E
F3E6
F484
F551
F582
F556
F563
F59C
F5AC
F5AD
F5DE
F600
F5B9
F575
F622
F7F4
F9E8
FACF
FA8A
F9ED
F9B3
F9D9
FA02
FA10
FA19
FA25
FA33
FA59
FA97
FAC1
FAB0
FA65
F9E7
F95F
F9A4
FC09
0115
0773
0CB0
0F3F
0F84
0EE8
0E50
0DD3
0D6A
0D0C
0C26
09DE
066F
0378
0265
02DA
0366
0357
032A
0343
0328
0260
0177
016B
0240
02F0
02D7
027A
0290
02EC
02EF
028B
0243
0265
02DC
0391
0459
04AD
0417
032C
0381
0611
09E4
0CE1
0DFF
0E01
0DFE
0E0D
0DC2
0D50
0D4D
0DCA
0E40
0E4E
0DFB
0D6C
0CEC
0D1A
0E39
0EEE
0C8E
05EA
FD90
F802
F735
F8D1
F968
F84D
F74C
F765
F784
F67E
F4E8
F428
F46E
F4BC
F497
F49D
F52C
F592
F52E
F497
F4C9
F5BD
F696
F6E3
F6EA
F6C9
F644
F57B
F522
F580
F5D7
F572
F4E8
F56D
F6D5
F778
F68A
F58A
F66A
F8FC
FB36
FBC1
FB2D
FA90
FA13
F96B
F8F7
F978
FABF
FBA7
FB98
FB36
FB1B
FAC6
F99F
F892
F9A6
FDE7
0443
0A73
0E9B
1017
0F7D
0E33
0D8D
0DAF
0D4A
0B04
0747
040A
02AC
02AF
02D8
02DF
033E
03DC
03FB
036A
02EE
0323
037B
02F9
01B2
00E2
016F
02CB
03B0
0388
02BF
0213
0201
0295
0362
03CB
03CD
0459
067F
0A1C
0DB4
0FAF
0FB3
0EA3
0D8D
0CE5
0CA5
0CBB
0D0F
0D62
0D76
0D3B
0CDE
0CD1
0D94
0ECE
0EA3
0AE5
03B3
FC4B
F867
F8A4
FA3B
FA68
F939
F882
F8CC
F8A9
F71B
F518
F41B
F428
F44E
F44F
F4BA
F588
F5E0
F563
F4DE
F520
F5C1
F5D9
F57D
F590
F62A
F64A
F57F
F4C5
F508
F5B6
F5C6
F56D
F5A6
F658
F643
F521
F4A5
F65F
F95A
FB01
FA59
F90C
F8EF
F9D4
FA82
FAC2
FB18
FB3F
FA76
F930
F90F
FA7F
FB8E
FA53
F81B
F8C5
FE7F
0704
0DC2
101D
0F04
0D1E
0C60
0D1B
0E2A
0DD3
0B2E
0734
041D
0359
043C
04F6
0496
03B0
031E
02E2
0296
025F
02A5
033F
037E
0317
0286
0275
0303
03BC
040C
03B5
02F8
0262
0259
02AF
02D3
02B4
0343
059C
0975
0CE3
0E1A
0D46
0C37
0C6D
0DB7
0EC5
0EA6
0DA2
0CB2
0C5D
0C4F
0C20
0C2E
0D2F
0EB7
0EA9
0AE8
03DD
FCCA
F8F2
F89B
F970
F99F
F97E
F9E1
FA2D
F917
F6C4
F4DF
F47D
F4DE
F4CB
F454
F46B
F535
F5D4
F5E5
F60C
F69E
F6C7
F5DE
F4C0
F4CF
F5FD
F6DD
F69C
F5F2
F5DD
F63F
F66B
F66F
F6C8
F719
F66A
F4FE
F4A5
F67A
F93D
FADD
FAFB
FACC
FAE7
FA9C
F994
F8D0
F921
F9A5
F908
F7F0
F873
FAC9
FC32
FA8B
F7EA
F8EC
FF61
080D
0E03
0F59
0E08
0CFD
0D68
0EA1
0F66
0EAC
0C06
0821
04AC
02FC
02D6
02FE
02BE
026D
028D
0302
0356
035F
0359
037B
03B4
03DB
03DC
03B6
037B
0365
039A
03D2
038D
02CD
022E
0204
01DC
0164
017B
037F
0773
0B62
0D34
0CDF
0C4F
0D0C
0E88
0F1E
0E49
0D39
0D41
0E35
0ECA
0E47
0D74
0D72
0DDA
0C78
0796
0054
FA21
F78A
F7F8
F8EE
F8F7
F8BE
F94B
FA1C
F9C6
F7EE
F5C8
F487
F42E
F43B
F496
F544
F5CA
F5AB
F546
F564
F5FB
F628
F594
F529
F5D2
F705
F763
F6AF
F60A
F626
F65C
F603
F5A7
F5FB
F668
F5E8
F4FC
F571
F7E0
FA79
FB30
FA48
F993
F9A8
F96D
F884
F857
F9B9
FB01
FA2E
F80C
F761
F8EF
FA3E
F957
F84F
FB39
02DC
0B35
0FC7
1000
0E8D
0DAB
0DA0
0DFC
0E74
0E55
0C81
08ED
055C
03C5
0431
04EB
04AC
03CE
0336
0308
02FF
0341
03EF
0466
03DE
02A5
01EF
0262
0366
040C
041E
03E9
037C
02C5
0235
026F
0339
0390
0342
03AB
0607
098E
0C28
0CEC
0CFF
0DBB
0EDC
0F17
0E27
0D4B
0D8B
0E45
0E1E
0D09
0C7A
0D5B
0E59
0CBD
0725
FF42
F8BE
F62C
F6FB
F886
F8F4
F8A1
F8CD
F994
F9BD
F864
F627
F487
F459
F52B
F5FD
F623
F59D
F4ED
F4C9
F56F
F62E
F61B
F557
F507
F5B2
F66D
F627
F552
F559
F696
F7B8
F79A
F6CD
F67B
F66F
F59E
F470
F4D4
F764
F9F8
FA43
F8D7
F829
F908
F9C1
F8FB
F7BD
F7B2
F88A
F8C6
F882
F952
FB1C
FB61
F927
F7C0
FB74
03F8
0C3B
0FF1
0FA0
0E8B
0E5E
0E6F
0E50
0EB2
0F52
0E31
0A47
05AA
0361
03CE
04B5
0484
03E9
0407
048A
0470
03C2
035F
035C
02F2
022B
0245
03BC
0514
04A3
02CE
0170
016E
0213
0288
02C8
02DF
0276
01DD
02B7
0652
0B66
0EC0
0EC2
0D33
0CD9
0E15
0F0C
0E99
0DAB
0D8E
0E04
0DEC
0D2D
0CE9
0D9A
0DB0
0ADE
04BB
FDA9
F8E9
F7D8
F90F
FA01
F966
F818
F7A6
F845
F8A8
F7C0
F608
F4C5
F47B
F49F
F48F
F450
F453
F4D6
F5B2
F680
F6CE
F65D
F582
F51C
F5B8
F6C0
F71C
F6A0
F627
F627
F615
F59B
F580
F674
F794
F743
F589
F471
F581
F7A1
F892
F7F4
F780
F84C
F966
F9B1
F998
F9EA
FA20
F959
F846
F876
F9BC
FA11
F8FA
F970
FE9C
0726
0DEF
0FDB
0EE9
0EA6
0F83
0F8C
0E60
0DDC
0EB3
0EC0
0BF1
0784
04A6
0463
04B4
03CB
027D
0275
0383
0436
0438
0474
0519
0506
03A5
0214
01D4
02DD
03D7
03E3
0353
02B6
0229
01D2
021B
02CE
02F8
028B
0340
069F
0B72
0E8D
0E6A
0CE4
0CB1
0E03
0EBC
0DAF
0C3F
0C30
0D2B
0D8C
0D11
0D2E
0E67
0EA4
0B23
03DD
FC2B
F7CA
F776
F8C9
F925
F83E
F79C
F830
F91F
F8F5
F76F
F5AE
F4B8
F464
F40A
F3BB
F424
F541
F602
F59E
F4AE
F478
F55A
F67B
F6E8
F67F
F5B7
F4F7
F476
F46E
F4F2
F5A4
F5FF
F602
F60C
F619
F5AC
F4C7
F468
F57A
F79E
F989
FA5E
FA43
F9C4
F930
F8BE
F8B8
F91B
F969
F967
F9A9
FAA0
FB5B
FA8C
F922
FA67
005E
08A3
0E63
0F6C
0E05
0D84
0E6D
0EFE
0E8D
0E59
0EDD
0E55
0B2F
06C3
0406
03F0
04B9
04A1
0420
0484
0588
0596
042C
02A8
0256
02BE
02A0
01EC
01C6
02D3
0468
055E
0522
03F9
02B1
0233
02CE
03BB
03CD
031F
0385
0690
0B26
0E36
0E31
0CC8
0C8F
0DBB
0E5C
0D82
0C85
0CCE
0D9B
0D3C
0BEA
0BBB
0D4B
0DD8
0A1E
0299
FBA2
F8F3
F9FB
FB29
FA33
F828
F767
F86D
F966
F89B
F671
F4B2
F45A
F4B2
F489
F3CB
F375
F41A
F508
F52F
F49C
F473
F565
F6B5
F715
F636
F4FE
F465
F47A
F4AB
F4A4
F496
F4C1
F522
F598
F607
F63C
F607
F5A1
F5C1
F6EB
F8C3
FA4F
FADD
FA86
F9E6
F98D
F9AE
FA24
FAA2
FADF
FAB8
FA31
F964
F8B0
F91C
FC11
01F8
090A
0E29
0F88
0E29
0C9B
0C79
0D93
0EF6
0FEA
0FD1
0DFE
0A7C
06B5
046B
03EA
03F3
039A
0364
040C
04FA
04EE
03D2
02EE
032B
03F3
0423
0394
02FE
02C0
028A
0242
0262
0314
03BE
03E2
03D8
03FF
03FD
0392
03C7
060E
0A19
0D88
0E74
0D9A
0D1A
0D86
0D83
0C66
0B90
0C5B
0DDE
0E40
0D93
0DAB
0ED4
0E54
0964
0117
F9F2
F75E
F872
F9A8
F8EE
F742
F6B0
F7C7
F935
F94A
F79E
F55F
F416
F41D
F477
F441
F3D7
F43E
F583
F666
F5E1
F49B
F425
F4F6
F5CE
F572
F43D
F380
F3E0
F4D7
F59A
F5DB
F5C1
F59F
F5B2
F5EB
F5EF
F5A2
F5A2
F6D1
F914
FAFA
FB31
FA27
F97C
F9E7
FA90
FAA8
FA94
FABF
FA5E
F8B4
F740
F924
FFA8
0832
0E83
10B6
1045
0F68
0ECA
0E27
0DDD
0E88
0F8A
0F34
0C90
087D
04E4
031F
0321
03C0
03C7
0305
026F
0307
048A
0574
04B4
02FF
01F1
01FD
0243
0252
02E2
0439
051A
0459
02C9
024D
0333
03D9
0351
0329
057D
09E1
0D9B
0EE9
0EA5
0E4D
0DF6
0D1F
0C4D
0C65
0D0F
0D36
0D04
0DB5
0F01
0E11
0875
FFAE
F864
F5CF
F6E2
F879
F8FC
F907
F963
F9E0
F9F6
F96F
F851
F6CC
F569
F4B5
F499
F477
F41B
F429
F512
F606
F5D5
F4C3
F479
F5AB
F6D8
F63D
F443
F2EE
F359
F4A6
F56D
F559
F511
F51C
F55E
F576
F544
F514
F57B
F6EE
F8FB
FA2D
F981
F7FB
F7B0
F912
FA52
FA0B
F93B
F96F
FA0F
F958
F801
F9C1
00E5
0A7C
10CD
1178
0F69
0E67
0EAF
0E56
0D34
0D23
0E93
0F1C
0C6A
0766
036A
02A5
042F
05A8
05C5
04EB
03FA
035E
0315
02F1
02DB
02F6
0362
03C8
03A7
0338
0364
0461
050C
044E
02BA
01EF
027E
034C
0378
03F3
0640
09F0
0CB7
0D43
0CC2
0CFB
0E0E
0EE7
0F02
0EAC
0E0D
0D3B
0CFE
0E12
0F2E
0D21
063C
FD2F
F70B
F62D
F830
F961
F8D7
F838
F8A1
F96C
F99F
F923
F84B
F72E
F5FB
F548
F579
F607
F602
F540
F475
F41D
F404
F41B
F4D0
F617
F6E1
F656
F511
F45D
F48B
F4DD
F4DC
F4F6
F597
F64F
F652
F58D
F4C3
F4BD
F5BF
F7A6
F9CE
FAF4
FA3A
F889
F7E4
F8E4
F9E6
F96E
F857
F858
F943
F976
F92B
FB60
020F
0A8F
0FBD
0FC1
0DC8
0D72
0E90
0ECA
0DDD
0DC3
0EEC
0ECD
0B2E
0591
01DB
01FC
0427
056F
04F4
03F0
0390
03E7
0480
04F5
04E1
040B
02CB
01DF
01BA
0239
02EB
0373
03B4
03D3
0404
043A
0416
0377
0310
041E
0716
0AC2
0D3E
0DE1
0D93
0D53
0D3D
0D29
0D51
0DBA
0DC1
0D32
0D20
0E70
0F97
0D43
062D
FD80
F81E
F797
F907
F912
F7AE
F713
F839
F9D9
FA70
F9D8
F8AD
F742
F5CB
F4D9
F4E9
F595
F5D6
F540
F478
F444
F48C
F4BC
F4AC
F4AB
F4FB
F59E
F659
F6AB
F615
F4DF
F420
F493
F59B
F5E6
F503
F3D4
F379
F43B
F5C8
F7E3
FA1E
FB58
FAAE
F8FB
F841
F933
FA5E
FA67
F9E4
F9EE
F9EB
F89E
F741
F97A
00F0
0A26
0F9A
0FC3
0E36
0E83
100C
1026
0E9E
0DC7
0E86
0E9C
0BC6
0710
03BC
0360
0470
049E
0397
02B3
02E4
03D2
04BA
0524
04D5
03D6
02C1
026F
0325
0437
04B1
043F
0371
0319
0366
03B4
0352
0287
0288
0455
0795
0AC7
0CAD
0D58
0D8D
0D9B
0D58
0D0E
0D60
0E14
0E11
0D25
0CCA
0E0F
0F26
0C95
0562
FCF0
F7D6
F738
F85C
F88C
F7F0
F812
F90C
F983
F8D0
F7BA
F705
F673
F589
F493
F437
F475
F4B4
F4C1
F518
F5F7
F6B6
F689
F593
F4CC
F4E0
F595
F625
F5E8
F4E2
F3E5
F3EC
F510
F651
F69B
F5E3
F507
F4DB
F595
F6FC
F8A6
F9DD
F9E4
F8F2
F872
F968
FAC8
FAA8
F91B
F86B
F9B1
FAC0
F93B
F6F0
F8EB
0143
0B92
112C
1050
0D59
0CDE
0EBD
0FE3
0F28
0E1D
0DBF
0CB7
09A3
059C
0332
035D
04A3
0538
04F3
04B4
04B0
0454
038A
0316
0386
045A
04A5
042A
038A
0373
03CA
03E3
0372
02FE
031B
036C
0314
0223
020F
0439
082C
0BD7
0DA5
0DE1
0DDB
0E25
0E62
0E5E
0E51
0E0E
0D11
0BE4
0C29
0E32
0F2F
0B7A
0309
FA6E
F675
F763
F96A
F971
F80F
F792
F898
F9B9
F9BE
F8CD
F785
F62C
F500
F491
F517
F5E0
F5F1
F525
F43D
F3CB
F396
F353
F35E
F435
F592
F692
F6BE
F668
F612
F5D6
F584
F520
F506
F57F
F64A
F6B8
F67E
F647
F715
F8EC
FA68
FA21
F86E
F73A
F7BF
F910
F993
F96B
FA22
FBD0
FC4D
FA5D
F89D
FB61
035C
0C05
102B
0F54
0D5D
0D5F
0E9C
0EE2
0E12
0DB2
0DE1
0CB3
0911
04D6
02ED
03E5
0566
051E
035A
023C
02E7
045D
051F
04F5
04BB
04D3
04AB
03D1
02D9
02B0
0342
037D
02E6
027C
035D
04DF
0523
03C2
02E0
04C7
090E
0CE8
0E42
0DA6
0CE9
0CEF
0D69
0E06
0EAD
0EB4
0D5C
0B89
0B7B
0DAB
0ED1
0AD9
01E7
F90E
F55C
F6EB
F9A8
FA45
F91D
F850
F8A0
F918
F8EF
F854
F79E
F6B4
F599
F4C0
F47E
F494
F494
F485
F4B9
F52A
F565
F52F
F4D8
F4B8
F4AB
F474
F451
F4B7
F595
F64A
F65D
F5FA
F59E
F579
F54E
F4F0
F4C9
F5A2
F79F
F9B1
FA67
F98E
F88B
F8D2
FA15
FAA6
F9CD
F8FC
F9D4
FB85
FB99
F9B6
F935
FDA3
0632
0DFD
1105
0FD6
0DD5
0D11
0CF6
0CA3
0CB1
0DC7
0E9D
0CFA
08A5
0437
0277
0389
052E
056B
0465
038F
039D
03E0
0383
02C5
0286
02F5
0355
031C
02C7
0324
0409
046B
03E3
0372
0406
04DB
0465
02E7
02D3
05D6
0A72
0D87
0DE0
0D23
0D37
0DF8
0E22
0D82
0CF7
0CBB
0C35
0BB6
0C9E
0EB3
0EBB
0992
007D
F8B9
F63F
F7F8
F9D3
F9A2
F8A3
F8A6
F967
F97A
F88C
F784
F6E2
F635
F540
F499
F4D2
F596
F60B
F5CE
F532
F4AA
F45B
F445
F47D
F4FA
F578
F5C0
F5E5
F600
F5EC
F587
F516
F507
F562
F5BE
F5AA
F524
F4B5
F51F
F6A5
F890
F9A8
F972
F8D0
F906
FA21
FAE3
FA88
F9FF
FA81
FB73
FB13
F99A
FA28
FF4E
0755
0D73
0ED8
0D50
0C6A
0D39
0E16
0DE9
0DC2
0E97
0F05
0CD3
0839
0424
02F3
03FC
04C9
0412
02C9
026A
0316
03BD
03A2
031E
02F1
0352
03DE
0430
043C
0422
03DD
0353
02C4
02D9
03C6
04A7
0451
030F
02D3
0535
0970
0D00
0E39
0DB8
0D2A
0D3C
0D5E
0D11
0C9C
0C53
0C2F
0C59
0D3D
0E49
0D4D
0867
00A4
F9C5
F6DA
F77D
F8E4
F92C
F8D1
F902
F9AE
F9DA
F921
F809
F701
F5F8
F4F0
F464
F4AC
F571
F600
F61B
F610
F60D
F5C2
F4E8
F3E6
F390
F43D
F561
F616
F5F5
F559
F4EC
F504
F55C
F584
F56D
F55D
F582
F5E4
F6B3
F833
FA14
FB44
FAF1
F9A6
F8E8
F981
FA9F
FB1C
FB06
FB0F
FAE6
F98D
F7C4
F8BC
FED1
0800
0F19
10E7
0F28
0DBF
0E05
0E45
0D47
0C5B
0CED
0DB5
0C04
078A
0336
01E0
033C
04BC
04C2
03E9
036F
038D
03C6
03EF
0433
0468
043B
03D6
03B2
03C6
038E
02EE
029A
032F
042E
0469
037D
027C
02F3
057D
094C
0CCE
0EA2
0E7C
0D6C
0D00
0DA1
0E16
0D15
0B3E
0AAF
0C44
0DC5
0BC5
0566
FD9F
F878
F75C
F882
F96A
F930
F898
F88E
F91B
F985
F912
F7AC
F5FD
F4EF
F4DB
F53A
F550
F523
F54F
F5F1
F640
F59C
F4A9
F4A8
F5C9
F6C9
F688
F577
F4F1
F561
F5E2
F5B2
F53A
F538
F57F
F566
F52A
F5E8
F7F3
F9FC
FA8F
F9EF
F997
FA09
FA28
F92C
F82E
F8B5
FA33
FA7A
F915
F8F6
FD63
05A3
0D12
0FE5
0EDF
0D8D
0DCD
0E78
0E2D
0DA7
0E3F
0F2D
0DFC
09DC
0524
02B5
02CC
0353
02EA
024C
0297
036C
03A2
0330
032F
0407
04B2
0447
035F
0336
03E2
045C
041F
03D5
041E
046D
03D0
028E
0241
042B
07E9
0BDD
0E7C
0F15
0E12
0CD5
0CC0
0DCF
0E8B
0DF2
0D05
0D73
0EA2
0D5E
0762
FEC0
F85D
F6EB
F876
F95E
F885
F78B
F7CD
F8A0
F8AF
F7C4
F6A0
F5C1
F52C
F50E
F5A7
F679
F684
F5A0
F4DA
F502
F58E
F596
F54B
F582
F621
F617
F504
F3FC
F40F
F4CA
F502
F4BB
F50B
F625
F6CE
F659
F5FD
F71E
F90D
F9D8
F92C
F8C8
F9CA
FADB
FA42
F8C7
F8C7
FA7B
FB2D
F944
F78F
FA84
0295
0B0E
0F31
0F0D
0E3B
0EE5
0FCE
0F3E
0DF0
0DD0
0EC3
0E64
0B30
06AB
03A3
0306
035B
0309
0235
0207
02E3
03F8
0475
045E
041F
03DB
038B
0372
03D8
0474
048A
03E3
0334
033D
03C1
03CB
0314
02B2
0416
076C
0B3B
0DA9
0E0F
0D5C
0D16
0DED
0F17
0F29
0DD6
0CAC
0D70
0F76
0F64
0A61
0197
F9BA
F6A8
F7E9
F9E1
F9F1
F89C
F7C2
F814
F8CA
F90E
F8A5
F78A
F5DE
F45F
F412
F512
F622
F613
F544
F50C
F5C6
F649
F5A5
F475
F3F1
F453
F4D8
F507
F516
F52A
F50C
F4CF
F505
F5CC
F63A
F596
F4D3
F5B2
F84A
FA89
FACD
F9E5
F99B
FA01
F9AD
F862
F7D5
F8FF
FA25
F928
F75E
F907
002D
096E
0F53
1018
0EB0
0E57
0EFD
0EC9
0D96
0D19
0DE1
0DED
0B37
06A8
0349
02C6
03DA
045C
03CB
034A
039D
043A
043D
039C
0304
02E7
032F
039D
0409
043B
03FD
0383
0362
03DF
0470
043D
033D
028D
0383
0673
0A52
0D74
0EB9
0E4D
0D73
0D64
0E11
0E4A
0D5B
0C51
0CEF
0F1C
0FF0
0C36
040E
FB68
F67C
F61C
F7CA
F8DD
F8DE
F8E1
F98D
FA5E
FA87
F9C6
F85B
F6AF
F551
F4CF
F532
F5BF
F5B1
F50A
F46E
F44B
F47C
F4C7
F53D
F5EC
F67A
F679
F603
F5A0
F58F
F58C
F56D
F56F
F5B3
F5CE
F575
F543
F62D
F818
F9A4
F9C3
F910
F8DF
F95F
F995
F93A
F97A
FB00
FC34
FAEC
F80B
F7D6
FD83
0705
0E9C
10AB
0EE0
0D3A
0D44
0D81
0CE0
0C9A
0DE0
0F27
0D8D
08B9
03CC
01DF
02AA
0397
035C
0312
03DF
0501
04F8
03CD
02F3
0320
0373
031A
02A9
031C
042A
049E
0425
03C4
0431
04A9
0414
02E7
02FB
056D
093E
0C5C
0D9F
0D6D
0CE5
0CDC
0D59
0DA8
0D16
0C01
0BE3
0D82
0F1D
0D47
0672
FD5C
F709
F612
F87B
FA57
F9DC
F84E
F79A
F816
F8AC
F865
F749
F614
F57B
F5AD
F62C
F630
F577
F4B4
F4CD
F5A1
F617
F58D
F4B6
F49C
F53A
F5AD
F587
F53B
F535
F538
F50D
F52B
F5FD
F6C3
F647
F4CF
F457
F635
F927
FAC2
FA6C
F9CA
FA29
FAC0
FA42
F93F
F96C
FAB7
FAE5
F8FB
F7D6
FB84
0418
0CB4
108B
0FB3
0E08
0E09
0EA3
0E18
0D24
0DA0
0EFC
0E2A
09AF
042F
019C
02A0
0442
0408
02CA
02BB
03EB
0467
0354
0243
02DD
0473
0508
0427
0358
03BC
047E
0459
0398
0381
042F
045E
0387
0330
0544
098A
0D89
0F06
0E1C
0CB9
0C89
0D8B
0E6B
0DE2
0C2B
0B21
0C63
0EDE
0EDD
098D
0085
F8E8
F687
F856
FA2A
F988
F7B1
F719
F831
F95C
F93C
F7E8
F62B
F4A3
F3D0
F40E
F50B
F5AC
F530
F43C
F42F
F564
F6BF
F719
F67C
F59B
F4DD
F461
F483
F565
F63D
F5F8
F4C7
F43B
F53F
F6AC
F6C4
F5B7
F585
F72C
F939
F9DE
F96D
F993
FA94
FAF5
FA10
F965
FA43
FB4F
FA4F
F848
F98F
008B
09D3
0F54
0F06
0CA7
0C8A
0E95
0FA6
0E9E
0D99
0E1A
0E44
0B82
069B
032C
032D
04AC
04B7
0316
01FC
02A6
03EE
044F
03E0
0392
0384
0331
02CF
032E
0438
04A6
03C6
02A8
02C1
03C8
0402
02CA
01DB
0369
077E
0BDA
0E33
0E1E
0CFD
0C95
0D9E
0F2A
0F81
0E0E
0C79
0D16
0FAD
108A
0BF7
02C9
FA50
F721
F8A5
FA8D
FA08
F832
F793
F898
F977
F8D4
F73F
F5FF
F574
F52E
F4EE
F4D5
F4D2
F4A2
F45D
F46E
F4D9
F516
F4CB
F46B
F4A7
F57C
F639
F664
F63B
F628
F630
F622
F5FD
F5CE
F567
F4C2
F489
F59F
F7E0
F9DB
FA5A
F9BF
F95D
F998
F99F
F91B
F91A
FA61
FB8A
FA75
F7DB
F7F7
FE16
07F8
0F5D
107D
0DBB
0C1D
0D63
0F2E
0F53
0EC7
0F42
0FC5
0D92
0865
038C
0206
030D
03B0
02DF
0229
02D4
03F3
0415
0380
037D
0422
0433
0349
029C
030F
03C1
0377
029F
02A0
0390
0402
034C
02CC
043D
0776
0AB0
0CAE
0DAC
0E44
0E7F
0E6C
0E7E
0EA7
0E10
0C99
0BD1
0D04
0E78
0C65
055B
FCBF
F79F
F772
F928
F96A
F837
F79D
F854
F914
F8C9
F7DE
F71F
F681
F5A8
F4E6
F4EF
F5B2
F64A
F61C
F57F
F505
F4C6
F4A9
F4DE
F56F
F5DC
F5B1
F54A
F558
F5C9
F5DB
F552
F4ED
F53C
F59E
F522
F436
F46B
F65C
F8A8
F9AA
F983
F985
FA05
FA01
F918
F8A3
F9E1
FBC0
FBE5
FA25
F9AF
FDB4
0558
0C37
0F0C
0EB4
0E3A
0EDE
0F5E
0EBB
0DFF
0E70
0F0B
0D63
0901
0494
02FC
03EF
04BA
03EE
02E3
0349
0486
04AC
0359
0245
02C2
03F4
042C
0350
02B7
02FD
0333
0291
01D9
0236
0362
0407
03D7
042C
0658
09E0
0CFC
0E6B
0E51
0D8A
0CD0
0C8C
0CC6
0D01
0CB1
0C2F
0C7C
0D6D
0CBE
0820
005A
F962
F6AB
F7CE
F97E
F975
F874
F85A
F966
FA1F
F96F
F7BA
F607
F4E1
F460
F497
F56B
F63F
F653
F59D
F4CD
F476
F477
F477
F485
F4F0
F5BB
F681
F6D6
F67F
F589
F471
F413
F4D4
F5EC
F600
F4E0
F424
F564
F810
F9E9
F9D3
F912
F947
FA1C
FA18
F941
F94B
FACB
FBC5
FA6F
F8B3
FAE9
027A
0B65
104D
101C
0E3A
0DBD
0E3F
0DF8
0D1E
0D6C
0ED2
0EB7
0B51
065E
0356
0364
047F
0466
0332
028A
0322
0419
046E
043C
0420
042B
03EF
0361
0303
032E
03A0
03EF
040B
0407
03BE
0312
0299
0396
06C5
0B18
0E33
0EB1
0DA1
0D49
0E5A
0F35
0E49
0C7A
0C29
0DAF
0DFE
09C1
018E
F9E4
F6AD
F7A8
F990
F9F5
F912
F865
F8A0
F941
F972
F8BC
F747
F5C7
F519
F578
F619
F60E
F588
F586
F633
F66F
F578
F432
F40D
F50E
F5D9
F591
F4D8
F4B3
F529
F577
F54D
F50F
F500
F502
F53B
F634
F7E2
F961
FA0B
FA2F
FA2A
F9AB
F890
F7CD
F854
F95C
F940
F861
F9DA
FFDD
0826
0DD6
0EEC
0E0A
0E3E
0F1E
0E98
0D07
0CEA
0EC5
0FAC
0CF1
07CF
03E7
02E2
032E
0312
02E9
0397
0464
0408
02F1
02C0
03C4
0481
03E7
02D0
02A1
0342
0369
029B
01F6
0292
03DB
044A
0381
0301
04B0
08C7
0D46
0F75
0E7B
0C66
0BFB
0D83
0EB8
0E29
0D50
0E20
0F52
0D08
05B5
FCEB
F7F8
F827
F9FE
FA07
F887
F7D5
F8AD
F9C5
F9F9
F944
F7E7
F610
F47C
F43E
F556
F652
F5FC
F4F8
F4D0
F5AD
F62E
F5A0
F507
F55F
F60D
F604
F586
F58B
F629
F69C
F69B
F688
F669
F5D3
F510
F569
F776
F9DC
FADA
FAA3
FAC5
FB56
FAC3
F8CC
F7A1
F8A2
F9EC
F94E
F893
FC0C
048B
0D25
1085
0EFB
0D46
0E19
0F88
0F3B
0E38
0E99
0F84
0E19
09D1
0571
037F
0386
03A6
034B
0338
039B
03AC
0332
0308
0393
03E6
0341
0267
0269
02E9
02C9
0213
01EB
02BD
038B
0353
0278
026E
0439
0787
0B01
0D3C
0DA3
0CF1
0CB4
0D9A
0E73
0DDF
0CB9
0D38
0F0D
0E55
0810
FE9E
F7E3
F6F4
F93A
FA4A
F8FF
F78B
F780
F7E7
F779
F6B0
F692
F6B8
F613
F4D8
F436
F48D
F51C
F55C
F598
F609
F642
F5ED
F57D
F590
F5F1
F5F2
F59D
F5A8
F629
F664
F62D
F646
F6DB
F6DD
F5CC
F50F
F638
F89C
FA05
F9A1
F8DD
F904
F978
F924
F89A
F907
F9BA
F906
F804
FAC1
02F7
0C76
112C
100C
0D97
0DBE
0F92
1015
0F17
0EF3
1025
0FE5
0C1E
06CE
03AD
03A0
0461
040E
0337
0330
03F3
0474
0434
03A0
032A
02BE
0245
0218
028D
0358
03D2
03B9
034C
02EE
02DF
032E
03C0
04BC
06CA
0A3F
0DEA
0FAF
0EF0
0D84
0D80
0E8A
0EA3
0D5E
0CCF
0E34
0EF2
0AF9
0236
F9B9
F655
F78B
F912
F855
F6A9
F664
F79C
F894
F83B
F724
F652
F60D
F61B
F646
F649
F5D5
F50F
F49D
F4BB
F4E7
F4CC
F4EF
F5B5
F676
F640
F54E
F4CC
F53B
F5D8
F5D6
F57D
F583
F5C3
F59E
F55C
F613
F7D9
F94B
F96E
F900
F912
F960
F91F
F8B7
F928
F9FB
F98A
F807
F8B7
FE73
075F
0E1E
0FB2
0E69
0E23
0F68
0FF2
0EEC
0E2D
0EEC
0F5A
0CEA
0803
03D1
0285
0324
0388
0344
0367
042B
0462
034A
01D3
0187
02C1
046A
053C
04F6
043A
03AB
0360
032D
0315
0326
033D
034C
03D6
05C1
0933
0CD0
0EA8
0E4C
0D6C
0DC0
0EC2
0E94
0D1E
0CBD
0ECA
10A4
0DDC
0586
FC03
F6C7
F6F6
F923
F9CC
F8AD
F79B
F797
F810
F846
F811
F780
F6A1
F5C8
F567
F56B
F54A
F4E1
F4D8
F5BA
F6F4
F752
F674
F545
F4CD
F51B
F5AA
F61D
F640
F5E3
F534
F4D8
F520
F575
F538
F4EB
F5B3
F79E
F939
F960
F8C7
F8D7
F978
F957
F850
F800
F938
FA63
F9F0
F972
FC61
0387
0B43
0F56
0F5B
0E57
0E79
0F14
0EF4
0EB5
0F69
1017
0E74
0A11
0557
02EB
0305
03DE
0415
03BD
0361
0303
027C
0224
0270
0323
0391
0378
0335
031A
0319
0316
0334
038E
03E4
03BF
031A
02E4
0473
081B
0C4C
0EB7
0E8D
0D60
0D4E
0E72
0EE5
0DA0
0C62
0D69
0F9C
0EC5
0864
FF2F
F87E
F6DA
F832
F93A
F904
F8B3
F8F6
F92E
F8D4
F83C
F7A0
F698
F532
F492
F574
F6C5
F6D4
F58D
F483
F4BE
F588
F5B5
F54C
F538
F5B3
F602
F5BB
F55E
F55C
F561
F51E
F4F8
F545
F59C
F592
F5B0
F6C0
F872
F998
F9B2
F96E
F96B
F95B
F8F7
F8EC
F9B6
FA1F
F8BE
F725
F971
014C
0AC7
1015
0FCF
0DC7
0DBC
0F3C
0FA9
0E8D
0DE6
0E8E
0E90
0BFD
07D0
0495
0341
02CA
0253
0237
02CD
037D
0393
0339
030C
0327
032A
0317
0362
0404
043C
039A
02C0
027C
02B4
02B9
027A
02BA
0444
0729
0A8F
0D09
0DB7
0D4C
0D84
0F09
1058
0F99
0D67
0C92
0E4C
0F8D
0C0F
03BE
FB72
F7A4
F7FD
F91D
F93E
F93D
F9D4
FA14
F90E
F77F
F6B8
F6A7
F63D
F55E
F50A
F575
F57F
F4AF
F453
F587
F741
F79D
F676
F554
F52F
F57F
F591
F58D
F5C0
F5C2
F53A
F4D5
F563
F642
F616
F536
F59E
F7EC
FA0F
FA1C
F8F2
F89C
F92D
F925
F864
F87C
F9BF
FA15
F876
F7FF
FCDB
0638
0E13
1019
0E58
0D7D
0E8F
0F10
0E09
0DA5
0F41
1082
0E3F
08FF
0483
0323
038F
0398
032E
0350
03B1
0338
0221
01C0
0264
02EB
02A4
0242
028F
030F
02CE
0203
01FD
0331
0452
03F2
028C
023A
048A
08FB
0D5B
0F7C
0F08
0DD9
0DE8
0EE1
0EB8
0CF6
0BFA
0DB0
0FEF
0E0A
0678
FD6A
F87A
F8A5
FA1D
F9B8
F860
F867
F9AB
FA29
F923
F7C5
F6F8
F64A
F54A
F48F
F4C6
F576
F597
F507
F49E
F4DD
F562
F5CA
F628
F656
F5DF
F523
F548
F66D
F706
F60F
F4CC
F50C
F65C
F6A4
F56E
F4DD
F6A3
F959
FA62
F9A5
F947
F9F7
F9F5
F894
F7F1
F987
FB33
FA60
F8F9
FBE6
043C
0CB6
0FC1
0E20
0D0B
0EB6
1011
0E86
0C6F
0D50
0FEF
0F81
0A59
044B
01C7
02C8
040C
03C6
0321
037B
042E
03F7
030F
02A7
02F6
0336
031C
031E
0357
0341
02B5
025C
02BB
0354
033B
0273
0266
0496
08D1
0CE9
0E9F
0DCF
0C95
0D08
0ED2
0F98
0E1E
0C46
0CB8
0EC0
0E33
0858
FF9F
F93F
F7AF
F8DC
F98A
F8F6
F871
F8A8
F8DF
F888
F82B
F823
F7B8
F650
F4BC
F450
F519
F5EB
F5F4
F579
F516
F4FB
F50F
F53E
F56A
F55E
F51E
F50F
F56C
F5C8
F59A
F531
F54F
F5D0
F5BE
F4F9
F4CB
F61E
F80F
F92C
F965
F9AA
FA0D
F9B3
F8C1
F8D7
FA92
FBC7
FA2C
F790
F8FA
009C
0A54
0FFA
1019
0E7B
0E95
0FB5
0F71
0DE6
0D71
0EBD
0F2D
0C2D
06BE
0283
01AD
0319
044C
0422
033E
02AF
02D8
0368
03EA
0425
0417
03D1
0370
031F
02F3
02D9
02BF
02BF
02FE
0350
0352
030B
0380
0604
0A69
0E62
0F89
0E23
0CCE
0D3C
0E4D
0E2C
0D5A
0DF6
0FF6
0FDC
0A78
0150
F9B2
F73F
F891
F9CF
F949
F855
F86D
F926
F93D
F877
F78B
F6D7
F601
F4E2
F40E
F41C
F4C8
F54F
F572
F598
F601
F64B
F5FE
F537
F49B
F4A8
F540
F5D7
F60D
F5FA
F5D1
F58A
F522
F50B
F5D9
F76A
F8CA
F93C
F90F
F917
F984
F9C6
F98F
F958
F979
F964
F8CE
F944
FD34
04B9
0C6C
106D
1034
0E88
0E09
0ECC
0F71
0F4D
0E83
0CCB
0994
058E
02C1
026A
037D
0422
03E0
0392
03A9
039F
0323
02C0
0304
0394
03BB
0372
0340
034E
034A
0338
0376
03C8
0382
0326
04AA
08FB
0DE6
1003
0EBA
0CFD
0D6F
0F08
0ED5
0C7F
0B19
0CCC
0F3A
0DBA
06C6
FDD5
F7B9
F632
F763
F89B
F8CA
F872
F84F
F87C
F89B
F838
F70C
F554
F3E6
F3A3
F48B
F5A0
F5DE
F545
F4B8
F4E2
F573
F59D
F536
F4FC
F583
F646
F658
F5BE
F56A
F5C7
F608
F575
F4B6
F522
F6D3
F85F
F8BD
F897
F90F
F9DC
F9D4
F91E
F93A
FA77
FAF9
F986
F849
FAFC
0244
0A64
0F33
1037
0FDD
0FAF
0F23
0DFC
0D89
0E64
0E94
0BBE
06A4
02B0
01FF
0339
03DF
0365
0305
034F
0382
033E
035C
0461
0547
04EE
03E6
03A0
043C
0478
03BE
030B
034F
03EF
03FB
0435
0681
0B07
0F2F
1067
0F20
0DF0
0E25
0E8D
0DD1
0CBD
0D1B
0EB6
0EA6
0A3D
0248
FABD
F70F
F730
F85F
F861
F77F
F753
F861
F94F
F89B
F670
F461
F399
F3DA
F456
F4BE
F528
F57B
F57D
F542
F509
F4D0
F46E
F421
F473
F559
F5E6
F56E
F4AC
F4DE
F5E2
F63D
F54D
F481
F58E
F815
FA1C
FA8E
FA29
F9E3
F98A
F8C3
F85D
F946
FA84
FA07
F81A
F853
FDB8
069C
0DE7
1053
0F2A
0DBA
0D87
0DE5
0E2E
0E7F
0E5C
0C5C
083F
0435
02C5
03D7
04FD
0490
0359
02E8
035E
03AA
0365
0355
040D
04F1
0510
0464
03A3
0339
030D
030D
034A
039B
03DC
0491
06A4
0A10
0D3E
0E6C
0DAD
0CE4
0D7B
0EBE
0F0B
0E45
0E04
0F1A
0FB8
0CF3
0623
FE25
F8D0
F766
F7FC
F833
F7CC
F806
F926
F9C1
F8A5
F68D
F53D
F546
F58E
F519
F464
F474
F521
F560
F4F9
F4E6
F5AB
F655
F5DE
F4CC
F47B
F520
F590
F52B
F4E3
F5BA
F6EE
F6E2
F58F
F4D7
F60E
F84C
F9CC
FA0C
F9AF
F916
F84D
F7FA
F8E4
FA44
FA00
F7BA
F6AA
FAA4
032F
0B48
0EBA
0E55
0DD5
0EDF
0FE1
0F6A
0E5A
0DF1
0D4C
0A7D
05C7
0207
0175
0327
0493
0490
03E5
0374
033C
0310
032D
03A6
0401
03DE
03A6
03F3
048C
0498
03D6
02F2
027E
0259
0296
043C
080F
0CD0
0FD2
0FBF
0E12
0D56
0E33
0F0A
0E78
0D59
0D83
0EC3
0E38
095A
013F
FA1E
F760
F874
F9E9
F959
F7AB
F737
F87A
F990
F8C9
F6BE
F549
F522
F55E
F50D
F478
F46E
F4FB
F56A
F561
F542
F56C
F5B9
F5E3
F5E8
F5C2
F540
F48B
F461
F530
F645
F685
F5F5
F5CE
F6DD
F862
F925
F929
F969
FA18
FA45
F997
F92B
F9D9
FA8C
F9AB
F80F
F90A
FEB6
0708
0D8C
0FC9
0F09
0DEA
0D88
0D83
0DA2
0E01
0DEF
0C17
0843
0435
0215
0246
0356
03D4
039E
035E
0366
0386
03A4
03DF
0427
0433
03E2
0366
0302
02E0
031A
03A6
0410
03CA
0305
031A
056A
09A1
0D7D
0EE5
0E09
0D04
0D57
0E59
0E7C
0D9F
0D3F
0E2E
0EB1
0BE9
0532
FD84
F8CF
F82C
F945
F96A
F870
F80E
F900
F9E7
F92C
F727
F593
F546
F560
F4E4
F42D
F430
F4E6
F54A
F4E0
F45C
F495
F558
F5CD
F5B4
F596
F5C7
F5F7
F5E3
F5D2
F5FE
F604
F586
F512
F5B0
F778
F93E
F9F6
F9DB
F9D0
FA06
FA06
F9D6
FA05
FA64
F9D1
F82B
F7C4
FB77
031C
0AEE
0F20
0F6B
0E68
0E16
0E38
0E05
0DD1
0E04
0D8B
0AD3
0652
02BD
0229
03C1
0504
04BE
03DB
037F
0383
0348
030A
037C
0479
04FA
046F
0361
02B3
02AF
0313
0384
03A7
0342
02E2
03FA
0774
0BF9
0EAA
0E37
0C8B
0C72
0E12
0F02
0DEB
0CB2
0DCF
103C
0FA4
0948
FFB2
F87A
F69F
F81E
F917
F836
F73F
F7F0
F993
FA09
F879
F632
F4F2
F506
F56E
F557
F4DE
F47F
F466
F478
F4A3
F4D1
F4DC
F4CB
F50E
F5F5
F701
F731
F64D
F56D
F59C
F660
F662
F582
F545
F6B0
F8BC
F9A6
F951
F930
F9EF
FA6F
F9B8
F8C1
F90C
FA12
F9F0
F8D7
F9F6
FFA2
07BA
0D85
0ED6
0DD3
0D84
0E4A
0EB0
0E65
0E68
0E8E
0CEB
08B5
042D
0245
031E
0448
042D
039D
03CB
0435
039F
024F
01EE
032F
04B5
04E4
03D2
02D6
02BD
0346
03DE
040F
037C
0270
025D
04D5
0979
0DA4
0EF1
0DD3
0CDA
0D6C
0E47
0DD0
0CC4
0D48
0F76
1031
0C3B
0402
FBB0
F764
F79E
F978
FA0B
F91C
F86E
F90C
F9FC
F993
F78B
F556
F463
F4A7
F504
F4D0
F459
F412
F404
F427
F4AB
F56D
F5BA
F527
F45B
F465
F563
F65A
F688
F641
F622
F5FA
F546
F47C
F4D8
F6A0
F894
F989
F9CB
FA32
FAAC
FA96
FA2A
FA42
FAB4
FA33
F8B6
F8EF
FDB8
061C
0D78
1034
0F2D
0DA9
0D3B
0D20
0CCD
0D12
0E22
0E30
0B72
06EB
03B2
0355
043A
0421
0321
02FD
0446
057F
053A
03DB
02DC
02F3
037C
0383
02D3
0201
01C0
024C
0328
0378
02F6
02B9
0470
085C
0C7B
0E63
0DD7
0CE0
0D41
0E76
0EAE
0D68
0C4A
0CED
0E48
0D1C
0771
FF3D
F902
F798
F995
FB2A
FA54
F89F
F897
FA40
FB21
F987
F6A1
F4CB
F4AA
F4F7
F4A5
F418
F40E
F44D
F432
F3F8
F467
F55E
F5BF
F51C
F47E
F4D1
F573
F53A
F470
F491
F610
F76F
F735
F5F9
F5A1
F6E3
F88A
F949
F938
F91E
F930
F94F
F9B8
FA79
FAB1
F9A2
F8A7
FAC6
0157
09B3
0F63
1084
0F23
0E2D
0E40
0E3A
0DAB
0D33
0CBE
0AF8
0751
038D
0244
03EA
0637
06AD
0529
037E
0309
0376
03C3
03B5
03D7
0463
04BB
041C
02C3
01EC
0279
03B7
03F7
02A0
014D
025E
065F
0B28
0DEF
0DFC
0CFF
0CD0
0D7B
0DCE
0D49
0CD4
0D5C
0E3F
0D6E
094B
0281
FBDB
F811
F78E
F87A
F8EC
F8C7
F928
FA42
FAA4
F90A
F668
F518
F5FC
F757
F70A
F524
F393
F3A1
F4B2
F581
F5B1
F5B1
F5A2
F533
F479
F41F
F484
F540
F5CF
F625
F641
F5D7
F501
F4C7
F622
F88C
FA60
FAC7
FA97
FAE6
FB76
FB62
FAEA
FB2E
FC15
FBFB
FA66
F9EC
FDBC
0576
0CE9
105E
1020
0F1F
0F01
0EFF
0E4D
0DD0
0E78
0F1E
0D88
0969
051B
0319
0389
04AF
052D
0517
050E
0522
04F9
048D
044A
046F
04CA
050B
0517
04F3
04AB
0456
0415
03FC
03FF
0400
0408
047B
05EF
0871
0B14
0C96
0CA9
0C58
0CC5
0DB9
0E02
0D57
0D0B
0E1A
0EF4
0C84
05E2
FE06
F90D
F836
F962
FA17
F9EE
F9DE
FA3F
FA7B
FA40
F9F8
F9D4
F948
F7F3
F66B
F57D
F51A
F4B1
F43E
F44C
F4E5
F549
F4E7
F43B
F434
F4FB
F5CB
F5FD
F5C2
F5A3
F5BE
F5C6
F57C
F4E3
F451
F474
F5D5
F810
F9EF
FAAB
FABE
FAFD
FB4A
FADF
F9DE
F98C
FA75
FB3F
FAA2
FA27
FD24
044F
0BE4
0F73
0EB9
0D46
0DBB
0F1C
0F42
0E3E
0DCD
0E1F
0D31
09CA
05A5
037A
03BB
0489
046F
03EB
0416
04F5
05A6
05A5
0526
0483
03E5
0392
03E0
049E
0501
049D
0410
042F
04C0
04B5
03BD
0303
041B
0742
0AEA
0D1E
0D61
0D00
0D6C
0E77
0EA9
0D5F
0BFA
0C4E
0DE5
0DB6
094A
01E0
FB8D
F91E
F9B6
FAB4
FAD1
FAA3
FABB
FAA6
F9ED
F8F9
F868
F7FB
F6FD
F589
F4A4
F4D5
F55C
F548
F4BF
F4A4
F549
F61D
F675
F62E
F5A1
F53E
F542
F578
F566
F4DD
F456
F478
F536
F5D2
F5FF
F68A
F82F
FA31
FB13
FABB
FAA7
FB97
FC4A
FB7B
FA14
F9F0
FAEA
FAF6
F9BD
FA50
FF98
07CC
0D9F
0E3B
0C3D
0BCB
0D80
0EDE
0EAA
0E4A
0EC9
0EA0
0BDE
0757
03FD
034B
03DC
03EE
03B2
043C
0537
053A
0401
02DE
02DC
037F
03DC
0403
0491
0557
0555
043A
0316
0304
03A1
03AE
0314
036A
060F
0A38
0D6E
0E10
0D0A
0CA1
0DA6
0E7D
0D71
0B71
0B48
0DB8
0F7F
0C76
0475
FC19
F838
F92C
FB4E
FB7E
FA04
F8F5
F933
F9D8
F9DD
F921
F7F7
F6A2
F55D
F475
F407
F3EC
F40B
F473
F50E
F574
F56A
F55D
F5DE
F6AD
F6F2
F670
F5E2
F5CE
F5D0
F57E
F53F
F597
F61F
F619
F5CD
F665
F83A
FA24
FB03
FB46
FBE9
FC8C
FBF5
FA6C
F9DC
FAE5
FB94
FA77
F9CA
FD4C
0507
0C3E
0E98
0CF4
0BAA
0CDB
0E95
0E9D
0DC0
0DE0
0E6C
0CF8
08F6
04E0
0335
03AF
0448
0403
03A4
03EC
0465
044B
03C9
0394
03CB
03FF
0418
0456
04A9
049B
0410
0396
03B5
043D
046D
03EA
0374
0471
0774
0B43
0DAC
0D9F
0C4A
0BCD
0CC0
0DA6
0D37
0C77
0D41
0EE0
0DBD
078F
FECC
F8A2
F7A3
F999
FAB2
F9B8
F864
F85D
F939
F99A
F91B
F853
F7AC
F6FD
F627
F55D
F4DE
F4C1
F4F5
F535
F51F
F4B6
F472
F4A4
F4EF
F4CC
F46C
F49D
F595
F666
F63A
F59C
F5B4
F66B
F67D
F5AA
F571
F6EF
F91F
FA3E
FA40
FA7E
FB4B
FB73
FA81
F9F5
FAF8
FC02
FAE4
F8FD
FADB
0267
0B6C
0FDF
0EB8
0C60
0CAB
0EA5
0F2D
0DBE
0C9A
0CE5
0CD6
0A81
06CA
042A
0383
03A8
0393
0397
042C
04CE
04B2
03F4
036A
0385
03DB
03ED
03D7
0407
0477
04AD
0451
038C
02C7
0263
0289
0348
04CC
075D
0AB2
0D71
0E3A
0D5A
0CAF
0D55
0E2B
0D85
0BEE
0BC1
0D91
0E44
0A34
0202
FA96
F7E1
F8E5
F9D7
F8FA
F7E3
F86F
FA28
FB2A
FA84
F8E7
F761
F647
F568
F4B2
F449
F445
F4AE
F557
F5AC
F531
F459
F441
F52E
F607
F5D1
F4FD
F4A0
F4D0
F4CA
F47E
F4DE
F63C
F755
F6F0
F5EB
F64D
F85F
FA2C
FA50
F9CB
FA0E
FAAC
FA5A
F974
F990
FABC
FB1E
FA35
FADA
0002
0826
0E1E
0F12
0D8C
0D80
0F14
0F5F
0D64
0BA2
0C34
0D7D
0C3E
080D
03F7
02AA
037F
0405
035F
02CD
034E
043E
0475
03D6
0337
032F
0389
03CB
03EB
043C
04BE
04E5
044A
0358
02E1
031E
0388
03E7
04FE
0797
0B06
0D56
0D8F
0D0D
0DAF
0F10
0F13
0D4C
0C27
0D76
0F05
0C87
04EE
FC41
F768
F72F
F884
F8DA
F893
F904
F9EB
FA16
F95F
F8A4
F839
F7A3
F6C2
F62E
F61D
F5DC
F4DA
F3A1
F337
F3BC
F466
F4BD
F505
F557
F540
F4BC
F4A7
F578
F657
F643
F599
F588
F642
F6CC
F6AA
F6C1
F7F4
F9A9
FA8C
FA79
FA79
FAF4
FB35
FB03
FB36
FBDC
FB64
F930
F815
FC0C
04F1
0D6A
104C
0E1F
0BCB
0C58
0E13
0E3C
0D3E
0D59
0E72
0DAB
0976
042E
018A
0273
0477
0512
043F
0393
03CD
0436
0411
039E
0386
03E6
0449
044F
0409
03CD
03D4
03FF
03FD
0396
02CF
020D
022B
041D
07E3
0BDD
0DE0
0D53
0BD9
0B71
0C1C
0C38
0B42
0B16
0D5C
1032
0F38
0881
FF4E
F8E5
F760
F88E
F970
F94A
F916
F94A
F95A
F8EF
F86A
F804
F762
F670
F5BC
F57D
F505
F3E2
F2F2
F34D
F48D
F51A
F444
F324
F318
F40C
F4EB
F547
F5A2
F635
F671
F617
F5CC
F603
F635
F5E6
F5C3
F6C3
F88D
F9C8
F9F8
FA0B
FABC
FB6E
FB59
FB08
FB67
FBCB
FABF
F928
FAA8
0156
0A28
0FA0
0FB9
0D85
0CAE
0D2F
0CD2
0B79
0B8B
0DF0
0FC4
0DA8
083D
038D
0254
035E
03F8
036D
0326
040A
0524
0521
042A
0397
040E
04D1
04DB
041D
035A
0339
03C5
049D
053B
0524
0439
0326
0340
0576
091D
0C2F
0D3D
0CED
0CF6
0DD0
0E31
0D29
0BEE
0C6E
0E46
0E42
09B7
01DF
FAED
F7EE
F84C
F97C
F9E8
F9A7
F941
F8EB
F8C3
F8D8
F8BA
F7BE
F606
F4BF
F4CE
F599
F5CD
F52F
F4C1
F509
F538
F491
F3BB
F3C9
F481
F4A6
F3E1
F354
F3F8
F53D
F5E7
F5C1
F598
F5C1
F5A7
F527
F53D
F6BC
F8FA
FA92
FAFE
FAB3
FA21
F971
F91F
F9BA
FAC6
FADA
F9E5
FA7D
FF6E
07BA
0E89
1007
0D5B
0AD8
0AF3
0C70
0D42
0D53
0DA2
0DD3
0C49
08AF
04FE
0358
039F
041B
03E5
03A3
03F0
043E
03CB
0302
030B
0429
0530
04FA
03E9
0373
043D
0544
052B
03E8
02AC
025F
02DA
03C2
056B
0843
0B7E
0D4D
0CF2
0BE9
0C26
0D74
0DC9
0C62
0B35
0C36
0DF9
0C9C
066A
FE66
F94D
F8A6
F9E2
FA1C
F943
F919
FA37
FB5D
FB35
F9C1
F7E1
F654
F569
F515
F4FC
F4A2
F410
F403
F4FD
F63A
F642
F4B9
F2F1
F256
F2DA
F376
F3B3
F3F1
F473
F4E5
F504
F50F
F54F
F598
F5C4
F65B
F805
FA52
FBCD
FBA0
FA9C
FA25
FA8E
FB0D
FAED
FA30
F94F
F90F
FA90
FEB2
04D1
0A92
0DB0
0E0C
0D6C
0D39
0D32
0CA8
0C00
0C19
0C9D
0BF8
094E
05BC
0343
02C6
0382
043C
046D
0426
0386
02C6
0286
0353
04CD
05CB
0596
04BF
0465
04D6
0538
04C1
03DE
03A4
0434
0454
0333
0215
0343
0719
0B24
0CBB
0BFA
0B3D
0BCE
0C75
0BE0
0B3E
0CB7
0F7C
0F6C
09B8
00C7
F9FF
F81F
F920
F9A6
F8E9
F86C
F8F7
F99B
F99C
F9AA
FA68
FAF6
FA03
F7D6
F60B
F57C
F577
F528
F4CB
F4EE
F52E
F4AA
F38E
F322
F40F
F544
F540
F3F3
F2B7
F2AF
F3C3
F51C
F5FC
F616
F58D
F4F0
F4E1
F57B
F63A
F6BC
F762
F8B3
FA40
FADC
FA30
F96A
F9B4
FA8C
FA75
F958
F95A
FCB0
0310
09A7
0DB0
0EA4
0DF8
0D48
0D2A
0D53
0D55
0D1C
0CF5
0D2C
0D6B
0CAC
0A24
0664
0335
020C
02A6
0389
03B7
0395
03F6
04BB
04FA
0446
0356
0313
037E
03DB
03C5
0394
03A3
03BB
0383
032A
0326
0356
0327
02D3
03C9
0700
0B32
0DA6
0D2F
0B8A
0B3D
0C98
0DC9
0DAF
0D46
0D8E
0D1E
0971
0292
FBFD
F904
F95C
FA2C
F9E4
F988
FA3F
FB29
FABE
F94B
F89D
F936
F969
F7E2
F5CC
F551
F699
F799
F6D9
F52C
F42D
F408
F3B7
F2FC
F2DC
F3FC
F577
F603
F589
F4F0
F4B1
F47B
F430
F44D
F52B
F64A
F6E4
F6D2
F696
F6A3
F722
F82E
F9AA
FACB
FA9F
F970
F8EC
FA1C
FBB7
FB8E
F9C9
F9A0
FE04
05F1
0CFE
0FAC
0E8A
0CC8
0C8F
0D64
0DBB
0D1F
0C75
0CA4
0D6F
0D88
0BBA
0819
0444
0237
0294
0406
0496
03B5
0299
029C
039A
044F
03EB
02EC
0262
02D9
0409
0531
0590
04D2
0379
02A8
0303
03C9
0394
025A
0209
0478
08EF
0C93
0D69
0C59
0BA8
0C1A
0C8B
0C42
0C49
0D9C
0EB7
0C6D
05B2
FD88
F854
F78A
F8D7
F960
F8C1
F85F
F8D6
F93A
F8D9
F86B
F8D9
F9A0
F959
F7BB
F61C
F5AE
F60A
F60B
F586
F544
F591
F5B6
F539
F4CC
F559
F66C
F68A
F52F
F3A1
F369
F478
F574
F583
F510
F4E1
F506
F511
F4E9
F50C
F602
F7E1
FA2B
FC01
FC8B
FBBA
FAA1
FA6E
FAE8
FAA1
F940
F8F0
FC84
03FD
0BBA
0FB7
0F50
0D53
0CA3
0D86
0E61
0E2A
0D79
0D67
0E1C
0E84
0D37
09B9
0528
01A0
0092
019E
031E
03D4
03DB
03D6
03D1
0364
02B4
0282
0307
0392
039D
0396
040C
0495
0466
03CB
03EE
04E2
0504
0352
01AD
0344
0863
0D59
0E74
0C36
0A4F
0AD9
0C55
0C9B
0C2A
0CED
0E75
0D66
0786
FF12
F8D5
F742
F88F
F992
F935
F880
F857
F86D
F860
F89F
F98A
FA5B
F9D4
F7EF
F61C
F599
F606
F61D
F568
F4A1
F47E
F4C0
F4CA
F4AB
F4FE
F5D6
F658
F5B5
F43A
F318
F31D
F404
F4EE
F551
F53A
F4F6
F4C1
F4C7
F53B
F656
F828
FA49
FBD5
FC01
FAFE
FA0E
FA3B
FAFE
FAB5
F8FB
F813
FB0F
024B
0A68
0F52
0FF0
0E74
0D75
0D84
0DA7
0D4C
0CF5
0D3E
0DE8
0E08
0CC9
09E3
05F2
0282
0126
01F9
035E
03BA
032C
030A
03E2
04BB
0492
03C6
0373
03D6
0443
0481
0511
05D7
05B9
0453
0316
0385
04D0
04C1
032B
02DD
060E
0AE2
0D50
0C3E
0ACE
0BE2
0E32
0E88
0CBB
0BEF
0DA2
0E9F
0AAC
0233
FA5A
F75A
F85C
F9A4
F94C
F862
F836
F878
F86F
F879
F93D
FA22
F9CA
F80B
F669
F627
F6BA
F6BF
F5F0
F539
F51D
F4FC
F43E
F36C
F37A
F456
F4EE
F496
F3DD
F3B1
F425
F494
F4A8
F4AD
F4F6
F557
F577
F55E
F56D
F5FD
F72E
F8D0
FA37
FA77
F966
F853
F8E4
FAE7
FC01
FA81
F848
F997
0055
093B
0EB8
0E96
0BD6
0AD1
0C8B
0E9A
0ECE
0DB4
0D45
0E26
0EEF
0DDB
0A97
0670
033D
021A
02A9
035A
02EA
01C8
0196
0306
04BE
04EA
0379
021A
0214
02F3
03A4
0409
04A4
0540
050A
0405
0345
034C
034A
02D8
036A
0699
0B3E
0DF9
0D31
0B4D
0B9C
0DF4
0F26
0DCA
0C4A
0D04
0E1E
0B6F
0431
FC9A
F90C
F951
F9EE
F91C
F85C
F928
FA51
F9E9
F864
F7F8
F929
F9E9
F886
F626
F529
F5F5
F6A6
F5EC
F4B9
F49E
F57C
F5EA
F55D
F4C8
F502
F5A0
F5C9
F585
F56C
F584
F53B
F487
F442
F4F7
F5EA
F5ED
F4E6
F3F5
F41E
F563
F731
F910
FA9B
FB4C
FB0B
FA97
FAB7
FAF7
FA25
F88E
F8D7
FD78
0563
0C49
0EB7
0D6E
0C05
0CAB
0E37
0E72
0D2A
0C3A
0CFC
0E9E
0F0A
0CF9
08FF
04F4
0293
0252
0326
0382
02D3
020A
0258
039E
0485
043C
0362
02FA
0318
0328
030F
033C
03B2
03D8
0382
036C
040A
0485
03FA
0370
0524
095F
0D57
0E44
0CCC
0BEC
0CDC
0DBB
0CDD
0BA7
0C6A
0E17
0C87
05C2
FD45
F870
F89A
FA5B
FA5B
F8F7
F86F
F92A
F981
F8AD
F7FD
F88A
F93F
F853
F5FC
F44F
F47D
F576
F5AF
F524
F4E5
F531
F52A
F466
F3D1
F46A
F5C1
F67E
F61A
F568
F54A
F5A7
F5DD
F5C1
F5A0
F57C
F4FF
F434
F3E1
F4CC
F6D3
F905
FA85
FB07
FAB3
F9FC
F984
F9AC
F9F8
F976
F849
F875
FC47
0381
0ACC
0E9D
0E7B
0CF6
0C81
0D21
0D65
0CDC
0C9E
0D89
0ECC
0EB1
0C6C
08BF
052B
02E3
024E
02EF
03C8
0418
03F9
0407
0463
0476
03D8
0320
0328
03C8
0400
0384
033D
03E0
04BC
04B0
03BE
02E2
0289
0256
029A
04C9
095F
0E06
0F84
0D9F
0B98
0C0E
0DDC
0E4B
0D49
0D4C
0EF4
0EFA
09EC
010E
F996
F70E
F80A
F8FD
F8A2
F84F
F8EC
F9A2
F99A
F95D
F9AD
F9EA
F8CD
F667
F450
F3AD
F3F3
F410
F400
F469
F524
F548
F49F
F429
F4B8
F5B5
F5DF
F503
F449
F4B0
F5CC
F661
F5F3
F532
F4EE
F524
F548
F529
F536
F5F4
F76A
F915
FA51
FACB
FAB5
FA83
FA70
FA19
F8EB
F72E
F6B4
F9BF
00AB
08D0
0E5F
0FAE
0E69
0D5C
0D7A
0D8E
0C99
0B83
0BF7
0DFA
0F7F
0E7F
0B03
06D5
03C8
028B
02AA
031C
0304
025B
01F9
029D
03F3
04D4
0495
03BD
0333
0321
031C
0325
03A5
046C
04A2
040F
0396
03DB
043A
0403
042B
066A
0A8D
0DEC
0E76
0D5C
0D4F
0EAC
0F39
0DF1
0CE4
0DE1
0EC1
0B68
035D
FB4A
F7F3
F911
FA7D
F99F
F7DC
F792
F8B1
F97E
F95E
F939
F970
F918
F78C
F591
F452
F3F1
F3C1
F386
F3AA
F439
F48D
F44B
F416
F4A7
F596
F5D3
F527
F47F
F4AB
F54B
F565
F4AB
F3E2
F3F6
F4E3
F5B4
F596
F4D8
F49D
F5AF
F7AD
F980
FA76
FACB
FB09
FB1C
FA74
F90A
F7E3
F85F
FB3D
0038
0622
0B32
0DD6
0DE4
0CE0
0C95
0D59
0E13
0DF5
0D8F
0DCF
0E52
0D97
0AF4
078D
0501
03BA
0312
02A2
029C
0314
03A2
03E8
0407
0452
04BC
04D8
044F
0336
0201
0148
017F
0284
0381
03C4
039A
03CA
043B
0410
0370
0416
0737
0B77
0E17
0E15
0D0C
0CBD
0D01
0CFE
0D46
0ECC
0FF6
0D1B
0539
FC81
F85A
F978
FBAD
FB6D
F996
F90E
FA4E
FB0B
F9DC
F837
F829
F97C
FA56
F9BF
F856
F6EA
F5AC
F4CB
F4B8
F56A
F5FD
F59F
F494
F3ED
F43F
F513
F59D
F598
F53C
F4CA
F481
F49F
F514
F564
F535
F4C2
F472
F448
F40C
F3CD
F3E2
F491
F5E6
F7C0
F9AB
FADE
FABF
F9A8
F8B1
F86D
F841
F7BE
F83D
FBE2
02AC
0997
0D78
0E12
0D77
0D2C
0D0A
0CBC
0CE1
0DF0
0EFB
0EAF
0D5A
0CA6
0D15
0CF5
0A94
06A1
035D
0203
01FD
025D
0301
03FF
04D3
04D2
0417
037D
038F
03F4
03FE
038D
030C
02D5
02DE
02DA
0291
024C
02C5
0436
057F
0538
03D3
03B4
0667
0A70
0CD9
0CB7
0BE6
0C2B
0CF1
0CD8
0C66
0D23
0E29
0BFA
04FB
FC93
F7F3
F86A
FA9C
FB1C
FA04
F972
FA08
FA76
F9F1
F95B
F99A
FA16
F9C8
F8D8
F82E
F7E2
F748
F639
F565
F547
F589
F5A1
F57F
F560
F54A
F50F
F4AB
F45F
F45D
F4AC
F55A
F64D
F6E6
F675
F53C
F46C
F4A8
F534
F511
F457
F3E7
F44D
F57A
F74E
F988
FB55
FBBA
FAD4
F9EA
F9B3
F94B
F7FE
F7B4
FB9D
03CC
0BE7
0F75
0E88
0CC4
0C91
0D15
0CD2
0C4D
0CE0
0E2D
0E87
0DA2
0D20
0DCD
0DEC
0B87
0766
0443
037A
03DC
03CA
0329
02D3
0309
033A
0315
02FE
034F
03AA
0378
02CF
025E
029E
035B
03F8
03FF
03AD
03D8
04DE
05BA
0509
033A
02AC
04FE
08E1
0B95
0C20
0BFE
0C8E
0D44
0D2C
0D0D
0E22
0EFD
0C09
043C
FB91
F732
F7FA
FA49
FACF
F9B9
F8F2
F90D
F91B
F8BC
F8B6
F965
F9ED
F981
F885
F7AA
F6C9
F584
F471
F482
F58F
F665
F639
F558
F479
F3F8
F3E5
F440
F4C5
F4DB
F43D
F39C
F3EC
F4FD
F59A
F525
F45B
F417
F434
F43E
F45C
F4DC
F577
F5EC
F6CB
F8AF
FADB
FBB4
FAD8
F9BD
F996
F9A3
F8EB
F906
FD06
04FC
0C9D
0FBE
0ECB
0D57
0D50
0D9D
0D2E
0CFE
0E1F
0F6C
0EF4
0D1B
0C60
0DAD
0EA0
0C99
083B
047A
02FE
02F6
0307
02F2
030D
0348
0352
0339
0351
03A5
03E1
03CC
0399
0390
03C9
0438
04A8
0498
03C5
02DA
02D1
037D
03AE
0346
03EB
06CA
0A8E
0CC8
0CE8
0C8A
0CE4
0D49
0CF7
0CE5
0E0F
0EA1
0B23
0349
FB7A
F82C
F91D
FAA1
FA98
FA16
FA6A
FAD3
F9EE
F831
F779
F899
FA6D
FB75
FB35
F9C8
F75C
F4C9
F386
F406
F4F1
F4EE
F46C
F4A3
F575
F59D
F4B1
F3C5
F3C1
F41D
F3ED
F37D
F3D0
F4CF
F53F
F4AE
F425
F460
F4AE
F45E
F41F
F4D1
F5FB
F6A9
F726
F874
FA5C
FB71
FB2C
FAA7
FA9F
FA08
F841
F7CB
FC41
051F
0CFD
0F5D
0D89
0BF3
0C6A
0D2A
0CD7
0CA3
0DCC
0F36
0F15
0DE2
0DA0
0E64
0DB9
0A36
05DB
038B
0376
039E
02F2
0239
0239
02AC
0316
0385
0405
042E
03B9
0321
0313
0375
0396
0350
0322
0327
02EA
0286
02C0
0389
03BE
0336
03AF
067F
0A50
0CA1
0CEF
0CE9
0D96
0E07
0D7D
0D34
0E32
0E4E
0A03
01B2
FA7B
F87A
FA24
FB1F
FA0D
F92F
FA1A
FB7A
FB89
FAAF
FA65
FAAB
FA3D
F8DB
F7A8
F718
F63C
F4C9
F413
F4EF
F60D
F5E9
F52D
F56C
F65C
F639
F4AC
F387
F421
F561
F57C
F4AA
F4A7
F5BC
F63A
F542
F444
F4A8
F58A
F545
F418
F3B7
F4F2
F71F
F970
FB6A
FC54
FB95
F9FB
F958
FA2F
FAC1
F9DF
F9D4
FE2A
0664
0D5B
0F2A
0D81
0C87
0D41
0D85
0C61
0B9F
0C95
0DE1
0DBC
0D00
0DC4
0F87
0F1D
0B11
05FB
0339
02F8
030C
0276
01FD
0210
0205
019C
01A4
0296
039A
03A9
030C
02E4
0372
03C4
034E
02CE
031F
0410
04E2
0519
0459
029D
0133
024F
0673
0B1D
0D4D
0CCE
0BD7
0BDB
0C3B
0C61
0D42
0F28
0F51
0A51
012D
F987
F776
F928
FA2B
F94B
F8D5
FA0E
FB3E
FA98
F903
F8A0
F9AF
FA7C
F9F2
F8AB
F750
F5AB
F402
F3B5
F545
F6F0
F6C3
F536
F444
F495
F505
F4DE
F4E4
F5CB
F6BD
F680
F563
F4E1
F561
F59A
F49A
F33D
F2D1
F354
F3E9
F45C
F517
F63E
F7B2
F967
FB0D
FBD2
FB65
FACF
FB3C
FC01
FB34
F8E6
F88A
FD75
0640
0D96
1002
0F0F
0E08
0DBF
0D2F
0C88
0D1A
0EA0
0F15
0DCB
0CCE
0DE1
0F5C
0DE5
090B
0431
0255
02BB
02EC
0261
026F
0380
045D
041E
0344
02A4
024A
01E9
01AD
01FD
02B2
032F
033F
034A
039A
03FB
043F
046A
0443
03A1
0379
055F
0944
0CCF
0DEF
0D2F
0C7F
0C80
0C77
0C70
0D7C
0F16
0DFD
07B6
FEA8
F87F
F7ED
FA01
FA8D
F93E
F899
F97E
FA31
F97D
F88A
F8D9
F9EF
FA20
F8F5
F783
F69C
F5ED
F523
F4AE
F4B6
F484
F3CF
F39F
F4C9
F653
F698
F58E
F4C0
F519
F5E0
F5FD
F578
F525
F55D
F5B8
F5E3
F5EE
F5CB
F53F
F498
F49A
F565
F644
F6FB
F812
F96B
F9E0
F928
F8E5
FA66
FC2F
FBB1
F988
F9FA
FFEF
08A3
0E57
0EE9
0D78
0D5E
0E24
0DCC
0CB1
0CAE
0DAA
0DB9
0C8E
0C4B
0E01
0F47
0D15
0814
0426
038A
0477
0444
0306
028D
0333
039F
032F
02C6
0316
0394
037A
02F2
02AF
02D9
02FE
02E0
02C2
02DA
030A
033F
0379
0367
02D3
02A3
0461
081C
0BD1
0DAF
0DFC
0DEE
0DAE
0CD1
0C25
0D0B
0EA2
0D4B
06AD
FD81
F77F
F733
F9A8
FAB5
F9CA
F91B
F9AE
FA5D
FA37
F9DA
FA08
FA4B
F9DE
F8FB
F86A
F81C
F74A
F5ED
F503
F50A
F534
F4C4
F43F
F475
F513
F547
F528
F574
F62D
F67E
F609
F584
F5B1
F656
F6A0
F644
F5AD
F52B
F4B8
F485
F4FD
F5F0
F6AF
F72F
F82A
F9A2
FA67
F9ED
F973
FA39
FB42
FAA5
F90B
FA17
0014
0868
0DEC
0EA7
0D4F
0D09
0DAE
0D7A
0C84
0C76
0D99
0E5D
0DF1
0D85
0E18
0E57
0C15
0773
0331
0196
0233
032C
03A9
03F8
042E
03EE
0364
033E
03A0
03E2
0391
0314
0306
0346
0323
0269
01CC
021B
0338
0428
0401
02CF
01AF
0228
04E7
08E7
0C2B
0D86
0D59
0C9D
0BE0
0B88
0C3B
0DE4
0EA3
0BE3
0534
FD7D
F8A1
F7EF
F969
FA7C
FA83
FA5E
FA8B
FA9F
FA40
F9CB
F9CB
FA4F
FACC
FA7C
F8F7
F6BC
F50B
F4D9
F5D2
F6A3
F664
F583
F50A
F532
F547
F4E8
F4A3
F50D
F5D5
F647
F641
F621
F607
F5BC
F534
F4AB
F461
F470
F4E2
F590
F5F2
F598
F50E
F5BB
F828
FACB
FB94
FA95
F9F4
FAC2
FB6B
FA51
F906
FB15
0182
08FB
0D37
0D61
0C32
0C3A
0D56
0DF8
0D9D
0D03
0CC7
0CD3
0CF3
0D25
0D5C
0D86
0DA5
0D78
0C43
098A
061E
03C8
0382
0457
0486
0391
029B
02A2
033C
0367
02F8
028F
0296
02F0
0366
03D8
0413
03F7
03B4
0388
0365
031C
02D5
02E7
0323
02C8
01C5
019E
040D
0894
0C63
0D3B
0BCF
0AA8
0B49
0CF5
0DC6
0C23
0796
0131
FB57
F855
F88A
FA14
FACD
FA55
F9BE
F99C
F96E
F8FD
F8F9
F9AE
FA43
FA14
F9E5
FA9C
FB68
FA90
F805
F5D9
F5AD
F68F
F669
F4E1
F38F
F378
F3D9
F3E4
F429
F53F
F638
F5CF
F478
F3E1
F4A9
F5BD
F615
F5FC
F61E
F64A
F5FC
F596
F5D3
F640
F5BB
F4AE
F526
F7CF
FA72
FACD
F9C1
F9E4
FB79
FC00
FA4F
F92B
FC55
03A0
0AC8
0E2C
0E40
0DB0
0DD1
0E1A
0E08
0DDE
0DCD
0DB0
0D9A
0DC6
0DEA
0D83
0CE2
0D11
0E12
0E01
0B17
0651
02E8
02AB
0416
04A5
03EE
0359
0394
03C4
032E
025C
023E
02D5
0358
0346
02DA
0286
0280
02D3
0362
03AE
033B
0268
0238
02DE
0352
02EF
02D4
04B3
0860
0B90
0C3D
0AD8
09CE
0AFA
0DB9
0F59
0D39
06FA
FF2F
F9B9
F89F
FA38
FB0B
F9AC
F7E4
F7D2
F91F
F9F1
F9B2
F97E
FA08
FA85
FA2E
F9AA
F9EC
FA3F
F8F7
F61E
F3FC
F43E
F5DD
F6BA
F64F
F5AC
F567
F514
F493
F495
F553
F5D5
F54A
F473
F4B1
F5E5
F67B
F5C0
F4E4
F508
F598
F584
F512
F53D
F5DA
F5DE
F55F
F5E2
F814
FA77
FB4A
FAF6
FB1E
FBAF
FAD5
F899
F876
FD98
0663
0D9A
0FED
0ED1
0DB2
0DCF
0DEB
0D1A
0C2E
0C3A
0CF3
0D5E
0D3C
0D0E
0D19
0D44
0D88
0DBB
0D19
0AEC
07B6
0508
03E3
03B9
0364
02AE
025B
02C4
0341
0321
02AC
029D
0310
037F
039B
0385
0366
033C
0319
032B
0364
0370
032E
02E6
02D3
02C0
0280
02C0
04A8
083E
0BB5
0D06
0C29
0B36
0C15
0E42
0EF5
0BA1
0479
FCA0
F7BB
F715
F8F3
FA9A
FAC8
FA2E
F9E4
FA07
FA14
FA07
FA53
FAD2
FAB6
F9CB
F903
F91F
F96A
F894
F6A3
F524
F53F
F642
F6A6
F5FF
F544
F53B
F58F
F59D
F568
F536
F4F3
F492
F47E
F506
F5AB
F5A2
F504
F4B5
F508
F53D
F4BD
F43D
F4BF
F5DD
F644
F5E2
F646
F841
FA68
FB02
FA74
FA61
FAE1
FA69
F8F9
F99F
FF23
07C8
0E43
0F5C
0D22
0BC3
0CA2
0DE1
0DD8
0D19
0CF0
0D64
0D99
0D4A
0CFE
0D11
0D48
0D73
0D8C
0D0F
0B10
0793
042C
027E
027F
02DB
02C6
029F
02EE
0387
03F0
0414
0425
041D
03D2
036D
0355
038F
03B4
03A0
03A4
03C9
0390
02DD
0275
02EB
0395
037A
031E
0451
07B6
0B57
0C9B
0B80
0ABF
0C64
0EE9
0E97
0989
01AE
FAFE
F823
F8C4
FA74
FAFE
FA09
F8D0
F887
F937
FA14
FA79
FA51
F9C6
F915
F8C0
F96D
FAF7
FBE2
FA93
F758
F474
F3C9
F4EB
F602
F5FC
F557
F503
F547
F5C0
F5F2
F5A6
F507
F4A1
F4FC
F5DD
F640
F592
F4B6
F4F2
F5FF
F647
F558
F4BA
F5A0
F6E2
F691
F505
F4B0
F6CC
F99E
FAE4
FAC6
FAE5
FB4A
FA7D
F904
FA55
00A6
0936
0EC2
0F50
0DAF
0D49
0E47
0EAE
0DD3
0D01
0D25
0D94
0D97
0DA1
0E23
0E5F
0D95
0C79
0C2C
0C2F
0AC8
078C
044A
02EF
0363
040C
03F9
0397
036B
0347
0305
0310
038B
03B6
02F9
01F5
01B5
0247
02EE
0359
03CE
042C
03DC
02FF
02C3
03C7
04C5
0423
02C0
0395
07D1
0CA1
0E3D
0C88
0B10
0C68
0EBE
0DE5
0807
FFB5
F958
F747
F86E
FA1C
FA81
F9A7
F8B2
F883
F8FC
F977
F9AD
F9D0
F9E1
F98E
F8F8
F8E9
F9AF
FA52
F988
F769
F588
F529
F5D8
F624
F56C
F46D
F421
F49B
F541
F585
F52E
F473
F410
F4B2
F5F8
F693
F5E1
F4D6
F4B9
F558
F570
F4AF
F44D
F527
F62C
F5D7
F4B3
F4EE
F743
F9D1
FAB7
FA67
FA40
FA32
F97B
F947
FC65
0390
0B71
0FC2
0FDA
0EA6
0E7D
0EC5
0E36
0D66
0DA3
0E7A
0E52
0CF8
0BFB
0C49
0CFB
0D0E
0D0C
0DCA
0E37
0C34
07BC
03AE
028A
039A
045A
03D0
0315
0327
03A0
03D7
03F0
043B
044A
0388
0264
01FE
029E
0363
03A2
03AE
03DF
03CA
0333
02E9
0398
0458
03C0
0277
0324
0713
0BE8
0E04
0CF6
0BFB
0D80
0F82
0DBC
06E9
FE7F
F915
F818
F96D
FA63
FA23
F977
F93B
F980
F9ED
FA49
FA83
FA90
FA6D
FA2E
F9F5
F9D8
F9C1
F961
F863
F6E0
F56B
F498
F47D
F4C1
F50A
F53C
F555
F543
F4F2
F479
F421
F439
F4C7
F57A
F5E4
F5D5
F583
F550
F54E
F532
F4DE
F4CC
F568
F62A
F606
F4EB
F43F
F549
F79E
F9AA
FAA7
FB17
FB4F
FAA8
F92D
F941
FDC5
062A
0DD9
10A3
0F01
0CE1
0CD6
0DDA
0DD7
0CC3
0C23
0C81
0CE7
0CBA
0C9B
0CFD
0D34
0CD3
0CD2
0DFA
0ED8
0CE0
07DF
02EC
0123
023D
0376
0337
0285
02B7
0360
034C
028B
022E
0284
02C6
0288
0261
02DE
0394
03CC
0394
0375
0379
033C
02E2
02FC
035C
032E
02C6
0418
082E
0CDF
0EBC
0D58
0C00
0D55
0F49
0D2D
05A9
FCF4
F860
F8D9
FAE0
FB3D
FA10
F94F
F9C6
FA86
FAA3
FA4D
FA2B
FA54
FA68
FA41
FA0C
F9D8
F974
F8C4
F7F0
F727
F686
F626
F60D
F609
F5BF
F518
F467
F416
F43E
F498
F4E2
F524
F576
F5B8
F5A5
F536
F4C3
F4A8
F4EB
F549
F583
F58B
F56C
F531
F502
F542
F643
F7CC
F91E
F9C0
FA09
FA77
FAB6
FA0D
F909
F9F9
FECC
0661
0CE2
0F52
0E65
0D2D
0D70
0E3B
0E16
0D3E
0CFF
0D97
0DFB
0D8E
0CF7
0CFC
0D61
0D81
0D76
0DB1
0DA0
0BD9
0813
0411
01E9
01DF
02A0
0320
036C
03C8
03FA
03C9
037B
0359
0302
0210
0122
016C
030A
0493
04CB
041F
03CC
040E
041B
0396
031A
0316
031D
02EA
036C
05D5
09A9
0CC9
0DE1
0DC8
0DCE
0D40
09F3
036B
FC5A
F852
F853
FA2F
FB2E
FAAC
F9E6
F9DF
FA3C
FA24
F992
F948
F9B6
FA5E
FA7B
F9FA
F986
F999
F9CA
F951
F80A
F6A9
F5D5
F57A
F527
F4C8
F4AB
F4EB
F538
F540
F517
F511
F544
F580
F59B
F593
F562
F4F9
F482
F462
F4B9
F533
F578
F595
F5BE
F5D8
F598
F51A
F50B
F61B
F849
FAB6
FC19
FB9C
F9BC
F88F
FAA2
0098
07ED
0CD9
0DD4
0CC9
0C74
0D61
0E1F
0DE5
0D9E
0E26
0EA8
0DCB
0C01
0B55
0CAD
0E71
0EA0
0D7C
0D0E
0E3A
0F68
0E55
0AA2
0620
02F7
01F1
0260
0314
0340
02D2
0254
0261
02FB
038E
03B2
03AB
03F7
048F
04F1
04CD
0454
03E0
038B
0335
02D7
02A7
02E1
0361
039E
0335
0296
02EF
0513
085D
0B05
0C0B
0C5F
0D5A
0E3A
0C5E
069A
FF56
FA66
F918
F974
F94A
F8CE
F95E
FAD0
FB63
FA5B
F91F
F92B
F9FD
FA0C
F919
F851
F877
F90D
F971
F9CC
FA48
FA2C
F8AA
F662
F4FA
F516
F58D
F533
F477
F487
F56E
F612
F5E4
F585
F599
F5B9
F521
F3F1
F322
F348
F3F6
F490
F50C
F5A0
F613
F607
F5A1
F572
F5B1
F5FC
F5DC
F565
F55C
F6AD
F976
FC5F
FD58
FBB1
F98A
FA79
FFFD
0783
0CAA
0DA1
0C87
0C5F
0D9A
0E6F
0DDF
0D01
0D32
0E18
0E43
0D58
0CAB
0D71
0F01
0F8D
0E54
0C93
0BF7
0C92
0CB3
0AC3
0723
03F1
02DB
0374
0406
03B5
032D
0336
0387
0374
032C
0369
0415
0432
0368
02DB
03A8
0512
054C
0404
02D7
02ED
0377
0348
02DA
035C
046E
0479
0379
03B7
06B4
0A87
0C22
0B8F
0BB7
0D71
0D3B
07AA
FEC4
F880
F813
FABD
FBD6
FA51
F8B3
F8D5
F9BE
F9E5
F986
F99E
F9F4
F9A8
F8FA
F909
F9EA
FA68
F9E9
F961
F9B7
FA23
F928
F6D7
F4EA
F484
F4E7
F4F1
F4CA
F526
F5AA
F545
F40E
F37B
F46F
F5F4
F67E
F5EA
F570
F5B3
F5DA
F4FB
F3A2
F33C
F433
F565
F59D
F4EC
F46A
F4CF
F5B4
F62C
F615
F67A
F856
FB08
FC8B
FBBB
FA3C
FB6F
00F3
0882
0DD1
0EB8
0D08
0C14
0D18
0E8D
0EA2
0D69
0C73
0CC5
0DCE
0E54
0E00
0D9E
0DE5
0E6D
0E3F
0D37
0C5E
0C90
0D11
0C21
0927
05BB
03EC
03DD
03EE
032F
0279
02C5
0381
0386
0306
0346
0470
04E8
038F
01AA
0162
02D5
0406
03D1
034A
03A4
0434
03CB
02FD
034F
0482
048E
02D2
01B6
03C1
0805
0B30
0BEA
0C07
0CC6
0C1B
077F
0039
FA99
F905
F9B5
F9C3
F8DE
F8B6
F9D5
FADE
FAE3
FAA4
FAE6
FAF0
F9EB
F8AB
F8A6
F9AF
FA2B
F98D
F921
F9E9
FADA
FA31
F7F0
F5E2
F529
F50F
F4AF
F478
F521
F5FB
F5A6
F43F
F381
F47F
F637
F6E1
F62A
F554
F555
F5B1
F579
F4CA
F4A0
F566
F656
F670
F59F
F4CF
F4E0
F5C1
F68B
F6C3
F726
F8BB
FB09
FC10
FAB4
F8DE
FA42
008E
0934
0F83
10F1
0EE8
0C97
0BD0
0C3B
0CBF
0CD9
0CB5
0CC0
0D27
0D9F
0DAD
0D44
0CEE
0D13
0D57
0D22
0CAE
0CE1
0DC6
0DBD
0B24
06B3
0321
022C
02E7
0367
0329
02EF
02F7
02A7
01EA
01C0
02CC
0429
047A
03B8
0311
0313
032F
031F
0388
048A
04EC
03C6
022F
01FD
031B
03A8
02E8
02AF
04E7
08B6
0B8D
0C9E
0D57
0E15
0C7A
069E
FEA8
F932
F847
F994
F9F4
F91F
F8E3
F9CC
FA5D
F980
F831
F7EF
F8B5
F96B
F9B0
F9F6
FA38
F9D8
F8EA
F885
F946
FA2A
F9A0
F792
F598
F510
F5A1
F5FA
F58B
F4E5
F4B3
F4FE
F584
F61A
F6A4
F6DE
F689
F5C0
F50B
F504
F5C2
F6AA
F6F6
F67A
F5C8
F58C
F5D8
F639
F667
F68E
F6BC
F684
F5C9
F595
F720
F9D6
FB57
FA55
F8D9
FA93
00BF
0882
0DBE
0EFF
0E14
0D58
0D6E
0DB4
0DC1
0DA8
0D72
0D20
0CFB
0D3D
0D94
0D88
0D42
0D56
0DC5
0DD5
0D3C
0CD1
0D4B
0DAA
0BFA
07F1
03CF
0202
029C
03CC
043D
040F
03C9
0371
0300
02E5
036B
040B
0408
0394
0381
03E3
03E9
0355
030C
0392
03F6
0333
0205
020B
0348
03DC
02CA
01C4
0323
06B5
0A13
0BF0
0D4C
0EA1
0DB8
0835
FFA8
F8F9
F75F
F932
FA79
F991
F81D
F7F4
F8C6
F945
F941
F981
FA1C
FA54
F9E7
F981
F9A2
F9D8
F992
F929
F96A
FA42
FA7B
F91E
F6B4
F4C7
F43F
F4A1
F4EB
F4B6
F467
F475
F4D8
F530
F54B
F55D
F594
F5BE
F59C
F567
F597
F61D
F645
F5AA
F4D1
F48F
F4FE
F591
F602
F69B
F749
F730
F602
F538
F6AF
F9D8
FBB0
FA78
F897
FA5D
00FF
08FB
0DD2
0E7B
0D64
0CED
0D36
0D5A
0D42
0D6A
0DC4
0DDA
0DA8
0D80
0D3C
0C83
0BC0
0BF5
0D44
0E6D
0E5D
0DB7
0DCC
0E4A
0D3C
09C5
05C8
03C6
03E9
0432
0364
026E
02AE
03DE
0498
0454
03DE
03DA
03E7
0391
0339
0363
03B6
037F
02E0
029F
02DF
02EB
0269
0213
0292
0348
030F
0227
0256
04D2
08CB
0C79
0EC8
0F42
0D0D
0783
FFFF
F9DF
F7AF
F8B7
FA12
F9FE
F93C
F92B
F9AC
F9BC
F93E
F919
F9A7
FA33
FA2B
FA15
FAAA
FB83
FB72
FA28
F8C3
F860
F8A4
F845
F6CE
F523
F44D
F44D
F46A
F43E
F40F
F437
F490
F4B6
F4B5
F502
F5B8
F634
F5DD
F517
F4F0
F5CC
F6D5
F709
F680
F623
F643
F62E
F580
F50F
F5B5
F6B3
F696
F5C0
F669
F95B
FC0F
FBAA
F965
F9FF
0026
08C9
0E50
0ECB
0D3E
0D07
0E0A
0E4A
0D6A
0CD6
0D3D
0DB6
0D7E
0D0A
0CF9
0D05
0CC9
0CCB
0DA1
0E82
0E17
0CB4
0C45
0D4C
0D7C
0A9B
05D2
0286
023A
032D
033B
029F
02F2
0462
0558
04D5
03C7
037A
03CB
03BD
0323
02B3
02C9
0315
035A
03AE
03DF
0364
023E
015D
01A6
02C9
038E
0360
0313
03FE
06AA
0A7D
0E09
0F55
0CB6
0656
FEE8
F9E8
F8C9
FA01
FAFD
FA9E
F9A9
F92E
F938
F92C
F8E6
F8E8
F973
FA16
FA3B
F9F0
F9C5
FA13
FA87
FA95
FA37
F9F1
FA09
F9F2
F8EF
F727
F5A3
F517
F51C
F4EE
F48A
F496
F538
F5A8
F536
F452
F3F7
F454
F4AF
F4AC
F4DD
F5AD
F65D
F5ED
F4B5
F435
F51B
F641
F63F
F553
F4F4
F5A6
F66A
F68F
F703
F8D0
FB0C
FBBA
FAFB
FBF5
0149
094C
0F2C
1009
0DD0
0C75
0D68
0EDA
0EE4
0DE1
0D50
0D8F
0DC0
0D66
0D0D
0D33
0D87
0D91
0D5B
0D07
0C6C
0BB2
0BAB
0CA2
0D34
0B70
074D
032C
0160
01D0
02A1
02C7
02D0
033D
0361
02A1
01B6
01C4
02B0
036B
0389
039A
03FA
0434
03E2
0378
0396
0408
041A
03CA
03B8
03D9
0344
01D8
0125
02D6
06A8
0ABC
0D5E
0DC4
0B77
066A
FFE8
FA96
F884
F954
FACD
FB33
FAA0
FA05
F9BC
F98F
F972
F988
F9B8
F9D1
F9E4
F9FC
F9DF
F978
F93A
F9A5
FA89
FB38
FB47
FAC1
F9AB
F7EA
F5DB
F488
F491
F527
F4F3
F3FF
F3AE
F495
F582
F557
F4B7
F4F0
F5EE
F67D
F634
F5DF
F5F7
F5D0
F4F8
F46F
F554
F6E0
F717
F5A2
F46A
F4D0
F5CB
F5E1
F5B1
F6D1
F8F1
FA17
F9F2
FB32
005D
0829
0E52
1015
0EBA
0D71
0DBE
0ED8
0F83
0F62
0EAE
0DB9
0CE4
0C65
0C17
0BCA
0BB6
0C2C
0CF2
0D59
0D14
0C99
0C82
0CC8
0CFA
0CFB
0CF2
0C72
0A80
06EC
0335
014B
019A
02D0
036A
031E
02AA
02B8
0329
0351
02D3
0216
01CB
0225
02AB
02E8
02F9
0344
03D2
0437
0436
041A
0433
0442
03F6
03AD
03EE
0446
03BF
02E7
040B
0837
0C9E
0C99
069F
FE56
F8FD
F84D
F9B5
FA21
F93B
F8A4
F942
FA6B
FB37
FB76
FB50
FACC
FA10
F98B
F986
F9BA
F99A
F8FD
F855
F831
F8AD
F966
FA0B
FAA3
FB37
FB62
FA7B
F858
F5DA
F46A
F4B9
F5FF
F6C4
F661
F573
F4E3
F501
F594
F630
F647
F577
F441
F3E5
F504
F6AC
F75A
F6D0
F63A
F668
F6B1
F630
F56C
F599
F671
F653
F4DB
F3E5
F4F9
F6F9
F7E3
F848
FB26
01E7
09E4
0EE0
0F77
0DEE
0CFE
0D16
0D24
0CC5
0C91
0CD9
0D47
0D85
0D97
0D82
0D3E
0CF5
0CDC
0CCA
0C78
0C1F
0C5A
0D32
0DC4
0D56
0C86
0C97
0D6C
0D23
0A4A
05F1
02BA
0200
02B7
0319
02B4
026A
02E3
039B
03A3
02E6
024B
0288
0342
03A6
037D
033A
0313
02B8
0215
01D4
028A
039C
03C6
02ED
0287
0379
0442
02DD
0063
00D0
05FE
0C11
0CBD
0626
FD13
F7DB
F832
FABB
FBC8
FAEB
F9E7
F9BB
F9ED
F9F3
F9E4
F9DB
F999
F919
F8E4
F969
FA61
FB19
FB37
FB08
FB00
FB14
FAC3
F9D5
F8D5
F892
F926
F9B2
F938
F7A7
F5EE
F50D
F523
F592
F5D3
F5CD
F587
F509
F4A8
F4D2
F562
F5B5
F5A3
F5C7
F675
F701
F6A9
F5CF
F57B
F5D6
F5F8
F572
F526
F5EB
F6E9
F69F
F54E
F4E8
F62D
F77A
F786
F80C
FBFF
0379
0AE7
0EA5
0E76
0D06
0CCB
0E16
0FAE
104C
0F5A
0D43
0B6D
0B3D
0C90
0DC6
0DBC
0D12
0CE1
0D21
0D2B
0D1B
0D91
0E50
0E4A
0D3B
0C5F
0CDF
0E05
0DBC
0AF9
06E1
0370
01A1
0148
01DB
02C3
036A
03AA
03C5
03AE
02EE
01AD
0110
01D0
030E
035C
029D
020E
027A
0346
0390
036E
0359
0305
0220
01AB
02D1
045C
03B7
0146
014F
0662
0C6C
0C54
0472
FAF6
F6ED
F8BB
FB3A
FAEE
F96E
F98C
FAFD
FB89
FAB5
F9EE
F9E4
F9DA
F971
F965
FA1A
FAB1
FA40
F92E
F8A5
F8FB
F956
F8FA
F84F
F83E
F908
FA17
FA91
F9CA
F7B5
F552
F41F
F48C
F576
F5A7
F547
F53C
F5AD
F5EE
F5A5
F53E
F540
F5AF
F63B
F6B1
F6E7
F696
F5C8
F53F
F5AD
F69C
F6E9
F669
F624
F68F
F6C5
F628
F599
F615
F706
F76C
F841
FBFB
0326
0AAA
0EA5
0E87
0D34
0D2E
0E15
0E4C
0D97
0CEE
0CC0
0CBA
0CD2
0D56
0E0C
0E41
0DD6
0D72
0D7A
0D87
0D42
0D2B
0DD3
0EA9
0E82
0D6C
0CE9
0DAD
0E11
0BE0
0756
0334
01C6
02A4
039F
034E
022D
0185
01D2
027B
02DD
0312
036D
03BA
0382
02DF
0283
02C2
0312
02D7
025F
0279
031A
032A
0244
01BD
02C9
041B
0346
00BB
0067
04B5
0A49
0AE2
049A
FC5C
F85D
F979
FB7D
FB1F
F96C
F902
FA0B
FAA2
FA08
F975
F9E0
FA89
FA4A
F945
F898
F8CF
F960
F98C
F949
F90D
F915
F93C
F965
F9AB
FA09
FA25
F990
F82E
F66F
F52A
F504
F5D2
F6C1
F72E
F714
F6B0
F623
F599
F55A
F56D
F57E
F563
F56D
F5E0
F65F
F65D
F5F2
F5D0
F634
F677
F612
F5A2
F617
F72A
F79C
F71D
F6BF
F70E
F728
F6A9
F789
FC44
0451
0BBA
0EEC
0E22
0C75
0C2F
0D0C
0DD5
0E3E
0E98
0EC5
0E70
0DC9
0D42
0CF0
0CC0
0CEB
0D72
0DAA
0D01
0C20
0C54
0DB4
0EB1
0DFD
0C64
0BDC
0CD2
0D51
0B64
078B
0421
02C4
030C
038C
0359
029C
0212
022C
028F
0293
0231
0216
0297
0323
0306
0277
0252
02F0
03BA
0424
0459
048E
0439
0305
0213
02D0
046A
0446
01E2
0081
032B
07E8
0925
0438
FCC4
F889
F901
FAB3
FA54
F883
F7D1
F8DE
FA12
FA54
FA3B
FA89
FAEB
FAA8
F9D3
F937
F963
FA18
FAA8
FAAA
FA43
F9D1
F97C
F936
F904
F91B
F998
FA12
F9BE
F84F
F693
F5BE
F5FC
F64F
F5FD
F56B
F547
F590
F5F1
F66A
F702
F733
F67F
F558
F4D9
F561
F605
F5C5
F4DF
F468
F4D2
F591
F618
F664
F66B
F603
F5B0
F64E
F77F
F7A7
F695
F71B
FC44
0516
0CB0
0F47
0DF9
0CC6
0D9D
0EE6
0EBB
0DA2
0D3C
0DB4
0DFE
0DBD
0D88
0D92
0D61
0CDE
0CA1
0CE2
0CF4
0C41
0B4B
0B15
0BBA
0C67
0CAD
0D17
0DE2
0DEC
0BCD
07C7
03E2
01FC
023C
0352
03E2
0395
0308
02D1
02B8
0236
017F
0174
0263
036F
0395
02F5
029B
030C
03B9
03F4
03EE
041A
0439
03E4
03B9
0490
0590
04CB
0277
01D0
04FD
092F
08F1
028F
FA84
F692
F7B0
FA15
FA8D
F9B1
F99B
FA7D
FAE8
FA62
F9DC
F9F4
FA2C
F9FF
F9A9
F9A1
F9DC
F9FB
F9DC
F9AB
F991
F98F
F995
F993
F97B
F95F
F97C
F9C8
F98C
F825
F647
F587
F647
F6FD
F63C
F4B6
F443
F563
F6B5
F6D9
F5FA
F52C
F4F6
F517
F565
F609
F6D1
F706
F665
F5AA
F5AA
F63F
F696
F632
F549
F482
F48E
F580
F651
F5D8
F4D9
F64F
FC7B
05A8
0D00
0F32
0DA4
0C53
0D1D
0E82
0EBC
0E48
0E7B
0F0E
0EA4
0D1F
0BF0
0C09
0CC2
0D0D
0CE1
0CE4
0D35
0D51
0D09
0CBE
0CA2
0C63
0C05
0C46
0D75
0E56
0D17
0974
053C
029D
023F
0317
03B3
0382
02FC
02BF
02CA
02B2
0264
0256
02DA
0395
03D8
0371
02E2
02CC
0346
03EA
0453
043F
038C
029D
0276
039C
04E2
047D
02B1
0223
047E
0783
0703
01D2
FB79
F85B
F90F
FA9A
FAA9
F9E3
F9DD
FA71
FA52
F950
F896
F8D9
F97F
F9C1
F9AA
F9BB
FA08
FA38
FA2E
FA35
FA8C
FAF7
FAF6
FA4C
F93C
F876
F8A2
F9A4
FA49
F94F
F6FB
F514
F4D4
F57B
F572
F473
F3C0
F460
F5DB
F6EE
F6FE
F687
F643
F664
F6A4
F6AA
F642
F577
F4C3
F4C3
F57D
F63F
F665
F604
F598
F57D
F5CA
F648
F65B
F5B1
F576
F816
FECB
0767
0DA2
0F20
0DA4
0CA5
0D49
0DE6
0D2D
0C1C
0C2C
0CFF
0D34
0CB1
0CA5
0D7B
0E24
0DBE
0CE7
0CB8
0D23
0D40
0CDA
0CAA
0CE1
0CAC
0BC6
0B70
0CC7
0EAC
0E93
0B68
06D4
0369
024C
02CC
03A8
040E
03B2
02BE
01DE
01E3
02D8
03BC
03A6
02DF
027C
02F2
03A6
03DC
039B
036B
037A
0362
02D7
0235
0224
02BD
0356
0369
034E
03A3
0407
0315
FFF6
FBD1
F906
F8CE
FA01
FA8A
F9C0
F8CC
F8D2
F985
F9E2
F9AD
F98A
F9DE
FA3D
FA1D
F998
F947
F993
FA63
FB49
FBC2
FB65
FA3E
F911
F8C7
F977
FA2C
FA02
F92D
F8A2
F8E9
F995
F9DA
F947
F7F0
F63D
F4D8
F46A
F505
F5D3
F5CF
F4F2
F44E
F4C2
F5EC
F6A8
F67E
F5FD
F5C4
F5B8
F58A
F56D
F5BE
F61A
F5AF
F491
F40F
F511
F6B3
F738
F64F
F569
F598
F616
F5EB
F670
FA7F
029E
0B3F
0FE9
0FB0
0D94
0CCA
0DAD
0E98
0E88
0DFF
0DC0
0DCA
0DC8
0D9B
0D2F
0C63
0BA6
0BE7
0D4E
0E9C
0E88
0D5A
0C75
0C87
0CEC
0CEF
0CC4
0CF5
0D6E
0DD1
0E43
0ED8
0E60
0B4F
0641
0252
01D9
03A4
04A0
03A3
0252
0270
03A2
046A
0444
03DF
03A4
0336
028C
0254
02CF
033A
0309
02D9
0360
0421
0431
03BD
03BE
044C
0458
035D
025B
027B
0334
02C2
0072
FD7B
FB53
FA20
F955
F8F8
F953
F9FD
FA2C
F9D8
F9B1
F9FB
FA32
F9ED
F98B
F99E
FA0C
FA2E
F9C3
F951
F95F
F9CB
FA20
FA2D
FA0D
F9E8
F9F2
FA3A
FA4D
F98C
F838
F79C
F88A
FA0D
FA54
F8CF
F6CA
F5CC
F5E3
F605
F59F
F526
F50F
F516
F4EC
F4EB
F589
F66C
F6BE
F63C
F582
F556
F5EB
F6A4
F68B
F555
F407
F40E
F57C
F6A3
F619
F4BB
F4AE
F638
F6E5
F518
F387
F709
006F
0A7D
0F56
0E9B
0CB9
0D10
0ECB
0F64
0E4F
0D08
0CAB
0CF1
0D77
0E60
0F65
0F81
0E58
0D0A
0CBC
0D14
0D0D
0C9A
0C72
0CBF
0D0C
0D4B
0DDE
0E7E
0E2E
0CDE
0C25
0D25
0E45
0C9B
07E3
035D
01F3
02D9
034D
0289
022D
0335
0464
043C
032A
02A8
02FF
0335
02EB
02FA
03BE
042E
038D
02E7
03A5
0537
0592
0404
023E
021B
034E
0425
03E9
0374
0355
0290
FFF2
FC16
F913
F838
F8D6
F97C
F9A8
F9D8
FA5E
FACE
FAA2
F9F2
F947
F8E6
F8A9
F889
F8D4
F996
FA3A
FA2D
F9C6
F9E3
FA9B
FAFD
FA5A
F962
F949
FA18
FA91
F9FA
F945
F9C6
FB2F
FBB3
FA56
F81A
F68A
F5F5
F5A9
F550
F52C
F542
F528
F4CC
F4B3
F52C
F5AE
F58B
F4F1
F499
F4A9
F4B6
F4C3
F550
F623
F630
F543
F4B8
F58E
F6AF
F65F
F50B
F4EF
F69D
F790
F5CF
F3EB
F6FB
001B
0A1F
0F00
0E4A
0C73
0CE4
0EBF
0F8C
0EE6
0E4B
0E72
0E90
0E18
0DB9
0E0F
0E7A
0E18
0D38
0CD7
0D22
0D6F
0D60
0D35
0D1C
0CEC
0CBA
0CEE
0D8F
0DED
0D98
0D27
0D53
0D75
0BED
086A
04CF
0321
0338
035C
02B6
0226
02A6
03E6
04D2
04E6
0476
03EA
036B
0333
0379
03DC
0396
02A5
0224
02DB
0404
0434
034C
0299
02E6
035A
02D0
01BA
01B1
030D
03ED
0237
FE2C
FA36
F84D
F843
F8AE
F8D5
F912
F9B6
FA4A
FA29
F97B
F919
F97A
FA21
FA49
F9D9
F959
F930
F946
F96F
F9C6
FA53
FAB5
FA73
F9B9
F94C
F9A2
FA48
FA83
FA5D
FA7E
FB03
FB07
F9B5
F771
F583
F4BB
F4CF
F4F4
F4BE
F458
F421
F44B
F4C2
F53B
F57A
F596
F5EE
F689
F6C7
F63A
F58E
F5D4
F6DE
F738
F63A
F52F
F596
F6DA
F70B
F5C7
F4EF
F5C1
F692
F54F
F3A2
F62F
FEC1
0917
0F2A
0F9B
0E2D
0E5A
0F9B
0F92
0E02
0CDE
0D25
0DB0
0D65
0CE8
0D3D
0DF6
0DFB
0D52
0CD7
0CB4
0C5F
0BEE
0C31
0D3C
0DE7
0D63
0C8B
0CAF
0D8D
0DC6
0D2F
0D22
0DF0
0DAA
0AAB
0654
03A1
0372
03D2
030A
01DD
01FE
035D
0447
03EA
0333
0307
02ED
0252
01EB
02B1
042A
04E0
045F
038C
031F
02CE
024D
0231
0305
0411
0411
0323
02CA
0397
03D2
0177
FCFB
F903
F770
F7B8
F841
F87E
F917
FA63
FB90
FB8D
FA62
F92F
F8E8
F96D
F9F0
F9F1
F9AD
F9AB
FA14
FA8F
FAB1
FA79
FA32
FA09
F9FE
FA2C
FA9C
FAE4
FA6F
F96F
F8FC
F9C9
FB03
FB04
F93C
F6E4
F596
F592
F5CD
F57D
F4EE
F4B9
F4E2
F511
F53F
F598
F604
F633
F605
F592
F501
F493
F496
F505
F561
F543
F4F4
F50A
F576
F577
F4E3
F4B6
F595
F646
F543
F3DF
F615
FDDA
07D2
0E37
0EDF
0CE5
0C5B
0DCD
0EE2
0E46
0D3B
0D50
0E31
0E97
0E3B
0DCF
0DB9
0DD6
0E16
0E6B
0E66
0DB0
0CCD
0CA5
0D3E
0DB2
0D88
0D76
0E23
0ED5
0E63
0D2E
0CCA
0D59
0CD0
09C1
05B6
0377
038F
040B
0366
0242
01E5
0235
0237
01EB
023C
0331
0392
02C9
01FD
0262
036F
03C6
035E
035E
041E
048F
03E6
02DE
0297
02E3
02B9
020F
0219
0343
03EE
0232
FE62
FAD9
F95B
F983
F9E5
F9F4
FA2F
FAE1
FB68
FAFB
F9D0
F906
F961
FA6B
FB0A
FAC6
FA27
F9EA
FA28
FA69
FA5F
FA2C
FA02
F9C5
F95E
F922
F97C
FA27
FA6E
FA38
FA4B
FB22
FBFA
FB91
F9A4
F734
F577
F4DE
F51E
F5AE
F608
F5C9
F516
F4AA
F509
F5B2
F5B6
F520
F4E8
F560
F59B
F4E9
F415
F44C
F550
F5D3
F569
F516
F591
F611
F5A3
F4DC
F4E0
F51F
F407
F267
F41A
FB9A
0605
0D72
0F25
0DDA
0D9E
0F08
0FB7
0E72
0CD9
0CCC
0DE5
0E83
0E36
0DEE
0E2E
0E68
0E17
0D80
0D3D
0D94
0E64
0F44
0F97
0EEE
0DAC
0CF2
0D65
0E42
0E42
0D52
0C87
0C33
0B0E
0813
045C
0221
0215
02CD
02B9
01F0
018C
01FD
029A
02BF
0288
0260
0260
0285
02F2
0390
03CA
0330
0229
0188
019C
021E
02CF
03A9
0466
0473
03AF
02EC
0317
03F1
0406
023B
FF03
FBDD
F9EF
F963
F9C9
FA8D
FB1B
FB1A
FAA3
FA27
F9FB
FA19
FA36
FA0E
F995
F904
F8C2
F918
F9E5
FA9F
FAD3
FA88
FA15
F998
F90E
F8CE
F962
FAA1
FB80
FB47
FA93
FA95
FB63
FBA6
FA39
F7A3
F58B
F4E4
F528
F55D
F54E
F564
F5C3
F616
F613
F5D5
F5B1
F5DF
F644
F672
F603
F521
F483
F4AA
F54A
F5AB
F585
F52E
F4EF
F49B
F423
F41E
F4F0
F5CF
F5A2
F52E
F71F
FD0F
051F
0B8E
0E76
0F07
0F28
0F15
0E15
0C9D
0C40
0D77
0ECB
0EC8
0DE2
0D8C
0E1F
0EAA
0E77
0DD7
0D66
0D46
0D5A
0DA5
0E13
0E40
0DF6
0DAC
0DE5
0E2C
0D96
0C4A
0B84
0B9A
0B07
0863
04AD
0267
0283
0365
0337
024A
0242
0376
0465
03DC
0290
01F1
0237
027E
024C
020D
0221
024D
0246
0238
0265
02A4
02B4
02C0
032B
03DF
0443
0417
03D2
03C7
0359
0184
FE37
FAA3
F846
F7D0
F8DB
FA54
FB2A
FAED
FA03
F945
F93B
F9B0
FA04
F9EC
F9BA
F9EB
FA8C
FB36
FB70
FB11
FA4D
F98F
F926
F902
F8EB
F8F2
F962
FA43
FB2D
FBB9
FBD1
FB53
F9E0
F774
F50E
F423
F510
F678
F6BA
F5C6
F4ED
F4FE
F564
F569
F568
F60B
F6FC
F734
F673
F595
F55A
F58B
F5A2
F5BE
F640
F6D8
F6CB
F62A
F5E1
F628
F5E6
F476
F378
F5AD
FC01
0458
0B6E
0F6E
109B
1022
0F07
0DF7
0D60
0D41
0D2F
0CF3
0CCE
0D04
0D5B
0D77
0D5A
0D3E
0D25
0CFB
0CF5
0D63
0E31
0ED5
0ED6
0E28
0D12
0C00
0B91
0C5F
0E1A
0F15
0D72
0937
049C
01F6
0198
0231
02A5
02EA
0340
0372
033D
02E5
02F0
0353
0362
02B9
01D0
0176
01E9
02AA
0317
02F3
027E
0236
0265
02CC
02FA
0301
0367
041A
03E2
0183
FD73
F9EE
F8E4
FA06
FB3E
FAFF
F99B
F869
F835
F8E0
F9EC
FAD9
FB1D
FA77
F94F
F87C
F87A
F90D
F9AF
FA1E
FA52
FA39
F9CC
F952
F931
F959
F94D
F8EF
F8EC
F9E4
FB5C
FBEE
FAB7
F844
F609
F50E
F533
F5A5
F5D0
F5BD
F5B9
F5C8
F5B5
F575
F55C
F5B6
F65B
F6CA
F6C6
F6A2
F6BF
F6F1
F6BE
F623
F5A0
F576
F563
F55A
F5E0
F70B
F796
F61A
F39B
F3DB
F9D9
0401
0CDC
102C
0EB8
0C9C
0C8E
0DBF
0E25
0D6A
0CE0
0D48
0DE0
0DC4
0D48
0D63
0E22
0E8D
0DFE
0CFA
0C7C
0CC5
0D4F
0DA2
0DD2
0E10
0E1E
0D9A
0CC3
0C83
0D56
0E46
0D71
09ED
0517
01AF
0158
030F
0457
03CE
025A
01B0
0249
030E
02EC
020B
0164
0184
022B
02E5
0382
03D8
039B
02D7
0240
028B
0374
03EA
035F
0295
02BC
03C1
03F5
01B7
FD63
F955
F7C5
F8C1
FA5A
FAB7
F9E0
F94C
F9F7
FB2F
FB8E
FAC3
F9E4
F9E7
FA69
FA4D
F934
F7EA
F772
F80A
F93D
FA76
FB49
FB6A
FADF
FA31
FA05
FA54
FA88
FA65
FA4C
FA61
FA09
F8C4
F71F
F622
F5E9
F591
F4A5
F3FB
F47E
F5B0
F642
F5F7
F5F1
F6BD
F755
F6AF
F587
F56F
F67F
F72C
F689
F594
F59B
F63E
F612
F503
F4A1
F5A0
F65D
F51F
F33A
F47D
FB0B
0494
0C41
0F18
0E35
0CEA
0D47
0EA9
0F43
0E69
0D16
0C90
0D02
0D9E
0DCE
0DE0
0E56
0EF3
0EF0
0E1E
0D38
0CDC
0CC6
0C68
0BE7
0BE4
0C72
0CEC
0CE7
0CD8
0D57
0DED
0D25
0A19
05C2
0260
017F
029F
03D5
03A7
0265
01A7
026C
03DF
0456
035F
022D
01F9
0293
0305
02FA
02D5
02B7
024E
01B9
01CE
02E1
03D4
0368
0246
0263
040D
04CA
0227
FD04
F8D9
F7EA
F93D
FA67
FA67
FA0E
FA3C
FABD
FAE2
FA78
F9C5
F918
F8CF
F942
FA31
FA9F
F9E8
F8BB
F880
F9AB
FB3B
FBDF
FB42
FA20
F95A
F943
F9AC
FA46
FAC8
FAF7
FAB8
FA1B
F92E
F7FD
F6BE
F5C4
F525
F4B5
F466
F469
F4C0
F517
F54E
F5BE
F692
F72E
F6C2
F56E
F45D
F46F
F53D
F5CB
F5DD
F5FD
F648
F636
F5C0
F5D4
F6E6
F7C5
F702
F567
F5FC
FAEF
02F6
0A3D
0DEC
0E53
0DBC
0DC0
0E2F
0E2D
0D9A
0D1A
0D20
0D5F
0D3E
0CB5
0C76
0D07
0DF1
0E38
0DA3
0D06
0D1D
0DA4
0DEA
0DE3
0DFE
0E21
0D92
0C35
0B43
0BF0
0D79
0D6E
0A52
057D
01D0
00E6
01FA
033D
03A1
0350
02F7
02FB
0339
036C
0392
03D4
042F
0463
0451
0430
042A
03E2
02D5
0157
00B8
01B6
0335
0379
029D
0290
03FE
048D
0185
FBCD
F79E
F7D8
FABD
FC4B
FB07
F916
F8C0
F990
F9BE
F90A
F8CC
F99A
FA67
FA3D
F99C
F988
F9F3
F9FA
F975
F95B
FA4A
FB6D
FB7C
FA6E
F981
F988
FA03
FA0B
F99E
F974
F9C3
F9CF
F8E0
F741
F5F7
F58C
F590
F56B
F537
F568
F5E6
F608
F58F
F512
F528
F59E
F5D3
F5AF
F5B9
F63B
F6C7
F6D5
F67A
F620
F5CE
F54E
F4E9
F542
F636
F699
F5D2
F542
F749
FCC6
03F7
09FD
0D2F
0DF6
0DCC
0DD5
0E53
0EDA
0EDC
0E31
0D53
0CE3
0CEC
0CED
0CB4
0CB7
0D4A
0DF8
0E12
0D9E
0D36
0D18
0CFA
0CC5
0CEA
0D8E
0DE7
0D22
0BD8
0BAD
0D14
0E26
0C88
0843
03EC
01F3
025D
0359
0388
0323
0303
0342
033F
02C6
0277
02CF
0341
02E1
01D4
014D
01F7
02EB
02D7
01F3
01D9
0327
043A
0353
0179
0180
03DD
0515
01AB
FADE
F5D1
F5E0
F920
FB30
FA68
F8EA
F907
FA56
FAF9
FA79
FA00
FA49
FAA7
FA43
F965
F8FD
F970
FA36
FA9A
FA67
F9E6
F971
F933
F941
F9A4
FA42
FACC
FAF7
FABD
FA78
FA8D
FAD0
FA5E
F885
F5E6
F417
F3FC
F4DD
F57D
F593
F5B0
F612
F644
F5FB
F5B4
F608
F6B5
F6DF
F642
F591
F57D
F5E6
F647
F66F
F67B
F67A
F687
F6D0
F72A
F6E6
F5CD
F520
F6F4
FC27
0336
0961
0CE3
0DE4
0D9F
0D2F
0D38
0DDC
0E9B
0EAB
0DF1
0D49
0D77
0E1F
0E5A
0DFA
0DAA
0DDB
0E2F
0E20
0DCD
0DA2
0D9B
0D55
0CE0
0CB8
0CDB
0C9E
0BD8
0B8F
0CA1
0E10
0D9F
0A5B
05EB
02EC
025C
02FE
0329
0287
01E5
01CF
0206
022F
0261
02C0
02F6
0291
01CD
017A
01FE
02B6
02C1
0241
0236
02EF
0352
0271
015A
0205
0432
049F
0094
F9AD
F4D2
F51F
F8B8
FB4F
FAF5
F962
F8E6
F994
FA15
F9F7
F9F5
FA66
FAA8
FA3A
F98C
F949
F974
F997
F9A1
F9EF
FA8F
FAF6
FAB5
FA23
F9F8
FA62
FAE5
FB08
FAD6
FAAC
FABC
FAB5
F9EC
F80D
F5C2
F456
F478
F581
F629
F5E7
F54E
F51E
F564
F5A6
F5B6
F5E6
F669
F6E7
F6EC
F674
F5DF
F578
F54A
F539
F511
F4BC
F476
F49E
F51E
F568
F559
F5ED
F87E
FD4F
0311
080C
0B73
0D73
0E56
0E4B
0DEA
0E09
0EB9
0F12
0E6C
0D68
0D14
0D7F
0DBF
0D5F
0CF3
0D2C
0DD9
0E54
0E7A
0EBA
0F2D
0F54
0EE5
0E3E
0DBF
0D39
0C8C
0C47
0CF6
0DE6
0D67
0AA8
06BF
039C
0225
01BF
018A
0171
01D7
02A6
0349
036E
0359
0356
034B
0307
02BA
02C5
0321
0342
02CD
0228
020A
027A
02AE
0242
0205
02EC
0434
0393
FFC3
FA62
F69C
F61E
F7D9
F9BD
FADC
FB77
FB99
FADA
F96F
F875
F8A7
F97A
FA03
FA41
FAC2
FB64
FB4B
FA33
F903
F8C1
F95D
F9EF
F9F0
F9B0
F9A1
F9B8
F9BE
F9BB
F9C9
F9D6
F9DE
F9FE
F9FF
F92D
F740
F523
F42D
F496
F536
F509
F469
F473
F564
F630
F5E3
F4D3
F423
F454
F4DF
F514
F4EB
F4CD
F4F9
F539
F538
F50B
F527
F5AD
F604
F59E
F521
F629
F991
FE72
032C
0711
0A77
0D51
0EB3
0E36
0D2A
0D49
0E71
0ED1
0D8D
0C07
0BDC
0CBE
0D41
0D19
0D3E
0E1C
0ED2
0E9B
0E02
0DF1
0E39
0DEF
0D08
0C76
0C9D
0CD9
0CEA
0D82
0E8C
0E29
0ACD
05CC
025D
0213
0374
044C
0442
0453
04B0
047A
038F
0316
03C0
049F
0496
03FB
03CD
03FF
03C0
02FF
0291
02D1
0325
031F
0319
0327
0216
FEAF
F9D9
F660
F60A
F7C6
F94D
F9AE
F97F
F94B
F8FF
F8B7
F8EE
F9A9
FA33
FA04
F995
F9BE
FA87
FB16
FAD3
FA16
F989
F94E
F92E
F93A
F9A5
FA36
FA67
FA0C
F996
F9A2
FA5C
FB25
FADE
F8F3
F63C
F47A
F490
F591
F5DC
F514
F45F
F4A5
F53D
F505
F441
F450
F57F
F666
F5F0
F4F0
F4DB
F5A0
F5F7
F57C
F52C
F597
F5D9
F51E
F486
F620
FA29
FE96
01C7
046E
07EA
0BB6
0DDF
0DBD
0CD2
0CBF
0D5C
0D7F
0CF9
0CCD
0D97
0EA5
0EF8
0E7D
0DCA
0D39
0CE0
0CF7
0D9A
0E40
0E35
0D9B
0D5F
0DE5
0E69
0E2D
0DBC
0E2B
0F12
0E66
0AEE
0630
0313
02CB
03EC
0480
0429
03D0
03EB
03F8
0398
0331
0335
036B
0365
0331
0318
0307
02CC
02AD
0320
03DB
03FB
035C
0309
0385
032F
FFB9
F982
F446
F379
F693
F9EB
FAE1
FA15
F989
F9DE
FA38
FA17
F9FD
FA47
FA6B
FA01
F9A0
F9F9
FA94
FA4D
F910
F81B
F86C
F989
FA39
FA0F
F9AB
F999
F992
F924
F8A9
F8F7
FA14
FAC9
F9E9
F7B4
F5B4
F522
F5AC
F5FC
F562
F499
F4B3
F5A0
F655
F639
F5B8
F55A
F50F
F4C3
F4E9
F5CB
F6AC
F67D
F572
F4F6
F59B
F601
F4E3
F3A0
F519
F9D3
FEEE
01C1
0328
05C3
09EA
0D28
0DCC
0D2E
0D8B
0EDA
0F3B
0E19
0D09
0D4E
0E06
0DCE
0CE8
0C8B
0CEA
0D48
0D90
0E68
0FA3
0FF7
0ED3
0D77
0D57
0DFF
0DD4
0CBB
0C66
0D8B
0E3B
0C47
085B
0540
0466
0490
0405
02DA
0257
02EB
039E
0378
02A1
01E1
01B0
0211
02CD
0368
034F
029F
024F
02F6
03C5
0386
0279
0235
034C
03D9
0152
FBC3
F664
F48B
F662
F922
FA42
F9B1
F8F5
F8F9
F950
F95A
F953
F9E9
FB0F
FBD8
FB9B
FACC
FA55
FA56
FA2A
F994
F927
F94A
F96B
F8D8
F7FD
F80F
F958
FA8E
FA77
F996
F965
FA07
F9F8
F83F
F604
F516
F598
F611
F59B
F4DF
F4C1
F4F8
F4C2
F452
F481
F541
F58A
F515
F500
F60E
F726
F6BB
F547
F4E1
F635
F73C
F617
F432
F507
F9B0
FF4C
029A
03E0
05FE
0A17
0DF8
0F1F
0DF5
0CEB
0D2E
0DA4
0D2F
0C78
0CC4
0DE4
0E83
0E1C
0D93
0DB3
0E1B
0E11
0DB7
0DB2
0DFA
0DD8
0D2C
0CBA
0CFF
0D6A
0D63
0D59
0DDE
0E0C
0C0A
078A
02EF
011E
0263
0458
04C3
03D4
0331
0395
0431
0411
0355
02CE
02EA
034C
0354
02DC
026E
02A3
0358
03A0
02E1
01E5
0235
03F1
04B7
01B1
FB12
F4C3
F2D9
F59B
F99D
FB88
FB03
F9EB
F9A1
F9DF
F9E0
F9A6
F9AB
F9EB
F9E2
F971
F920
F967
F9FF
FA44
FA03
F9AA
F9A6
F9E6
FA0D
FA11
FA42
FAAF
FAD3
FA4D
F99E
F9A8
FA4F
FA3E
F875
F5CA
F43E
F4CC
F65C
F736
F6F6
F670
F61E
F5AA
F50B
F50E
F60F
F709
F6B7
F559
F467
F495
F515
F52A
F567
F676
F75C
F688
F4A4
F4CA
F8DB
FECF
02F2
0454
057A
088E
0C61
0E3B
0D99
0CA8
0D1F
0E27
0E09
0CDC
0C44
0D03
0E11
0E31
0D84
0D03
0D16
0D4D
0D3D
0D04
0CE0
0CCF
0CD2
0D0F
0D72
0D71
0CCB
0C2B
0C6F
0D35
0CCC
0A06
05D4
02A0
01E8
02E5
03AA
034A
0290
0295
034B
03A3
02FC
01F7
01B1
026C
034C
037D
033D
035C
03EC
03FF
0307
01F1
023E
03C8
0424
00F2
FAC4
F532
F39B
F60D
F981
FB04
FA26
F897
F7F3
F870
F94C
F9F5
FA64
FAB9
FAE5
FAC7
FA5A
F9BC
F91E
F8C2
F8E6
F986
FA3E
FA8F
FA59
FA0C
FA2D
FAB0
FAF0
FA7B
F9CC
F9CB
FA97
FB04
F9C6
F70F
F4A2
F409
F4FA
F5E5
F5E3
F576
F561
F585
F55C
F514
F56B
F673
F730
F6D0
F5C3
F52A
F569
F5F9
F661
F690
F643
F524
F410
F535
F9BF
FFBD
03AD
0473
04B6
0775
0C0D
0F07
0E9C
0CDC
0CB1
0E20
0ED8
0DC0
0C60
0C85
0DDA
0EA7
0E36
0D77
0D68
0DE5
0E3E
0E35
0DE7
0D4D
0C83
0C13
0C52
0CAD
0C5C
0BAD
0BCA
0CEC
0D78
0B9E
07AF
041C
02E3
0396
0445
03E1
030B
02C5
0312
032F
02AC
01F6
01C7
024D
0304
035F
0363
0360
0350
02D7
020C
01DE
030C
04B3
0468
0079
FA18
F4B5
F2F2
F483
F71C
F8E4
F98E
F9A8
F9A8
F9BB
F9E9
FA06
F9C6
F939
F8FB
F98D
FA80
FAC0
F9E8
F8CD
F87D
F90C
F9B7
F9ED
F9C3
F99A
F9B5
FA11
FA6C
FA65
F9EF
F993
F9E8
FA99
FA5B
F861
F5A7
F41A
F469
F566
F5C6
F5AB
F5DB
F63B
F601
F529
F4BE
F56E
F689
F6F6
F69C
F62F
F602
F5E2
F603
F6C9
F78A
F6DC
F50D
F504
F923
FFAF
0414
0448
0364
05B8
0B35
0F83
0F99
0D46
0C55
0DAC
0EFD
0E84
0D2C
0CB4
0D3A
0D8E
0D2E
0CC9
0CF2
0D55
0D80
0D89
0D91
0D44
0C86
0C13
0CA2
0DAC
0DFA
0D69
0D2E
0DFD
0E96
0D02
0910
04EE
02EB
0327
03E2
03BF
0303
02BD
0347
03F8
040C
0379
02D0
0281
026F
0257
0252
0296
02DA
027F
0192
0136
025C
041D
03F1
002A
FA0C
F4E8
F30A
F408
F5FF
F7AE
F8EF
F9CF
FA1D
F9E5
F99A
F98A
F98A
F967
F95C
F9BF
FA56
FA7E
FA07
F97C
F95D
F98F
F9C1
F9F6
FA45
FA78
FA5F
FA30
FA32
FA2F
F9CC
F944
F949
F9D1
F9B2
F800
F598
F45D
F4F0
F605
F63D
F5C5
F588
F5A7
F59D
F57B
F5D1
F676
F66C
F565
F48E
F500
F608
F627
F56F
F562
F64A
F674
F530
F504
F8E2
FFAB
048E
04B6
02EA
0414
0917
0DF3
0F13
0D73
0C80
0D70
0E83
0E2B
0D04
0C73
0CAA
0CFC
0D36
0DAC
0E32
0E16
0D4E
0CCB
0D37
0DF7
0E12
0D92
0D3C
0D4B
0D3E
0CEC
0CE7
0D8C
0E1D
0D53
0ABD
0744
0459
02D3
029E
0320
03B1
03EF
03EC
03F5
040B
03E0
036D
032A
0371
03DA
03BA
0309
026C
0259
029F
02DF
0313
0333
027D
FFE2
FB69
F6B4
F3C1
F349
F497
F68D
F85E
F9A4
FA3C
FA46
FA08
F9B1
F962
F945
F979
F9CB
F9CD
F964
F912
F954
F9D5
F9CE
F928
F8B7
F8FB
F96A
F94E
F8DC
F8D8
F96A
FA0C
FA78
FAF7
FB82
FB3D
F977
F6DF
F4FE
F474
F48A
F493
F4CA
F56D
F5EE
F5CB
F580
F5CD
F661
F64B
F5A2
F598
F683
F6F0
F5A4
F3E1
F405
F606
F738
F64D
F5C6
F8D2
FEB5
036B
04CC
051B
07AB
0C4F
0FC2
1006
0E90
0DCA
0E03
0DF5
0D36
0CA2
0CC6
0D29
0D50
0D6C
0DB5
0DD6
0D71
0CD9
0CBD
0D39
0DBC
0DD6
0DA3
0D5F
0D19
0D0B
0D70
0DAC
0C54
08E6
04F6
02CC
02E4
03A9
03A0
0310
0317
03C6
041B
03A9
033F
0384
03E1
0379
02AC
029B
0370
0402
0385
02C5
0326
049B
052D
02D3
FD98
F7C9
F414
F394
F55F
F7A5
F912
F965
F908
F86A
F7D7
F7A7
F817
F8E0
F965
F97C
F9A5
FA32
FAA2
FA3E
F937
F8A5
F935
FA44
FA9E
F9F4
F911
F8BB
F8F1
F95A
F9C7
F9FD
F97F
F827
F6A9
F5EC
F60A
F64C
F625
F5BE
F577
F55D
F55F
F5A1
F617
F61A
F534
F433
F480
F61A
F73C
F6A4
F554
F512
F5C9
F5D3
F50E
F5F6
FA83
00DD
04F7
057D
0573
0816
0C93
0F52
0EC1
0D10
0D02
0E8C
0F8C
0EE4
0DAB
0D58
0DED
0E67
0E3B
0DA7
0D08
0C8C
0C5C
0C80
0CC0
0CF2
0D41
0DB6
0DD6
0D35
0C60
0C57
0CE1
0C28
08E4
0488
0225
02E4
04AA
04D7
0370
027C
02F4
03AC
0358
0270
0240
02F8
0399
03B0
03F0
04C3
0548
0491
0352
0322
042C
046A
01B4
FC31
F66E
F339
F37C
F5F5
F897
FA0C
FA3A
F9C9
F95B
F91B
F8E6
F8BA
F8C1
F904
F948
F95A
F951
F952
F95E
F96F
F997
F9C9
F9BA
F946
F8C2
F8B1
F924
F9AC
F9F4
FA2E
FA99
FAD7
FA2B
F879
F696
F570
F538
F581
F5CF
F5D4
F57C
F516
F522
F5A7
F604
F5BD
F540
F557
F5EF
F60E
F561
F4F2
F59B
F657
F599
F44C
F5B2
FB3F
01F2
055A
04DC
0449
06F6
0BC8
0F05
0F1E
0DFD
0DD3
0E6E
0E67
0D98
0D15
0D59
0DD9
0E16
0E29
0E1D
0DB4
0D12
0CE3
0D6E
0E08
0DFB
0DA3
0DBF
0DF7
0D3E
0BCC
0B61
0CA4
0D6D
0B21
064B
025B
01B3
031D
03E0
0338
02A7
0331
03EC
03A8
02D1
02A2
033C
03AA
0380
0358
0390
039D
0314
02A8
0345
0456
03C7
003A
FAC8
F625
F438
F4D3
F68A
F823
F91C
F96A
F92C
F8A1
F830
F834
F8B3
F959
F9C9
F9F5
FA04
F9F5
F9A7
F93A
F924
F99C
FA2D
FA26
F98C
F945
F9F9
FB06
FB2B
FA2F
F93D
F962
FA1F
FA0E
F897
F68B
F52B
F4F9
F58E
F63C
F68C
F666
F601
F5B2
F58C
F546
F4CE
F4B1
F561
F63A
F620
F532
F4DC
F5B0
F632
F50E
F3E2
F624
FC9A
035D
05E5
0472
03B7
06E6
0BF5
0EB7
0E25
0CDB
0D14
0E3C
0EAE
0E44
0DF9
0E0A
0DCC
0D36
0D32
0DFE
0E80
0DE2
0CED
0CD8
0D77
0DA8
0D1A
0C94
0C85
0C76
0C37
0C72
0D5E
0D7C
0AFE
0674
02C6
0210
035B
043E
03D8
0322
02F5
030C
02F6
02DE
02F5
02E2
0267
021E
02C0
03D8
041E
035F
0300
03EE
04D7
035E
FEED
F976
F573
F3D8
F40E
F52B
F6A6
F820
F92F
F99D
F9A3
F998
F993
F97D
F954
F933
F93A
F98D
FA29
FAA0
FA6D
F9B5
F950
F9BD
FA6B
FA7D
F9FC
F9BD
FA14
FA52
F9DE
F94C
F9A8
FAC0
FB0A
F98F
F736
F5B0
F58B
F5F0
F5F7
F596
F542
F53F
F571
F59F
F5B7
F5DA
F629
F679
F655
F58C
F4CF
F529
F676
F6FB
F5AA
F47C
F6E0
FD34
034B
04E2
02D5
0232
0619
0C19
0F7B
0EE5
0D1B
0CCB
0D93
0DC7
0D52
0D56
0E00
0E5D
0E0B
0DB5
0DB9
0D88
0CC7
0C30
0C91
0D6B
0D87
0CBF
0C39
0CA2
0D5B
0DBC
0E0F
0E68
0D89
0A47
05A9
0256
01C0
02C7
037E
035C
0316
0301
02BF
026B
02B6
038D
03C8
02EE
0236
02C0
03AD
0355
01F4
019C
031A
0442
0246
FD32
F7EE
F4F0
F42C
F473
F573
F74C
F937
F9F9
F991
F942
F9DA
FABB
FAE9
FA59
F9C4
F99E
F9BD
F9EE
FA37
FA72
FA4D
F9ED
F9FF
FABE
FB67
FB3D
FA8F
FA2E
FA2A
F9F0
F970
F95A
F9EB
FA31
F921
F71B
F5A9
F59C
F627
F61F
F58F
F562
F5EC
F687
F68E
F626
F5EA
F618
F64E
F608
F55B
F507
F58D
F64B
F609
F4CC
F4BC
F842
FED7
047A
059C
0358
0281
0611
0BCA
0F33
0ECE
0D1B
0CD7
0DF1
0E9B
0E1A
0D49
0CE9
0CC9
0CB5
0D16
0DF8
0E82
0E1C
0D65
0D35
0D4F
0CF8
0C6E
0CA6
0DAA
0E46
0DD1
0D3F
0D85
0D98
0B6E
070E
0325
01E8
0293
02F7
0273
021D
0295
0329
0329
02DA
02A5
0245
0197
0170
0284
03CA
0388
0211
01BB
034C
0412
011B
FB50
F699
F525
F565
F524
F4CA
F621
F8E5
FA9E
FA16
F907
F96E
FAB0
FAD5
F99E
F8A8
F8E5
F97E
F984
F963
F9F3
FAED
FB51
FAF6
FAB7
FB01
FB24
FA96
F9E1
F9B6
F9D8
F9BC
F997
F9D1
F9DC
F8BD
F6AF
F545
F57A
F665
F67A
F5AE
F563
F642
F734
F6F6
F5DE
F53A
F57A
F5DC
F5BF
F569
F562
F592
F558
F479
F3E8
F562
F9D0
FFD6
0455
0528
037B
0302
0625
0B55
0ED5
0EF1
0D70
0CBF
0D21
0D65
0D30
0D36
0DB5
0E01
0DBD
0D7F
0DBD
0DED
0D72
0CDC
0D2B
0E0C
0E19
0D06
0C42
0CC8
0DAD
0DC1
0D7C
0DD1
0DE4
0BA8
0704
02C9
019D
02E0
03CD
032A
0254
02A2
0370
0398
034A
0343
034F
02DF
025E
028A
02F4
029B
0208
0310
05A3
0667
0240
FACA
F536
F458
F5DA
F63D
F592
F647
F8B5
FA6E
F9E3
F88F
F893
F9BC
FA38
F981
F8F0
F95C
F9DC
F988
F914
F99A
FAB6
FB1C
FA8F
F9F2
F9C5
F9B0
F97B
F977
F9B4
F9A6
F91C
F8E1
F99F
FA6A
F98F
F6F8
F4A2
F427
F4DE
F53D
F514
F555
F615
F643
F556
F43B
F411
F4AF
F508
F4B3
F46F
F4E3
F59C
F5B2
F524
F52A
F735
FBA1
0101
04B6
0520
0391
035D
065D
0AF4
0E0E
0E99
0E13
0E0D
0E50
0DEA
0D19
0CF6
0DA5
0E15
0DCA
0DA6
0E55
0F0F
0ECC
0DE9
0D7B
0D98
0D62
0C9B
0C16
0C6D
0D25
0D9D
0E08
0E9E
0E59
0BD4
0795
042A
0354
0412
0450
0394
02DA
02A2
026A
0208
022D
0324
0405
03D7
02FA
028E
02C2
02CB
0286
02CF
0396
02F7
FF63
FA0B
F5D1
F42A
F419
F442
F4B7
F63C
F88B
FA50
FAC6
FA74
FA2F
FA16
F9F3
F9E5
FA17
FA3E
FA07
F9B2
F9B2
F9EF
F9F7
F9D1
F9F9
FA95
FB1F
FB24
FAD1
FA8B
FA39
F98C
F8DF
F902
F9E7
FA3A
F8D2
F63F
F433
F3AC
F42E
F4BC
F4F1
F505
F531
F56D
F5A4
F5D0
F5DC
F597
F506
F496
F4C5
F57C
F5E9
F53F
F3CC
F366
F639
FC83
036D
0702
05F3
0305
0259
0564
09F8
0D16
0DE9
0DC5
0DF4
0E55
0E26
0D5E
0CB6
0CBE
0D60
0E24
0E96
0E7E
0E07
0DA6
0DAE
0E0B
0E7B
0EE0
0F1F
0EF3
0E3E
0D7B
0D6E
0E00
0DCA
0B69
0750
03BD
0286
034C
042F
03FA
0313
0283
02A2
02F5
02FE
02C5
02A3
02AD
02A6
026A
0241
027E
02CA
0205
FF2A
FA86
F5DF
F314
F296
F372
F4BC
F651
F821
F97B
F9B0
F91F
F8F4
F9BE
FAC1
FAF1
FA3F
F985
F96A
F9B8
F9F5
FA03
F9FC
F9D7
F992
F983
F9FD
FABD
FB0E
FA96
F9BE
F93A
F950
F99E
F978
F883
F705
F5B7
F53D
F5A1
F653
F6AE
F68D
F63D
F5FD
F5D1
F5C1
F5EB
F635
F657
F653
F66C
F682
F5F6
F4DD
F4D7
F7D8
FDB2
0372
05FA
052A
03E9
04F8
084C
0BBB
0D8D
0DCD
0D8F
0DA9
0E27
0E80
0E2D
0D46
0C83
0C7C
0CFA
0D4C
0D48
0D7A
0E36
0ED6
0E8E
0DC3
0DB8
0EB2
0F63
0EBA
0D84
0D53
0E1C
0DF3
0B68
0767
043F
0324
0334
02F4
0210
0172
01DD
0309
03F4
03E2
0308
024D
0247
0282
0233
0190
01A5
0284
0254
FF27
F98D
F478
F247
F28F
F350
F3C3
F4DC
F725
F95F
F9FD
F92C
F877
F8BD
F970
F9C1
F9B5
F9CE
FA29
FA63
FA31
F9B7
F942
F8FD
F8F2
F91C
F955
F969
F967
F98D
F9DF
FA13
FA10
FA05
F9CF
F8DE
F716
F56A
F4F7
F5AB
F65D
F63C
F5B0
F589
F5D2
F5F7
F5D5
F5D9
F61E
F633
F605
F61D
F686
F658
F54D
F52B
F856
FEB3
04EB
077A
0628
0404
0415
06C3
0A54
0D01
0E2F
0E39
0DF6
0E22
0EBB
0F03
0E74
0D83
0D07
0D28
0D64
0D7F
0DD2
0E76
0EBB
0E0E
0D12
0D12
0E3C
0F3C
0F03
0E31
0E00
0E3A
0D47
0A49
0674
03E7
0380
0429
0440
0357
0264
0265
0324
0386
02F3
0223
0241
035B
0417
0375
0262
0295
03D1
036F
FF65
F90F
F404
F259
F2FE
F3D3
F457
F575
F762
F8F1
F936
F8C8
F8C4
F939
F963
F910
F8EE
F96D
FA1A
FA3C
F9BC
F91C
F8D3
F8EB
F92E
F967
F97C
F96B
F953
F95E
F98D
F9C6
FA16
FA77
FA65
F92D
F6FD
F520
F4BD
F58B
F648
F63D
F5D0
F59F
F5A5
F591
F581
F5D2
F652
F668
F601
F5B6
F5B7
F576
F4F1
F5B7
F970
FF73
04A6
0653
04DF
0349
042E
0793
0B7A
0DEF
0E77
0DE4
0D69
0D9E
0E1A
0E0D
0D5A
0CCF
0D1D
0DE0
0E20
0D97
0D03
0D1C
0DB7
0E26
0E22
0DED
0DA0
0D00
0C2F
0BF0
0CAE
0D74
0C96
098B
05C5
0371
0365
0469
049E
0373
021F
0213
033E
0434
03FF
033F
0327
03BD
03CB
02C4
01E2
028D
03EC
0340
FF11
F93F
F51A
F3FC
F48A
F518
F59D
F6DC
F891
F97B
F924
F89C
F906
FA0D
FA7A
F9E3
F922
F91A
F9B0
FA2C
FA31
F9FE
F9EC
F9FB
FA00
FA0A
FA51
FACB
FB00
FA8C
F9B7
F956
F9DF
FAAF
FA7A
F8A9
F631
F4A5
F493
F526
F573
F575
F59A
F5DA
F5D3
F596
F5A0
F5EA
F5BD
F4C7
F3F1
F45D
F5B4
F671
F622
F688
F9A8
FF05
03B4
054D
0448
034E
048F
0801
0BE0
0E6B
0F23
0EC1
0E55
0E4A
0E2A
0D63
0C3C
0BAB
0C30
0D29
0DA4
0D7E
0D45
0D48
0D43
0CFF
0CC8
0CF4
0D44
0D34
0CD7
0CD9
0D75
0DBD
0C63
0939
058F
0318
027D
02F3
0329
029D
0219
02A1
0406
04F5
048C
037A
0316
0393
03DA
0345
02C0
035A
041F
029E
FDFD
F875
F505
F44A
F48A
F475
F4AD
F640
F89F
FA17
F9F7
F952
F967
FA12
FA57
F9E8
F965
F955
F992
F9C6
F9F2
FA46
FAAB
FAC6
FA63
F9D0
F9A1
FA0D
FA94
FA81
F9C6
F932
F97E
FA40
FA1E
F861
F602
F4A0
F49F
F4FC
F4FF
F529
F5FE
F6D3
F6A3
F5AD
F530
F597
F5E4
F558
F4CA
F54E
F628
F59E
F40D
F49F
F9B5
015F
06D0
073E
0471
0287
03F3
07FC
0C38
0EBC
0F1C
0E3F
0D86
0DB1
0E40
0E32
0D73
0CF0
0D24
0D50
0CBD
0C09
0C4F
0D76
0E39
0DE8
0D41
0D2E
0D65
0D04
0C32
0C19
0D09
0D89
0BF8
088A
0513
031C
02C9
033D
0384
0336
02AF
02AA
0355
03EA
038E
0285
01FC
0283
0344
034F
031B
03A6
0431
026D
FD8C
F7FE
F4F6
F4E2
F58F
F579
F57C
F6F2
F94A
FAA2
FA43
F960
F92E
F96C
F94C
F8E8
F8F8
F988
F9F5
F9FC
F9FD
FA40
FA8E
FA98
FA67
FA3B
FA33
FA3A
FA1D
F9BC
F92D
F8DA
F92D
F9DA
F9BF
F815
F5BE
F486
F4F6
F5BE
F5A2
F509
F4FA
F567
F585
F554
F5A6
F689
F6DE
F60A
F531
F590
F651
F59E
F409
F4EC
FA42
016F
05B8
0575
0372
0350
05E7
0974
0C26
0D88
0DF9
0DE9
0DC9
0DDB
0DCE
0D2D
0C6F
0CAE
0DF2
0EB1
0DD9
0C79
0C57
0D6D
0E0C
0D59
0C6E
0C9A
0D7A
0DB7
0D2B
0D0C
0DC5
0DE3
0BDF
0834
04D2
0304
02A1
02E6
0342
037B
03AD
041F
04BD
04E2
041A
02F6
0290
030C
034E
02AC
0244
0365
04DE
0385
FE24
F795
F3C9
F392
F4A2
F518
F576
F6E8
F904
FA57
FA75
FA53
FA99
FAB1
FA00
F915
F8E1
F95E
F9C3
F9C0
F9B5
F9DC
F9FB
F9DA
F991
F953
F945
F978
F9DB
FA21
FA09
F9BF
F9AF
F9C1
F921
F753
F54B
F493
F549
F5E2
F557
F479
F491
F575
F606
F5EC
F5C2
F5C9
F582
F4EE
F50E
F650
F74E
F680
F51C
F684
FC15
02C5
0634
0563
0347
0335
05DD
09A8
0CC0
0E36
0E11
0D23
0C98
0D07
0DCB
0DD5
0D21
0CB2
0CF8
0D30
0CC7
0C6B
0CE8
0DBB
0DCE
0D2E
0CF7
0D87
0DD6
0D09
0BE9
0BEE
0D0B
0D69
0B87
07FE
04AF
02D8
0269
02AA
02E6
02C9
02A7
0316
03FB
0458
039D
02A8
02C2
03C0
042C
0369
02C7
0370
03F1
0177
FBAF
F5F4
F3AA
F48B
F5B7
F5AC
F59E
F6FF
F937
FA92
FA86
FA0F
FA0B
FA33
F9FE
F99E
F99A
F9E8
FA1C
FA2E
FA56
FA74
FA1C
F94E
F89D
F89C
F95A
FA5B
FAF3
FABC
F9F8
F969
F989
F9DC
F949
F773
F577
F4CD
F587
F644
F607
F558
F53A
F5AB
F5DF
F582
F514
F511
F571
F5FA
F686
F6B2
F5F6
F4A3
F47B
F75F
FCFE
0292
0563
053F
042F
0442
061F
0934
0C5F
0E7B
0EF6
0E53
0DBE
0DD9
0E23
0DCE
0CF2
0C7C
0CE7
0DA2
0DEA
0DBC
0D92
0D94
0D8F
0D78
0D66
0D38
0CBA
0C34
0C56
0D62
0E7D
0E2E
0BA4
0788
0390
015C
0166
02B7
03A2
0343
0253
0230
0309
03A6
0332
026F
028C
035A
03A9
0342
0351
0442
0424
0096
FA29
F48F
F2C3
F400
F54A
F548
F549
F6B6
F8E2
FA12
F9D7
F960
F9AD
FA58
FA7B
FA09
F9B2
F9C4
F9E4
F9D8
F9E2
FA27
FA39
F9A2
F8AC
F83B
F8C9
F9C7
FA3F
F9ED
F980
F99F
FA01
F9AF
F830
F635
F4F8
F500
F5B3
F614
F5D3
F570
F572
F5C2
F5E8
F5B9
F586
F59D
F5D8
F5BE
F530
F4EE
F648
F9F9
FF1E
0375
0518
043A
0320
0425
0797
0B97
0DFD
0E3C
0D73
0CFF
0D46
0DC9
0DF7
0DC6
0D8C
0D89
0DA7
0DAA
0D78
0D2B
0CF3
0CF1
0D33
0DA7
0E0F
0E25
0DE3
0DA1
0DAD
0D92
0C32
0901
0510
026F
0229
033E
03E5
0381
02E9
02E0
030D
02CB
0265
02AB
0389
03F5
0382
032B
03BA
03F7
019B
FC52
F6CA
F40F
F44E
F530
F517
F4F3
F65A
F8EB
FAA4
FA84
F9AD
F9A1
FA4B
FA86
F9F9
F97E
F9A8
F9ED
F9A6
F934
F960
FA0D
FA57
F9F5
F9B1
FA2C
FAD4
FAB7
F9F7
F9A9
FA29
FA66
F941
F71E
F576
F51C
F583
F5B8
F578
F520
F500
F514
F543
F57B
F59C
F599
F5A6
F5EE
F613
F581
F4A4
F536
F8AA
FE3C
0322
0505
0421
02DE
038D
0683
0A4A
0D22
0E50
0E43
0DE4
0DB7
0D97
0D40
0CEB
0D17
0DB8
0E0A
0D8B
0CBA
0C83
0D04
0D69
0D10
0C5D
0C1B
0C6D
0CE0
0D4E
0DF4
0E62
0D3F
09CA
0555
025C
0204
0311
039E
034C
0326
03BC
0440
03CD
02D2
027B
02F7
0337
02A8
0243
0326
046F
038C
FF1E
F8F6
F481
F359
F41B
F4C0
F525
F67E
F8DB
FA91
FA62
F938
F8E9
F9C5
FA68
F9E6
F919
F947
FA37
FA9F
FA1C
F9AE
FA13
FAAA
FA95
FA26
FA45
FADC
FAEB
FA29
F996
F9F7
FA75
F99E
F777
F5A7
F563
F615
F675
F623
F5A1
F532
F4B4
F45C
F4B1
F59E
F645
F61C
F5A6
F59A
F5B5
F552
F515
F6EF
FBB8
0170
04DB
04C5
0324
02F1
0569
0960
0CBF
0E42
0E1C
0D66
0D1D
0D6D
0DC7
0DB1
0D65
0D68
0DB1
0DB3
0D54
0D36
0DAC
0E0F
0DA1
0CC3
0C81
0D04
0D4F
0CD6
0C7B
0D25
0DC1
0C14
07BB
0348
0186
0253
0341
02DF
0228
0283
0388
03C9
030D
028E
02F3
0347
02AB
0200
02AD
0411
0386
FF89
F9DD
F5D7
F4C8
F51A
F4EB
F480
F576
F81A
FAA0
FB41
FA45
F966
F99C
FA42
FA5E
F9F8
F9C9
FA00
FA17
F9C3
F984
F9D7
FA66
FA78
FA13
F9FD
FA8E
FB0D
FAB0
F9CF
F980
FA00
FA2F
F8E5
F686
F4AF
F476
F557
F605
F5D6
F52E
F4DA
F542
F622
F6C1
F688
F5A5
F50A
F56A
F642
F66C
F5DD
F662
F9D8
FF94
0457
0563
0363
01C2
0338
0766
0BBD
0E23
0E6A
0DB0
0CFE
0CB6
0CD9
0D4F
0DDA
0E27
0E05
0D97
0D34
0D18
0D23
0CFE
0C94
0C4E
0C97
0D24
0D36
0CA7
0C68
0D44
0E44
0D2C
0919
0421
017D
020C
0399
03CC
02DE
0296
0360
03C5
02D5
01C1
021C
036A
03C3
02C3
0239
0341
03EE
0158
FB7B
F5B5
F316
F358
F42F
F497
F590
F7C2
F9FF
FABE
FA35
F9D8
FA3F
FA98
FA39
F9BA
F9F3
FA93
FA8E
F9B5
F91C
F9AE
FAEB
FB97
FB40
FA93
FA4A
FA64
FA8B
FAB1
FAEE
FB02
FA60
F8D6
F6F1
F592
F51F
F543
F561
F52A
F4CF
F4B7
F513
F5A0
F5EB
F5CB
F59E
F5D5
F64D
F64A
F562
F465
F51E
F8C3
FE73
037F
0588
0498
031F
03BE
06F5
0AF2
0D7E
0DFE
0D8A
0D67
0DC8
0E10
0DE9
0DA3
0DA2
0DC5
0DAB
0D4D
0D04
0CF9
0CE8
0CA8
0C98
0D2D
0E0E
0E3D
0D61
0C7E
0CBF
0DA1
0D0F
09C9
0541
0255
0241
0380
03E7
0333
02BA
031F
0374
02EA
0246
02C2
03FC
044D
0332
0240
02D8
03B4
01FB
FCE9
F735
F42B
F420
F4BF
F472
F439
F5C2
F8A6
FAAF
FA89
F940
F8A9
F931
F9D0
F9C8
F981
F99F
F9F6
F9F3
F99B
F98D
FA09
FA8D
FA98
FA64
FA7C
FADA
FAF4
FA96
FA37
FA3B
FA44
F994
F81D
F69D
F5C3
F57A
F54B
F51E
F535
F59E
F601
F60E
F5D3
F591
F57B
F5A7
F60A
F64A
F5E4
F4FA
F4EB
F76F
FC91
01F1
04AC
042B
02B6
032E
0651
0A5D
0D15
0DC8
0D76
0D60
0DD3
0E3A
0E0E
0D80
0D36
0D74
0DBB
0D75
0CD0
0C8C
0CF2
0D62
0D38
0CBB
0CB1
0D35
0D93
0D73
0D67
0DC3
0D6C
0AD5
0663
02B3
01DF
0321
03FA
0358
027D
02B9
037C
0361
027E
0247
0341
0415
0395
02A4
02DE
03D5
0307
FEF5
F957
F55B
F441
F492
F49E
F49D
F5C6
F812
F9EB
FA28
F965
F90A
F98D
FA24
FA0A
F983
F95D
F9DD
FA72
FA7C
F9FB
F975
F966
F9D8
FA80
FAF8
FAFC
FA93
FA12
F9E6
FA26
FA66
F9FF
F8B8
F713
F5E2
F587
F5B9
F5EE
F5E6
F5BC
F59A
F57F
F55A
F53A
F544
F597
F619
F66F
F629
F54A
F4CE
F659
FABD
0099
04F2
05C0
03FF
02DB
04A7
08BC
0C7B
0E09
0DC9
0D49
0D5D
0DA9
0DA2
0D69
0D75
0DCB
0DEC
0D8D
0D07
0CE2
0D1E
0D30
0CD4
0C80
0CC5
0D69
0D9B
0D19
0CAA
0CF9
0D31
0B82
0774
0320
0152
027B
0444
0457
02E0
01C6
01FD
029F
02A8
0271
02CD
0369
033F
027A
028E
03DB
043F
0138
FB43
F5D5
F3B9
F44F
F511
F50A
F595
F7C3
FA51
FB18
F9D3
F860
F85D
F96E
FA2D
FA14
F9CD
F9F4
FA41
FA24
F9A2
F941
F956
F9C7
FA51
FAB1
FAA9
FA30
F9B0
F9BA
FA55
FACE
FA5D
F8F8
F74B
F607
F55F
F530
F54D
F584
F59B
F589
F58E
F5D0
F60F
F5FB
F5CA
F611
F6DA
F74B
F6A8
F5A6
F64C
F9FC
FFAC
0467
05D1
0440
0270
031C
06AC
0B0A
0DB7
0E04
0D4C
0D30
0DE9
0E81
0E53
0DCD
0DA7
0DD4
0DC2
0D59
0D27
0D6D
0D96
0D12
0C52
0C46
0CF9
0D63
0CE6
0C51
0CC5
0DBF
0D36
0A00
058F
029F
0252
0345
0394
0301
02A4
02FE
0346
02C4
0205
0212
02D6
0331
02AB
023A
02B3
0304
0101
FC32
F6ED
F412
F415
F504
F540
F553
F693
F8D2
FA56
FA1D
F920
F8EC
F99D
FA02
F97D
F8E0
F935
FA45
FAE1
FA6C
F984
F91D
F969
F9EB
FA3E
FA66
FA70
FA48
F9FD
F9DD
FA0C
FA1C
F957
F791
F57F
F431
F42C
F506
F5EE
F65C
F65B
F633
F600
F5AE
F545
F513
F561
F5FA
F634
F5B5
F536
F63D
F9C2
FEF6
0385
055E
048A
0330
03B6
06AD
0A8B
0D50
0E42
0E1D
0DE0
0DCB
0D8E
0D17
0CD5
0D25
0DD1
0E45
0E2B
0DAF
0D2C
0CE7
0CFB
0D61
0DD4
0DD5
0D26
0C40
0C19
0D0E
0E0B
0D39
09E9
05AF
0315
0324
046F
04D7
03DE
02CE
02C1
0339
0328
02AB
02C9
03A4
0408
0344
027F
0333
04A2
0415
0003
FA2C
F5CF
F437
F416
F413
F49F
F6AE
F993
FB60
FB3B
FA46
FA06
FAA9
FB54
FB94
FBBD
FC0C
FC22
FBAF
FB15
FAEE
FB35
FB64
FB48
FB40
FB95
FC0C
FC22
FBAE
FB13
FAE2
FB3F
FB8B
FAE0
F902
F6CE
F592
F5BF
F680
F6B4
F630
F5B7
F5CA
F616
F627
F60E
F601
F5E3
F59E
F59A
F62C
F6C8
F68C
F5EA
F6F5
FB31
013C
059F
0644
0490
03AB
0546
088E
0BB0
0D88
0DFD
0D94
0D0E
0D0B
0D91
0E0C
0E04
0DBC
0DC1
0E0A
0DFB
0D5F
0CCA
0CC0
0CEF
0CC9
0C73
0C82
0CFB
0D41
0D0D
0CEB
0D55
0DA8
0C8E
0991
05F0
0386
0314
03C1
042F
03C4
02FB
02AE
0319
0398
038E
033A
0355
03D2
03D0
0302
0282
035D
0480
0333
FE3C
F7D9
F3C2
F355
F4B2
F5AF
F652
F7C4
F9E1
FB2E
FB01
FA68
FA95
FB4C
FB82
FB01
FA9D
FAD4
FB28
FB0F
FAE0
FB2E
FBC1
FBDE
FB5D
FAD7
FAC7
FB06
FB36
FB45
FB60
FB8B
FB86
FB07
F9F3
F875
F6FB
F610
F5F5
F650
F684
F665
F648
F654
F649
F602
F5CF
F5DF
F5E2
F5A0
F58F
F625
F6CE
F682
F5AE
F6B4
FB68
023C
0712
0766
04F5
03AB
057E
0913
0C01
0D4F
0D96
0D9E
0D94
0D66
0D2E
0D23
0D57
0DBC
0E31
0E70
0E32
0D9A
0D28
0D1B
0D25
0D01
0CEE
0D35
0D72
0CFF
0C11
0BC4
0CAB
0D9A
0C92
0905
04BF
023D
023E
035E
03E8
038E
032C
0352
0389
0322
0255
0222
02E8
03AE
035E
0269
026B
03D3
04A5
025B
FCEC
F731
F408
F39D
F41E
F477
F567
F7B1
FA68
FBD5
FB90
FAD4
FAC8
FB3D
FB52
FACC
FA45
FA49
FAB3
FB09
FB21
FB28
FB41
FB58
FB51
FB29
FAEA
FAAC
FA80
FA64
FA59
FA86
FAF7
FB34
FA78
F89F
F690
F56B
F561
F5A9
F59A
F557
F54F
F570
F561
F541
F581
F5FC
F5F7
F554
F4F8
F57C
F613
F5C0
F555
F733
FC6D
02E2
06E9
06F2
04E9
03FC
05A3
08F2
0C21
0E01
0E60
0DD2
0D36
0D17
0D53
0D7D
0D7F
0D98
0DD0
0DD9
0D87
0D25
0D11
0D28
0D08
0CC2
0CD6
0D51
0D7B
0CDF
0C23
0C46
0D21
0D3A
0B4A
07AA
042B
027C
02C2
03AB
03DA
032D
02A2
02FD
03D4
0420
03A4
0340
0392
03DD
0327
0218
0279
045C
0501
01BC
FB75
F608
F422
F4BA
F52E
F4C9
F515
F70E
F987
FAD0
FADF
FADF
FB59
FBCC
FBCE
FB9A
FB75
FB46
FAFB
FAE0
FB2F
FB95
FB8F
FB1F
FAC7
FAD0
FB00
FB12
FB0C
FAF1
FAB6
FAA3
FB2B
FBE2
FB69
F90E
F616
F490
F4F8
F5C5
F579
F469
F400
F4AC
F576
F57B
F4EC
F461
F418
F44B
F54A
F69C
F6D9
F580
F48D
F6EA
FCF2
0365
0673
0587
037C
0369
05F7
09BA
0CFE
0EB6
0EA4
0D8A
0CD1
0D3B
0E02
0DE5
0CDF
0C18
0C43
0CC2
0CB3
0C3E
0C36
0CBA
0CFA
0C7E
0BDA
0BC1
0C04
0C1B
0C2A
0CAF
0D51
0CD8
0A79
06E2
03C0
0256
0290
0345
035D
02C4
024A
02A4
0390
0425
03FF
03C0
0404
0445
03A3
02A3
02DE
0464
04B1
0156
FB40
F60F
F417
F438
F422
F3B6
F4CD
F805
FB5F
FC90
FBAB
FA89
FA53
FAB2
FB0A
FB49
FB79
FB57
FAD7
FA7F
FACF
FB84
FBE3
FBB2
FB6E
FB7D
FBAE
FBAD
FB8E
FB7D
FB6A
FB47
FB3A
FB10
FA0C
F7D8
F563
F427
F481
F551
F569
F4EE
F4D6
F572
F609
F5F6
F569
F4ED
F4C0
F4FA
F5A5
F644
F5ED
F4B6
F48B
F796
FD89
034F
05E0
0528
03C5
0437
06D2
0A3E
0CFF
0E40
0DED
0CD8
0C56
0CFC
0DF3
0DFC
0D12
0C5F
0CAB
0D60
0D6E
0CA4
0BBC
0B4E
0B40
0B58
0BB0
0C3E
0C7F
0C16
0B85
0B9F
0C45
0C34
0A47
06C5
0355
01A4
0200
0334
03CF
037D
030A
0325
0371
0324
024F
01FF
02C4
03B5
03AC
0318
0372
04A7
044D
005C
FA20
F533
F3A8
F43B
F49F
F487
F574
F808
FACD
FC0A
FBC2
FB39
FB22
FB29
FAF4
FAB4
FAA0
FAA0
FAA0
FAD1
FB4E
FBB8
FB96
FB05
FAA9
FAF0
FB8F
FBFA
FC00
FBD7
FBBA
FBBD
FBB7
FB2D
F9A3
F751
F540
F45E
F486
F4D2
F4B6
F48A
F4DA
F59D
F644
F66A
F61C
F599
F535
F557
F611
F692
F5D4
F452
F45C
F7E7
FE0D
036D
0558
0449
0310
03F7
06F8
0A71
0CDF
0DC6
0D99
0D34
0D3D
0D94
0D81
0CAF
0BC2
0B9B
0C38
0CC6
0CB5
0C54
0C3C
0C6E
0C71
0C18
0BBD
0BAB
0BB4
0B9E
0BA5
0C1A
0C9D
0C20
09EB
067D
035E
01F5
0264
037A
03DF
0359
02C2
02CE
033C
0361
033B
0352
03A6
036F
0261
01AD
02A8
0473
0421
FFF9
F9D1
F553
F422
F4B1
F4DD
F4A9
F5A9
F858
FB24
FC4A
FBC3
FAE1
FA8D
FAA8
FACD
FAF3
FB20
FB27
FAE4
FA8B
FA72
FAA0
FAD1
FADB
FAE9
FB32
FB9D
FBCD
FB93
FB2B
FAFE
FB2C
FB4B
FAA8
F8FD
F6E2
F556
F4C3
F4BB
F4BD
F4D0
F530
F5A4
F5AC
F543
F4FE
F549
F5DE
F63E
F667
F68F
F668
F571
F44A
F4F5
F8E6
FEF2
03E8
0572
0431
02EC
03F8
0766
0B69
0E0B
0E91
0DAD
0CAE
0C60
0C92
0C99
0C4F
0C2F
0C89
0CEB
0CC6
0C3E
0BFF
0C4A
0CA0
0C7B
0C08
0BDE
0C2B
0C85
0C94
0C85
0C94
0C5D
0B0F
0856
04F4
024A
0151
01E0
02E8
0370
0367
0361
03AA
03EC
03C6
036C
033D
030A
0253
0160
0172
031D
04BE
038C
FEAA
F881
F46E
F383
F422
F48F
F4F0
F662
F8E3
FAFA
FB79
FACB
FA3D
FA6B
FAE9
FB2A
FB29
FB1E
FB0C
FAD4
FA92
FA92
FAF1
FB62
FB76
FB1E
FAC1
FAC3
FB14
FB47
FB2A
FAFD
FB11
FB2B
FA9D
F910
F70D
F587
F4F2
F500
F545
F59D
F5D9
F597
F4C1
F3FF
F41D
F503
F5BF
F5C0
F590
F5F2
F695
F67A
F5AB
F5E8
F8DC
FDFF
02CA
0515
04FE
0474
054F
07E5
0B17
0D5E
0DE5
0D0D
0C0E
0BF2
0CB5
0D7B
0D98
0D36
0CDC
0CB1
0C83
0C4F
0C56
0CA7
0CEE
0CE1
0CAE
0CAE
0CE1
0CE9
0CA5
0C6C
0C82
0C6A
0B38
088E
0539
02AD
01E8
02AE
03D5
0443
03CA
0310
02C7
030E
0383
03BC
038E
0300
0251
0208
029C
03B2
03DC
01A4
FD1E
F821
F4A7
F334
F2F8
F348
F458
F66A
F8D9
FA70
FAAA
FA33
FA03
FA51
FA98
FA80
FA4C
FA68
FAD6
FB35
FB44
FB24
FB18
FB26
FB0F
FAAF
FA46
FA36
FA94
FB14
FB6C
FB92
FB84
FB00
F9B0
F7BC
F5EB
F504
F50B
F55D
F57A
F56F
F569
F54B
F4E6
F462
F41D
F435
F480
F4FA
F5C7
F695
F67B
F513
F3AF
F4B4
F92A
FF3B
039F
04A7
03A6
0356
053D
08A6
0BC0
0D51
0D60
0CC7
0C6C
0CA8
0D25
0D3C
0CB2
0C0E
0C09
0CAF
0D3E
0D02
0C24
0B77
0B90
0C3F
0CEE
0D43
0D46
0D13
0CC4
0C9B
0CF4
0DAC
0DD8
0C6E
0962
05F0
0398
02DA
0306
032A
02F8
02C5
02EA
0358
03BE
03D3
0383
0302
02B7
02F0
0388
03FD
03FD
03A0
02F6
0182
FE95
FA52
F604
F331
F25D
F2EA
F41A
F5BB
F7CA
F9CD
FAFD
FB0A
FA67
F9D3
F9BE
FA1F
FAA8
FB0B
FB2C
FB2A
FB36
FB4A
FB24
FAAA
FA41
FA67
FB04
FB66
FB24
FA96
FA58
FA82
FABF
FAE2
FAFA
FAC7
F9B8
F7B9
F5B9
F4E0
F542
F5D4
F5B6
F51E
F4B1
F48A
F463
F452
F4BD
F584
F5DD
F550
F47A
F44F
F4CA
F4F9
F483
F4A1
F707
FBDE
0136
0498
0505
03A9
02C7
0405
0743
0AE7
0D30
0D8D
0CCC
0C34
0C60
0CED
0D18
0CA1
0BFF
0BD7
0C4F
0CE9
0D0D
0CA7
0C3C
0C3C
0C76
0C77
0C53
0C96
0D4C
0DB0
0D2B
0C57
0C50
0D08
0CE2
0A81
06A0
0385
029A
0328
038D
0328
0295
0288
0302
0389
03B8
037F
0322
0300
0330
0351
0308
02A3
02CF
034E
0270
FEC1
F92B
F49A
F302
F382
F407
F40C
F4D7
F732
FA08
FBA6
FBA5
FB00
FA9C
FA81
FA84
FAC6
FB3C
FB60
FAE8
FA5E
FA69
FAE3
FB2B
FB1B
FB09
FAFE
FA8F
F9B3
F927
F98E
FA91
FB55
FBA2
FBCF
FB9E
FA2D
F77F
F526
F49C
F562
F5C0
F50C
F457
F4A9
F585
F5AA
F4D6
F3EB
F396
F3A6
F3E4
F4A6
F5E6
F690
F5AA
F40F
F422
F779
FD3A
02CC
05E8
0609
0469
030D
038C
062E
09BC
0C6E
0D50
0CD9
0C25
0BE3
0C15
0C79
0CD1
0D00
0D0E
0D08
0CCB
0C2E
0B87
0B91
0C88
0D9C
0DCC
0D2C
0CC8
0D10
0D11
0BE7
0A7B
0AAC
0C84
0D7E
0B58
06E4
0325
01FA
0296
032B
0318
0303
036F
0406
042B
03B0
02DE
022D
021B
02BD
0367
036A
0332
03B1
0452
02B5
FD82
F6F0
F308
F34E
F542
F5C0
F4CF
F4E8
F723
F9BE
FACA
FAA4
FAC7
FB5D
FB6A
FABF
FA57
FAB9
FB33
FB10
FAB3
FAD0
FB27
FAE3
FA06
F98A
F9EA
FA7C
FAA1
FAA9
FAE5
FADC
FA35
F9C8
FA88
FBAF
FB4B
F8C5
F5EE
F4CE
F534
F550
F458
F366
F384
F431
F483
F4AF
F551
F5F9
F5AA
F49D
F433
F4FB
F5BA
F526
F402
F4A8
F85F
FDDF
0293
04D3
04AC
0346
0244
0319
060B
09CA
0C87
0D7C
0D37
0CAE
0C63
0C5F
0C76
0C74
0C3C
0BF9
0C01
0C5E
0C9D
0C75
0C5E
0CE7
0D9F
0D78
0C7C
0C02
0CB6
0D5B
0C84
0AE3
0A91
0C0A
0D04
0B1C
06DF
0341
0235
02EE
039A
03A5
039F
03C4
03CB
039E
037C
0377
036A
0351
0329
02BE
021F
0211
0328
042F
0280
FD11
F6A4
F365
F437
F5EB
F5AE
F49D
F598
F8D9
FB94
FBD2
FAB6
FA55
FACA
FAB1
F9C8
F961
FA23
FAE9
FA9B
F9DE
F9DF
FA75
FAA3
FA58
FA64
FAEA
FB1F
FAB1
FA5A
FA9D
FAD3
FA45
F9A5
FA26
FB41
FAD5
F805
F4C3
F37B
F439
F533
F560
F53F
F549
F52D
F4D2
F4F5
F5F8
F6CC
F62B
F4A0
F40A
F4ED
F597
F4C0
F3D6
F570
F9FB
FF33
02B4
0404
040D
03B8
03A1
046E
067E
0934
0B52
0C40
0C91
0CF2
0D46
0D28
0CB6
0C4F
0C00
0BBF
0BD6
0C78
0D34
0D6B
0D2E
0D0A
0D0B
0C9F
0BB2
0B3E
0C07
0D28
0D07
0BA8
0AEE
0BE0
0CE2
0B9E
0813
0494
0300
02FD
0323
02E6
02BD
02F0
0315
02D5
027D
027E
02CD
0317
0325
02EF
02B6
031C
0441
049D
01E8
FBFE
F619
F3D4
F52D
F6B0
F5E1
F43E
F4DA
F7F6
FAAB
FAE9
F9E7
F9C0
FA70
FA88
F9E3
F9C8
FAA3
FB3E
FAB2
F9DB
FA06
FAF0
FB3D
FA93
FA05
FA3C
FA81
FA2F
F9E5
FA53
FAD5
FA6E
F98A
F96D
FA0D
F9D3
F7D2
F546
F418
F484
F52A
F533
F51E
F563
F58E
F558
F569
F625
F696
F5D1
F4AD
F4B4
F5A5
F583
F3AD
F29D
F53E
FB19
008C
02F4
0324
0350
03FD
0462
04B3
063F
0954
0C60
0DC4
0D95
0D1B
0D13
0D35
0D24
0CFD
0CD6
0C76
0BE8
0BBE
0C3D
0CD0
0CDB
0C94
0C81
0C84
0C2E
0BC1
0C05
0D07
0DC5
0D7F
0CC7
0C89
0C5C
0AC4
076A
0406
027F
02BE
032A
02DB
0265
028C
0319
0347
02E5
0293
02D7
036B
0397
0329
02D3
0356
0448
03CF
002E
F9FD
F476
F29F
F412
F586
F4DE
F397
F475
F7A9
FA90
FB20
FA2F
F9CD
FA70
FAE9
FAA1
FA72
FAEB
FB41
FAB0
F9E0
F9EF
FAB3
FB20
FB00
FB21
FBC2
FBEF
FAF7
F9AB
F958
F9F5
FA57
FA26
FA42
FAF2
FAE8
F910
F660
F4BD
F4A1
F4E9
F4BB
F480
F4C2
F531
F557
F57A
F5FA
F62F
F536
F3B9
F368
F463
F4B8
F388
F341
F6F3
FDF9
0417
0632
0558
047C
0484
0441
03A0
0494
0817
0C14
0DB4
0CDA
0BCE
0C05
0CBB
0CCA
0C6D
0C7B
0CDF
0CD4
0C46
0BF9
0C42
0C82
0C41
0BF5
0C1E
0C53
0BFB
0B69
0B62
0BE0
0C32
0C30
0C5A
0C8F
0B88
086B
0476
021D
0257
03A2
0413
0387
0322
034B
0343
028F
01D3
01E1
029A
0330
0352
038B
0435
0468
0272
FDAF
F7B1
F352
F24F
F3B8
F4F1
F476
F36C
F411
F6D4
F9B8
FAC4
FA2E
F999
F9D9
FA54
FA64
FA4E
FA9A
FB0E
FB10
FAAE
FA8F
FADD
FB13
FB01
FB2C
FBD0
FC40
FBE8
FB40
FB08
FB0C
FA8F
F9C6
F9DC
FB0E
FBB3
FA10
F6C3
F448
F40A
F505
F598
F594
F5AE
F5FE
F608
F5DD
F5FE
F647
F602
F531
F4CE
F53D
F572
F4B5
F4A9
F7D6
FE01
038C
0579
04AA
0410
04AD
0525
04DD
056C
082C
0BC4
0DA0
0D3C
0C7F
0CC1
0D20
0C6E
0B5B
0B54
0C32
0C85
0BE6
0B87
0C3A
0D1D
0CE4
0BB9
0AEF
0B2A
0BBB
0BDB
0BA8
0B80
0B59
0B3B
0B8E
0C1A
0B71
0882
047B
0206
025A
03F3
0496
03F1
0364
03A5
03D5
0326
023A
0213
0268
0224
0140
00F9
01EA
02BB
0155
FD2B
F7F6
F42A
F2F3
F397
F486
F4C3
F48C
F4E3
F66C
F8A5
FA55
FACE
FA85
FA48
FA47
FA1F
F9A0
F911
F8D5
F914
F9BC
FA92
FB3F
FB7C
FB60
FB5D
FBBB
FC32
FC46
FBF0
FB8D
FB34
FAA4
FA06
F9FF
FAA4
FAEA
F9C2
F793
F5DB
F56B
F593
F55A
F4DD
F4EE
F596
F5F4
F59E
F54A
F5B6
F684
F6DA
F688
F5FE
F582
F54C
F631
F931
FDFA
0279
04A8
048F
03DB
03C3
0434
050A
06DC
09C3
0C59
0D0A
0C23
0B81
0C3A
0D6A
0DB2
0D0D
0C73
0C44
0BFE
0B89
0BA2
0C8D
0D44
0CC7
0B9B
0B24
0BBA
0C4E
0BF5
0B0B
0A94
0B06
0C18
0D32
0D7A
0BDD
080A
03A4
0156
0221
0425
04CE
03B6
0282
0257
029B
0267
020D
025A
0302
02F7
024A
0266
03CA
047A
01E1
FC0F
F619
F31D
F377
F516
F5D8
F52F
F3E2
F31A
F3B6
F5D3
F87C
FA30
FA33
F953
F8F6
F98E
FA59
FA96
FA70
FA84
FADD
FAE4
FA44
F97D
F950
F9E2
FAA2
FAFE
FAF7
FAF2
FB2F
FB93
FBCA
FB9A
FB14
FA8D
FA5A
FA8E
FAD3
FA91
F958
F74C
F543
F435
F47A
F57B
F639
F630
F5AD
F556
F56F
F5BE
F607
F649
F67B
F64C
F592
F4F0
F5B6
F8C4
FD7A
01EE
0461
0493
03B3
0316
030E
031A
0304
0384
0590
0907
0C63
0E09
0DC8
0CE2
0C93
0CEE
0D47
0D47
0D2F
0D2A
0CE7
0C2D
0B67
0B34
0B8F
0BCD
0B98
0B61
0BAA
0C47
0CB2
0CC3
0CBA
0CA3
0C50
0BF9
0C41
0D0F
0CEC
0A62
060F
027E
0189
0276
0339
02F6
0282
02A2
02E3
029F
023E
0299
036E
03A1
030C
02E2
03A8
03AE
00C0
FB1A
F5AE
F32E
F394
F4D6
F55A
F4F2
F40A
F310
F2D8
F470
F7B6
FAC2
FBA1
FA7B
F942
F952
FA28
FA97
FA79
FA80
FAE2
FB0D
FAB7
FA65
FA8B
FAC3
FA80
FA07
FA0D
FA9D
FB0B
FAFB
FAD0
FAF2
FB29
FB15
FAF0
FB2F
FB8A
FAF9
F904
F686
F4D3
F469
F4D3
F574
F5E7
F5E7
F571
F4FD
F522
F5D3
F65E
F653
F617
F61A
F5FF
F563
F546
F7A6
FCDF
025B
04DA
03EE
0246
0262
03E2
04A3
03E4
035C
04FA
087C
0BC7
0D49
0D53
0D26
0D59
0D83
0D1A
0C46
0BB9
0BDE
0C66
0CB0
0C84
0C26
0BDA
0B9F
0B7B
0BB0
0C59
0D1B
0D68
0D2D
0CD9
0CA8
0C4C
0BAD
0B82
0C56
0D0F
0B98
0783
0330
0174
0284
0400
03F6
02DB
023B
026E
0294
024E
0242
02C1
032B
0335
039E
04A4
0496
0153
FB31
F54C
F27A
F2B5
F3F8
F4DB
F562
F59F
F51D
F412
F3F5
F5D7
F8C3
FAB2
FAE3
FA5D
FA49
FAB5
FB12
FB27
FB0D
FAB0
FA0D
F9B2
FA35
FB27
FB55
FA6B
F98A
F9C3
FAA4
FB13
FAF3
FB10
FB99
FBC1
FB13
FA5F
FA9D
FB68
FB55
F9CB
F7A7
F607
F529
F4E8
F556
F63C
F6A1
F5D0
F480
F429
F520
F63F
F689
F659
F660
F646
F566
F4C4
F6B7
FBEA
01B6
04A2
0417
02A7
02B8
0409
04C4
0429
036B
041C
0674
094D
0B63
0C43
0C4C
0C29
0C46
0C83
0C94
0C96
0CE9
0D66
0D48
0C37
0B01
0AB9
0B6C
0C2B
0C5A
0C49
0C79
0CC6
0CCC
0CAF
0CC0
0CAA
0BE2
0AF0
0B20
0C53
0C50
0960
04E2
0211
0246
0394
038F
0248
01A0
024F
0321
0313
02BD
02F6
0357
032E
02EE
0348
034C
00F4
FBF3
F6C1
F41D
F428
F4D2
F4C1
F48D
F4FC
F582
F54B
F4E1
F595
F792
F9A1
FAB6
FAF4
FB08
FB39
FB60
FB54
FAFB
FA33
F92C
F8B1
F96E
FAE5
FBC1
FB73
FAD2
FABF
FAEE
FAB1
FA50
FAA6
FB9E
FC08
FB24
F9C1
F949
FA0D
FAFF
FB02
F9DD
F805
F61E
F4E5
F4E9
F5CA
F662
F619
F5A4
F5DC
F673
F685
F60F
F5ED
F64C
F639
F54C
F516
F7B4
FCFF
0232
04CB
04E5
0443
03EF
03B3
0343
02D6
02C4
035B
0512
0828
0BB5
0DED
0DDB
0C84
0BB2
0BD6
0BFF
0BCA
0C07
0D0C
0DB1
0CE8
0B89
0B37
0C16
0CB9
0C58
0BCD
0BFF
0C68
0C12
0B63
0B8E
0C6F
0C98
0BC6
0B9E
0CE8
0D8B
0AFB
05FB
0220
018D
02B4
02F2
020A
01B8
029E
036A
0320
028E
02A7
02E4
0282
0242
0322
03E4
01BC
FC02
F5C8
F2C9
F36F
F4F8
F530
F49F
F4BE
F584
F5D6
F59E
F608
F7AF
F9AC
FAB6
FA95
FA09
F9CC
F9FE
FA69
FADA
FB27
FB21
FAC0
FA42
F9FE
FA12
FA65
FACB
FB07
FAEF
FAA5
FA85
FA9F
FA9A
FA3A
F9CC
F9D1
FA6B
FB42
FBC6
FB5F
F9B1
F71D
F4EB
F462
F55F
F643
F5C6
F49C
F47B
F5B1
F6B0
F65C
F59B
F5D2
F695
F640
F4C6
F484
F79F
FD34
0214
041C
03F1
037D
03BA
0468
04F7
04F4
0427
032D
0398
0671
0A9D
0D8C
0DDF
0CC0
0C3C
0CCC
0D47
0CF4
0C7C
0C95
0CD2
0C8A
0C18
0C4B
0CFD
0D3B
0CC5
0C71
0CCC
0D2E
0CC2
0BF4
0BDC
0C7C
0CAC
0BFF
0B95
0C3E
0CBD
0B10
0728
034B
0180
019A
0227
027F
02FA
039F
03C7
034A
02F4
033E
0376
02FB
028D
032A
03D9
01FF
FC93
F621
F281
F2E4
F4FE
F61C
F5DB
F56F
F549
F4D8
F420
F448
F613
F89E
FA4C
FA9B
FA69
FA91
FAEE
FAED
FA8E
FA57
FA81
FAC0
FAD1
FAC8
FAC2
FAA1
FA38
F99C
F927
F92F
F9C1
FA96
FB3D
FB69
FB11
FA7B
FA1A
FA48
FAEB
FB60
FAD3
F8F4
F688
F500
F529
F641
F6CE
F64B
F591
F577
F5B7
F59B
F53B
F541
F596
F540
F41F
F410
F734
FD1B
029D
04F9
0467
0333
02FD
039A
0421
041B
039E
0323
038D
05B4
093D
0C54
0D48
0C74
0BCE
0C6B
0D5D
0D5C
0CAC
0C78
0CEF
0D17
0C6D
0BB9
0BE1
0C9C
0CEA
0C85
0C1D
0C3F
0CA8
0CF0
0D17
0D15
0C8F
0B8F
0AFD
0B89
0C57
0B99
08AC
04FE
029A
0225
02AB
0303
02D4
0258
01E3
01DA
028D
039E
0424
03D2
0381
03D2
03B5
0141
FC32
F6CF
F3C6
F383
F440
F477
F458
F4AF
F546
F53F
F4A2
F497
F5F3
F825
F9EA
FAA0
FAA4
FA8B
FA79
FA4F
FA25
FA40
FAA3
FAF4
FAEF
FABB
FAB0
FAEB
FB28
FB1A
FAD4
FABE
FB0D
FB6C
FB62
FAFA
FAB6
FAD6
FB11
FB1E
FB2D
FB6A
FB4C
F9F5
F779
F53B
F484
F507
F567
F515
F4E1
F578
F63E
F645
F5C2
F5A3
F5E3
F572
F436
F432
F782
FD7A
02D6
0513
04BB
03F7
03DC
03F8
03DC
03D2
03F7
03DC
039C
0482
0780
0B60
0DA4
0D70
0C85
0CCF
0DF6
0E39
0D1D
0BF5
0BDA
0C45
0C3B
0BE9
0C32
0CFE
0D28
0C42
0B5A
0B81
0C3F
0C5F
0BB4
0B2A
0B50
0BB9
0BF6
0C4C
0CD7
0CA0
0A6B
068D
0315
01D3
028F
03A0
03CA
031B
024F
0202
0257
02F4
0348
032D
0314
0334
029F
FFDD
FAD9
F5C1
F32B
F36E
F48F
F4DA
F4B0
F527
F5F0
F5BC
F46E
F3AF
F4F4
F7A5
F9D3
FA74
FA2C
FA10
FA58
FA9E
FABA
FAD7
FAEB
FAC7
FA92
FAA6
FB02
FB31
FADB
FA3F
F9EB
FA2B
FAC9
FB50
FB72
FB3C
FAE8
FAA4
FA85
FA9C
FAFC
FB8A
FBBA
FAC4
F884
F605
F49F
F47D
F498
F444
F407
F47A
F51F
F510
F48D
F4C3
F5F0
F6BF
F645
F5F5
F844
FD5C
0271
04DE
04D0
043A
0420
0422
0406
0439
04AA
0476
0379
034F
0599
0993
0C95
0D2A
0C87
0C75
0CED
0CD0
0C15
0BDE
0CA0
0D6D
0D50
0C92
0C1B
0C2B
0C55
0C6E
0CAF
0CF8
0CB4
0BE4
0B80
0C35
0D53
0D9E
0CE3
0C0B
0BE3
0C4A
0C76
0B8E
0933
05F8
035B
02A8
038D
043A
0377
023D
025F
03D5
04A1
03BE
02B2
0325
03DE
01CE
FC1B
F5B5
F247
F269
F3BE
F437
F408
F44B
F513
F5A3
F5BD
F5AF
F56A
F494
F396
F3B5
F5AD
F8A9
FAFA
FBB8
FB5E
FAF1
FAE8
FB10
FB1B
FAF9
FAB6
FA64
FA2C
FA3A
FA88
FAD8
FAF1
FAD5
FABD
FAE7
FB38
FB3B
FA9B
F9B7
F955
F9BA
FA4F
FA78
FA6A
FACE
FB82
FB50
F950
F653
F44D
F447
F55C
F5FA
F598
F4DD
F482
F499
F4CB
F4CC
F48E
F47A
F587
F8AC
FDA7
029D
056A
058F
047D
03DB
03EC
03E7
0371
031A
036F
0424
046B
03F5
0368
03DA
05D9
08E1
0BA5
0D04
0CEB
0C5E
0C6A
0D14
0D87
0D40
0CB4
0CA3
0D0A
0D3F
0CE0
0C45
0BEC
0BE2
0BF6
0C3A
0CC6
0D2F
0CCD
0BAF
0AE3
0B42
0C58
0CF8
0CD8
0CD6
0D60
0D4A
0B0E
0713
03BB
02D0
038B
03D9
030D
026F
02FD
03CA
0362
0226
01ED
0338
03D3
0136
FBB5
F66B
F3F9
F42A
F502
F53F
F528
F547
F572
F54B
F50C
F51F
F551
F511
F47B
F482
F5E2
F826
FA0C
FAC1
FA84
FA26
FA27
FA69
FA93
FA88
FA6F
FA6D
FA7B
FA6B
FA2B
F9ED
FA03
FA81
FB24
FB98
FBC4
FBB6
FB80
FB34
FAE5
FA9A
FA47
FA02
FA12
FAA9
FB6D
FB87
FA55
F818
F5DC
F4A2
F4A2
F547
F5B7
F56F
F4AE
F44D
F4DC
F5D2
F610
F583
F5D4
F8D3
FE28
0321
0531
045B
02DE
0298
0361
03F2
03C3
036C
039B
0433
0489
0431
0383
0385
052C
085F
0BB5
0D88
0D71
0CA5
0C85
0D21
0D75
0CFC
0C5B
0C56
0CB6
0CC4
0C6C
0C41
0C6F
0C71
0BFA
0B97
0BF4
0CC8
0D19
0C8E
0BEF
0BFC
0C60
0C56
0BFE
0C43
0D33
0D4A
0AFD
06CC
031E
01D9
028D
0359
0346
030A
036F
03DE
034D
021B
01DE
02F9
0351
006D
FAAC
F56B
F380
F45A
F538
F4B5
F3F2
F44D
F53B
F54B
F471
F407
F4A6
F53E
F4D2
F443
F55A
F844
FB0C
FBDA
FB04
FA44
FA74
FAE1
FAAD
FA07
F9BE
FA20
FAC0
FB1E
FB2D
FB23
FB19
FB06
FAED
FAE0
FAE0
FAE8
FB03
FB38
FB63
FB54
FB0B
FAC6
FACD
FB35
FBC3
FBDB
FAC8
F85E
F57C
F3A9
F3DD
F57A
F6C4
F68E
F565
F4D5
F57E
F64A
F5D8
F491
F4BB
F827
FDEE
02E7
049C
038B
0242
028E
03F2
04DB
04A0
03FB
03CC
0413
0421
0392
02D1
02E1
0493
07CE
0B4B
0D5D
0D5B
0C54
0C02
0CEF
0E07
0E26
0D7A
0D04
0D1E
0D38
0CE6
0C88
0C99
0CDB
0CC1
0C5F
0C45
0C73
0C44
0B95
0B45
0BF4
0CCE
0C84
0B54
0B07
0C72
0DCC
0C77
0843
03E9
0212
0296
034E
0307
027F
02A0
02FB
02AB
0211
0267
038E
035B
FFE6
FA2A
F571
F3EF
F4A8
F522
F474
F3D6
F457
F53C
F532
F45C
F42F
F53F
F646
F5E6
F4B9
F4C5
F6E5
F9B1
FB3D
FB38
FAC5
FABE
FAE2
FAB3
FA4F
FA13
F9F9
F9C9
F9BD
FA45
FB37
FBBD
FB61
FAB8
FA9D
FB1D
FB8A
FB7F
FB44
FB32
FB2F
FAE8
FA5D
F9E5
F9CC
FA1D
FA9D
FAAF
F98E
F726
F4C3
F42C
F5A1
F73E
F714
F57F
F49E
F574
F680
F5E6
F465
F4F6
F941
FF5D
03B3
04A6
03B3
0324
03B3
0488
04DE
04C3
048E
0448
03DB
0369
031C
02F7
032E
046B
072B
0AC2
0D8D
0E6A
0DCA
0D06
0CCC
0CB4
0C47
0BE0
0C25
0CF8
0D7E
0D32
0C7E
0C14
0C13
0C2C
0C47
0C8A
0CC4
0C70
0B97
0B2B
0BF0
0D3C
0D94
0C91
0B8E
0BD2
0C9B
0BC8
0894
04C2
02A6
0293
02F2
029E
0218
0248
02ED
0328
0309
036D
041B
0323
FEFF
F8EB
F420
F299
F357
F413
F3F8
F3F9
F4D5
F5DC
F5FB
F553
F4F8
F560
F5CB
F571
F4B5
F4C5
F630
F846
F9D8
FA5B
FA2E
F9FD
FA1F
FA81
FAE0
FB04
FAE0
FA97
FA6B
FA89
FAE0
FB29
FB25
FAE8
FAD9
FB40
FBDA
FBFF
FB61
FA7E
FA24
FA8B
FB22
FB55
FB57
FBBF
FC70
FC4C
FA63
F74D
F4DC
F45A
F53B
F5D2
F53B
F44C
F473
F5C5
F6BB
F625
F506
F5EF
FA2A
0000
042C
0506
03DE
031B
03A0
046C
0471
03E2
0382
0381
0384
036B
0366
037C
03A5
0463
068D
0A04
0D23
0E3A
0D7C
0CAC
0CE2
0D58
0CF1
0C08
0BDC
0CA4
0D2E
0CA5
0BC5
0BC1
0C86
0CFA
0CA4
0C45
0C7A
0CBC
0C4E
0B92
0B82
0C17
0C33
0B62
0AC6
0B95
0D14
0D0A
0A4F
0642
034E
0272
02D1
0348
0392
03BD
0379
02A2
0202
0285
037F
02A8
FE94
F8CF
F4B0
F3E8
F4EC
F52B
F423
F35E
F3D5
F48D
F454
F3AF
F40A
F55D
F5E8
F4B5
F34F
F40E
F71B
FA2D
FB46
FABD
FA29
FA31
FA55
FA4D
FA88
FB2C
FB94
FB33
FA90
FA9E
FB64
FBE3
FB71
FA94
FA3B
FA94
FB18
FB5D
FB6D
FB71
FB74
FB80
FB8F
FB74
FB1D
FAD8
FAF8
FB0D
FA0A
F792
F4F4
F3FE
F4DC
F5D4
F584
F4A0
F4C4
F5F6
F671
F535
F3D7
F50E
F99C
FF5E
0374
04E0
04BC
0473
0474
0477
0456
042F
041E
0423
043F
0466
0451
03C1
0315
036C
05B6
0971
0CBD
0DF9
0D52
0C5F
0C4E
0CD1
0CF3
0C8A
0C4D
0CAE
0D2D
0D17
0C8E
0C3E
0C52
0C4A
0BF0
0BCB
0C48
0CF2
0D0C
0CA3
0C65
0C7D
0C45
0B75
0AEA
0B8E
0CB3
0C74
09EE
066A
03DE
02DB
0299
0281
02C2
0351
036B
02C3
0269
0379
04EE
03E6
FEDE
F806
F372
F2FE
F4C2
F5B4
F4FA
F404
F406
F473
F43E
F3A9
F3E2
F51B
F602
F578
F444
F44A
F644
F8E7
FA72
FA8C
FA45
FA8D
FB42
FBB6
FB9A
FB31
FAD8
FAC0
FAF1
FB4C
FB7E
FB3F
FAC0
FA97
FB0C
FBB5
FBF1
FB9D
FB1C
FAD1
FAD2
FB00
FB2E
FB27
FADB
FA91
FAAA
FAEB
FA67
F886
F617
F4B1
F4DB
F56C
F52D
F482
F4AF
F5B9
F616
F4EC
F3E2
F5AC
FAC9
0083
03A6
03A4
029C
0290
0377
0427
0436
0452
04FA
05AB
0598
04B3
03AC
030D
02EA
0380
0565
08A6
0BF5
0D9B
0D47
0C6A
0C7C
0D55
0DBB
0D37
0C90
0C7D
0C8C
0C07
0B4D
0B72
0C86
0D4F
0CF9
0C31
0BF2
0C11
0BBB
0B10
0B10
0BE5
0C59
0BA2
0AE5
0BC2
0DAC
0E04
0B4E
0719
040D
02E6
027C
0205
01F2
0284
02E7
0280
0230
030F
042D
02E4
FE04
F7CB
F3C7
F337
F451
F4D3
F452
F3DB
F41E
F4B4
F4EC
F4B8
F4A1
F502
F592
F5BE
F55B
F4FC
F587
F75E
F9C7
FB6A
FB8E
FACD
FA5D
FAD2
FBB1
FC2E
FBFD
FB6C
FAEC
FAB8
FAD6
FB45
FBEB
FC63
FC32
FB66
FABE
FAED
FBA8
FBEF
FB58
FAAB
FADC
FB9B
FB9B
FA6D
F95B
F9B7
FACD
FA92
F870
F628
F57C
F5F2
F5EC
F539
F52A
F61A
F672
F514
F3CE
F5D1
FBA0
01EC
0513
04CB
038F
0352
03E4
044A
0441
0420
041F
0438
046E
04A0
0467
03A6
030C
0368
0464
04D1
047A
04E2
075A
0AF7
0D5A
0D68
0C59
0BF5
0C81
0CDF
0C54
0B6D
0B29
0BB7
0C70
0CBB
0C96
0C58
0C4E
0C8E
0CF0
0D2E
0D1B
0CC2
0C3D
0BC0
0BA9
0C2B
0CC4
0C8D
0B60
0A5A
0AA4
0BCD
0BE6
0996
05C3
02B9
01CB
0253
02F2
031D
032C
0371
03B4
0339
010A
FCC4
F788
F3B5
F2E7
F44A
F57D
F52E
F443
F435
F4FA
F546
F491
F3BD
F3A6
F404
F45A
F4E0
F5CB
F654
F5AB
F488
F4C1
F70B
FA00
FBB9
FBD8
FB6A
FB2E
FAFE
FABE
FADF
FB75
FBBE
FB47
FAC7
FB14
FBC4
FBBF
FAF1
FA69
FAC6
FB52
FB0F
FA1B
F971
F998
FA28
FAA5
FB08
FB48
FB27
FACE
FAE7
FB78
FB77
FA19
F80A
F68F
F5DE
F542
F4B0
F4FB
F61C
F65C
F487
F274
F3D7
F9EC
016F
05D4
05D2
03DF
02D9
0364
045C
04B5
0469
0413
043B
04DE
0575
057D
0510
04D3
04FF
04D3
03A8
0284
0379
070F
0B1F
0D18
0CBF
0BE5
0BDD
0C48
0C56
0C24
0C52
0CD1
0D02
0CC9
0CBE
0D18
0D35
0C9C
0BD0
0B97
0BE9
0C2F
0C35
0C3C
0C45
0C0E
0BA5
0B7F
0BBC
0BE7
0BB8
0BA2
0C11
0C3F
0AB0
072B
0395
0212
02B0
0387
0320
020E
01FB
035F
048A
0301
FE05
F7B0
F35B
F2B5
F47A
F5FF
F5DD
F4D3
F44B
F490
F4DE
F4B3
F45E
F439
F42D
F434
F4A3
F570
F5CA
F525
F460
F505
F761
FA01
FB4D
FB37
FADE
FAED
FB12
FAF4
FAE9
FB43
FB9C
FB63
FAC2
FA61
FA82
FAD4
FB09
FB19
FB10
FAEC
FACD
FAD7
FAE9
FAAC
FA20
F9D7
FA3F
FAF4
FB45
FB45
FB95
FC0E
FB8E
F99A
F75C
F63C
F615
F5BD
F503
F4F4
F5E7
F669
F539
F3BE
F51C
FA6E
00F4
04D5
04F7
0372
02C0
0381
04C1
0573
054C
04B9
0465
049A
04E4
0481
0374
02C4
033C
042B
042C
0356
039D
0664
0A68
0CFE
0D11
0C0E
0BD0
0C94
0D47
0D45
0CF3
0CD0
0CBC
0C62
0BED
0BC6
0BEC
0C01
0BDC
0BB2
0BC5
0C27
0CB1
0D08
0CD6
0C3D
0BDD
0C24
0C9E
0C77
0BAC
0B49
0BFF
0CC6
0BA5
0815
0400
01D0
01E3
027C
022A
017D
020F
0427
05C2
0448
FF24
F8A0
F3F9
F2AB
F395
F49B
F4C2
F48E
F4AD
F4E7
F49F
F3F0
F395
F3DD
F450
F49A
F50D
F5D7
F654
F5D5
F4E5
F4FA
F6BC
F92D
FAC7
FB16
FAD8
FAC4
FAD7
FAE1
FAFD
FB3B
FB5B
FB41
FB42
FB8D
FBB9
FB60
FAE5
FAEC
FB4D
FB33
FA6D
F9FA
FAB6
FBF6
FC39
FB24
F9FC
F9EF
FABD
FB81
FBF2
FC16
FB77
F9A5
F746
F5BD
F588
F5CA
F5B7
F5AC
F627
F65A
F528
F395
F4A4
F9D6
00AD
04FF
0552
03E1
037B
048A
058C
058A
04FD
04AD
0495
044D
03CF
036C
0342
0340
0356
0358
031A
030D
044B
075C
0B16
0D6A
0D76
0C5B
0BC0
0C05
0C51
0C1F
0BE2
0C14
0C5C
0C33
0BD8
0BF2
0C79
0CA5
0C0C
0B3E
0B16
0BAB
0C3F
0C23
0B7E
0B19
0B7A
0C4B
0CB2
0C3A
0B69
0B34
0BBE
0BC7
09DE
063B
02F6
01FA
0301
040A
03B3
02A5
028C
03E5
0512
03B3
FEF8
F89D
F3A8
F20A
F33A
F503
F5A8
F534
F4CA
F4FC
F54E
F52A
F4B5
F46B
F476
F4CA
F579
F665
F6DA
F62C
F4E0
F499
F658
F91A
FADE
FAEA
FA60
FA80
FB17
FB2D
FA9B
FA24
FA3D
FA82
FA87
FA81
FAE0
FB84
FBD4
FB87
FAF5
FA90
FA73
FA85
FABF
FB0D
FB3A
FB44
FB70
FBD4
FC14
FBE5
FB8F
FB75
FB4D
FA4B
F83D
F609
F4D2
F4D7
F57E
F639
F6C0
F69E
F577
F435
F50B
F961
FFCA
04E5
0678
054D
03E6
03D3
04A1
050C
0494
03C6
035F
0394
03FF
0412
03AF
035B
039C
0425
041E
0388
03CE
0647
0A53
0D99
0E6C
0D6E
0C7A
0C66
0C84
0C3C
0C0E
0C99
0D55
0D2F
0C28
0B77
0BEE
0CE5
0D23
0C73
0BC3
0BD9
0C6E
0CC4
0CA1
0C5D
0C2D
0BE9
0B76
0B12
0B0B
0B64
0BC2
0B8F
0A34
0786
0453
0227
0201
0320
039F
02A1
0172
01E6
0391
038F
FFA7
F93A
F43E
F337
F4EB
F653
F608
F504
F485
F46D
F410
F3A6
F3F8
F4F3
F5A0
F5A7
F5C5
F667
F6AA
F5A8
F443
F47C
F6EF
F9DE
FB37
FAE0
FA59
FA8A
FAE3
FAB7
FA58
FA5C
FA99
FA93
FA6E
FAA2
FB11
FB27
FADE
FAD6
FB3C
FB55
FA9F
F9E5
FA46
FB71
FBE3
FB13
FA4F
FAD2
FBFB
FC52
FBB8
FB58
FB9A
FB61
F9B6
F756
F5C2
F553
F534
F50B
F566
F63F
F674
F5AF
F5D4
F91A
FEEB
03EB
057F
045D
0328
0343
03DD
03D6
035D
034E
03C0
0412
03F3
03AE
0391
038F
037E
0342
02D8
0292
0343
0595
0914
0C2A
0D7B
0D36
0CA2
0C8A
0C91
0C39
0BDC
0C24
0CEF
0D62
0D0C
0C69
0C38
0C9F
0D29
0D58
0D10
0C8A
0C16
0BED
0C1F
0C82
0CD5
0CEA
0CAA
0C0F
0B54
0B10
0B93
0C12
0B03
07E6
044C
0275
02D8
03A8
030E
0171
00E7
026F
0458
03C2
FF81
F93C
F3F5
F1BD
F27B
F471
F5C2
F5CB
F53D
F505
F540
F55C
F502
F493
F4A1
F529
F5A2
F5B0
F573
F52E
F503
F535
F638
F81B
FA0E
FB03
FACA
FA41
FA52
FAF3
FB67
FB3E
FACA
FA93
FAAA
FABC
FAA3
FA92
FAC5
FB31
FB93
FBAE
FB70
FAF5
FA73
FA1C
FA06
FA2C
FA70
FAA4
FABC
FAF1
FB8D
FC63
FCA0
FB6F
F8EF
F661
F50E
F51D
F5B7
F62F
F68F
F6E5
F6C9
F62C
F650
F8FE
FE45
03A1
0621
0557
03A2
035A
0459
04C5
03C4
0285
0285
039A
0453
03F5
034E
0369
040A
0404
02E9
01D8
026C
0514
08BE
0BE1
0D9E
0E00
0D88
0CCB
0C38
0C00
0C09
0C25
0C4A
0C85
0CC0
0CB4
0C41
0BB2
0B83
0BE6
0C8B
0D03
0D23
0D10
0D06
0D27
0D67
0D7F
0D1D
0C4F
0BA7
0BBA
0C5A
0C80
0B29
0865
0564
0373
02E9
0311
02FE
0269
01EA
023F
0330
0339
00C9
FC09
F71F
F44C
F3D9
F43E
F429
F3CE
F3FC
F491
F4AC
F42D
F401
F4A8
F54E
F505
F452
F480
F5A6
F662
F5D6
F51F
F5F1
F842
FA3F
FAAE
FA4E
FA75
FB27
FB69
FAF8
FAA1
FAEF
FB60
FB41
FAC1
FA9B
FAEC
FB05
FA81
F9E4
F9F1
FAA7
FB53
FB5F
FAD4
FA38
FA2A
FAD3
FB8D
FB6E
FA82
FA03
FAE6
FC50
FC34
F9C1
F691
F4EB
F541
F630
F6A8
F6E0
F6EF
F600
F40A
F347
F663
FCF8
0339
05C5
0507
0406
0481
057A
057A
04BB
0452
0467
0461
044A
04B0
054F
050D
03AF
0288
02BE
0391
0360
0252
029D
05B2
0A19
0CF3
0D2A
0C20
0B99
0BF4
0C98
0D21
0D7C
0D62
0C8C
0B6B
0AF7
0B84
0C45
0C5F
0C09
0C11
0C9A
0CF0
0C94
0BEA
0B9F
0BC4
0BD6
0B8C
0B44
0B7F
0C26
0C92
0C47
0B8C
0B19
0B1E
0AC7
08EE
059C
028C
01A0
02BD
03CA
0331
01C2
017E
0294
02A3
FF67
F9AD
F4C8
F320
F3F7
F4DE
F496
F3DE
F3D8
F483
F502
F4D6
F461
F44C
F4C0
F552
F58C
F569
F542
F550
F561
F523
F4D4
F556
F72E
F98E
FAE3
FA9C
F9E2
FA1D
FB3A
FBE0
FB51
FA57
FA1E
FAAB
FB04
FAB4
FA5D
FAAC
FB6B
FBF0
FC03
FBCF
FB5B
FA9C
F9EC
F9DD
FA74
FB14
FB4A
FB4F
FB6A
FB45
FA85
F9CC
FA36
FB93
FC1A
FA78
F797
F591
F536
F588
F59B
F5C8
F681
F6F4
F61D
F505
F65B
FB3E
015D
0540
05E5
052A
04F7
0536
04E7
040E
03A1
0407
049E
04DC
0500
0549
0545
0492
03CC
03E1
04A1
04DC
0419
0386
04B6
07C1
0B26
0D54
0DEE
0D89
0CD1
0C43
0C45
0CDB
0D67
0D38
0C5A
0B87
0B46
0B58
0B3D
0AEC
0ACE
0B12
0B62
0B5D
0B24
0B27
0B89
0BEF
0BF9
0BBB
0BA3
0BFA
0C82
0CB4
0C66
0BFF
0BC0
0AFE
08B4
050D
01E9
0124
026D
037E
02D0
0181
01BC
0371
03CF
0075
FA80
F593
F40E
F50F
F61F
F605
F567
F531
F559
F54E
F4F8
F4B7
F4B7
F4B9
F47C
F40E
F3B7
F3BD
F437
F4D6
F51A
F4EE
F506
F648
F89F
FAC4
FB79
FAE5
FA56
FAA1
FB50
FB8A
FB56
FB68
FBF9
FC5F
FBEF
FAD7
F9E3
F99A
F9D9
FA2F
FA5E
FA6F
FA92
FAED
FB67
FB9C
FB48
FACA
FAD4
FB6C
FBB7
FB1E
FA51
FA81
FB9F
FC11
FAA1
F824
F67C
F645
F65B
F5DB
F56B
F5E6
F68A
F5DA
F442
F47D
F88C
FEE7
03CB
052D
0471
0410
04A1
0503
04A3
044A
04AE
0544
052A
047D
0411
041D
040D
03B8
03D3
04C0
0585
04F3
039D
03B5
0697
0AF9
0E1D
0E94
0D64
0C78
0C8F
0CF5
0CE0
0C72
0C5B
0CDB
0D75
0D71
0CA0
0B9A
0B30
0BA0
0C5C
0CA2
0C49
0BDA
0BDC
0C30
0C43
0BCF
0B3B
0B17
0B74
0BDB
0BDD
0B96
0B7A
0BB2
0B99
0A21
06FF
0371
015E
0165
0223
01DD
00BD
00AE
0299
046B
02DF
FD57
F6FC
F38D
F3AB
F4ED
F522
F47C
F454
F4F1
F55F
F51F
F4DF
F54B
F5DE
F59E
F492
F3D4
F42F
F523
F584
F4D2
F3BB
F381
F4E1
F777
FA10
FB90
FBC6
FB62
FB1E
FB0C
FADC
FAA5
FAE9
FBC6
FC8B
FC7B
FBAA
FAD1
FA5C
FA25
F9F1
F9E1
FA27
FA9A
FAE0
FAD4
FA8A
FA15
F99B
F99E
FA7F
FBB4
FC1F
FB83
FB02
FB93
FC5D
FB96
F8EE
F646
F570
F601
F636
F590
F535
F5B3
F5D6
F4C4
F428
F6BC
FCA0
029F
0586
056D
04C9
050A
055F
04CC
03ED
03F2
04BD
0533
04EA
0490
04A5
04D6
04DA
0512
05A8
05B1
0448
025D
025B
0568
09CC
0CBF
0D5F
0D0A
0D22
0D87
0D6E
0CD7
0C76
0C8B
0C9C
0C58
0C16
0C22
0C2F
0BE3
0B93
0BD3
0C7F
0CD7
0C8E
0C3B
0C6A
0CB8
0C54
0B42
0A87
0AE2
0BC9
0C11
0B70
0AD4
0B19
0BB5
0B0B
0832
0443
01A9
01C9
0380
0449
0315
017D
01AE
034F
034D
FF3D
F885
F353
F255
F431
F583
F4C5
F367
F368
F4DC
F635
F65F
F5BE
F53B
F4FB
F47F
F3A4
F2FE
F333
F440
F57E
F63F
F66E
F6A4
F796
F949
FAF2
FBB2
FB7D
FB10
FB1B
FB8D
FBDF
FBCB
FB8F
FB70
FB51
FAF4
FA66
F9FC
F9F9
FA5C
FAEC
FB5A
FB76
FB55
FB37
FB2C
FB02
FAA5
FA6A
FAB5
FB45
FB51
FAA6
FA31
FAD9
FBF0
FBB2
F986
F6F6
F5D3
F604
F610
F56C
F523
F5D5
F64F
F54B
F407
F58E
FAF5
0181
0579
05FF
052C
04E4
04F8
048D
03F8
0431
0517
057D
04F9
0488
04F0
0580
0532
045E
0435
04CF
04E5
03DA
0312
0481
0827
0BD6
0D85
0D3E
0C79
0C34
0C4E
0C5C
0C65
0C9A
0CDF
0CEC
0CA7
0C46
0C13
0C33
0C88
0CB4
0C60
0B9D
0AFC
0B01
0B82
0BC1
0B64
0B00
0B6B
0C9A
0D86
0D4A
0C2E
0B69
0BBF
0C79
0BDB
08E6
04AD
0199
0127
0270
0334
027B
01A8
027E
0458
0447
0046
F9D3
F4A2
F2F7
F3DD
F4E2
F4E1
F48F
F4C7
F539
F50E
F434
F384
F3AB
F469
F4F4
F4CD
F433
F3D6
F427
F4E1
F54F
F525
F505
F5EC
F7FD
FA29
FB30
FAF9
FA8E
FAC2
FB45
FB4A
FAB2
FA30
FA5E
FB1A
FBC5
FBF2
FB9E
FB00
FA5D
F9FE
FA02
FA38
FA55
FA5D
FA98
FB10
FB6B
FB63
FB2C
FB0F
FAF9
FABA
FA9A
FB21
FC11
FC2B
FA71
F78E
F550
F4C2
F545
F5BF
F5F2
F627
F61A
F549
F46A
F584
F9D3
FFE0
0490
061D
057A
04A8
0478
0474
043C
041E
0450
0483
0479
0479
04C4
04F9
04A5
0435
0476
052E
0507
0384
024B
0398
0782
0BAF
0DDB
0DFF
0D95
0D6F
0D23
0C61
0BCE
0C0B
0CA9
0CBC
0C2D
0BB5
0BC0
0BF5
0C09
0C5F
0D55
0E60
0E73
0D56
0C08
0B91
0BDE
0C24
0BFF
0BBE
0BAC
0BA7
0B82
0B79
0BD2
0C2C
0B80
0918
0596
02B9
01EA
02E1
03F4
03D6
0306
031D
047F
0537
02C4
FD1E
F73E
F433
F435
F505
F4CF
F3E5
F38E
F40B
F47F
F468
F446
F49F
F51C
F51C
F4AE
F471
F4A2
F4DE
F4C5
F476
F456
F4B0
F5AF
F755
F941
FAB1
FB21
FAEB
FAD1
FAF1
FAAE
F9C9
F915
F97B
FAB6
FB97
FB6D
FABC
FA63
FA91
FAD0
FAD6
FAD5
FB05
FB49
FB67
FB59
FB31
FB0A
FB20
FB9E
FC26
FC09
FB3D
FABA
FB3C
FC00
FB6F
F928
F6B4
F5B7
F5FE
F615
F57E
F520
F572
F586
F4D0
F4E3
F7ED
FDA8
02F5
051A
0489
03C4
0432
050C
053E
04EC
04B6
047B
03E3
035D
039F
0453
0461
0396
0315
03B2
0497
046F
038A
03D4
0667
0A04
0C94
0D6E
0D87
0DC0
0E06
0DEF
0D7B
0CF2
0C89
0C5F
0C8D
0CD8
0CB5
0BF4
0B51
0BB6
0CE0
0D78
0CC9
0BB6
0B87
0C3A
0CC5
0CA7
0C67
0C7C
0C7B
0BDF
0B14
0B1D
0C2D
0D29
0CC1
0A9E
0760
041D
0205
01D2
02F0
03B7
0323
021D
0234
0326
0295
FEC3
F90A
F4BC
F3A6
F483
F512
F4B1
F45D
F4C5
F56F
F593
F50D
F44D
F3CB
F3BF
F412
F462
F44D
F3F1
F3E5
F468
F4E0
F4B5
F490
F5D0
F891
FB11
FBB6
FAFF
FAAA
FB47
FBAD
FAEA
F9B8
F974
FA34
FACA
FA8B
FA1A
FA31
FA8B
FA8E
FA57
FA59
FA70
FA25
F9AF
F9E0
FAEE
FBF8
FC26
FBBD
FB97
FBDA
FBE6
FB7F
FB34
FB5D
FB76
FAED
F9F1
F8D4
F764
F58F
F44D
F4B5
F628
F692
F52F
F439
F6B2
FC93
0271
053A
052F
048F
047F
0471
03FE
03D2
0462
04F4
049D
03AA
0334
0385
03CE
0387
032E
0348
037E
0353
031E
0371
03F4
03CE
0339
03A9
060D
096A
0BDD
0CAC
0CB6
0CE3
0D12
0CCE
0C5E
0C5E
0CC6
0D0A
0CFD
0CFC
0D35
0D55
0D12
0CAA
0C87
0CA9
0CBC
0CA8
0CAF
0CF7
0D42
0D51
0D2F
0CFB
0CBE
0C9D
0CC5
0CF9
0CAD
0BF6
0BC3
0C8D
0D0C
0B45
0716
0301
0193
0284
0361
02E1
0234
0278
0257
FF81
FA1E
F540
F38A
F468
F544
F4C4
F3DF
F3EF
F4C3
F52D
F4B8
F401
F3B7
F3E6
F438
F45F
F439
F3E4
F3C1
F41E
F4D7
F579
F5CC
F5FF
F637
F64F
F64F
F6DC
F88C
FACB
FC18
FBB4
FA8D
FA04
FA4A
FA89
FA63
FA66
FAFF
FBA3
FB93
FB01
FAD0
FB3D
FB86
FB19
FA71
FA54
FAB0
FAD7
FA96
FA71
FACD
FB67
FBBB
FBA0
FB43
FACE
FA6D
FA70
FB0D
FBDB
FC03
FB10
F953
F765
F5AF
F489
F44E
F4CA
F518
F4B6
F4A7
F6BE
FB6A
00AE
03D7
041F
031E
02C4
037B
0478
050A
0516
04A9
03E4
0337
0328
03AF
0437
0454
0433
0418
03DA
0343
02BE
02E9
038E
03B5
032F
0359
05A0
097C
0CC5
0E06
0DD7
0DBA
0E1D
0E39
0D91
0CD1
0CCC
0D46
0D42
0C66
0B73
0B4B
0BF1
0CAE
0CFC
0CF6
0CFA
0D02
0CAB
0BDB
0B26
0B3D
0C12
0CD0
0CC5
0C2F
0BD4
0BF5
0C14
0BDD
0BCE
0C5B
0CB1
0B41
07C3
0404
0216
0226
02CC
0325
039A
044C
03C4
0051
FA94
F58A
F39A
F43D
F51D
F4E3
F42D
F405
F46A
F4B0
F49A
F484
F4AA
F4D9
F4F0
F527
F5A2
F609
F5EA
F550
F4BC
F485
F491
F49A
F482
F47B
F4F5
F650
F861
FA58
FB53
FB32
FAB1
FA96
FAEE
FB35
FB28
FAFF
FAF2
FADB
FAA1
FA84
FABB
FB09
FB0D
FAE5
FB05
FB82
FBD5
FB83
FAC9
FA50
FA5F
FAAC
FAEF
FB2E
FB6C
FB75
FB35
FAF0
FAE3
FAE3
FAA9
FA33
F982
F84B
F66F
F4A3
F403
F49D
F50C
F451
F3B9
F5E1
FB71
01B9
053B
0526
0399
02D5
032F
03C9
0437
04A8
04F6
0490
037F
02A9
02B8
033F
0379
036E
03B6
045C
04BF
0493
0460
04A5
0509
04EB
049D
056B
080C
0B7A
0DBC
0DD9
0CAB
0BCB
0C03
0CD2
0D3B
0CE1
0C4D
0C27
0C62
0C5C
0BCC
0B27
0B09
0B7D
0C16
0C8F
0CF6
0D3F
0D23
0CAB
0C74
0CEC
0D7B
0D34
0C41
0BD5
0C5F
0CC1
0BF9
0ADB
0AFF
0C24
0BF2
08FC
04FC
02DA
0308
0352
026B
01CD
0300
0456
025C
FC67
F60B
F342
F43A
F5D9
F5CE
F4A9
F40C
F43F
F471
F45F
F47B
F4C7
F4A6
F3FF
F3A6
F43E
F53A
F57D
F4C9
F408
F426
F4FE
F5A5
F57E
F4E2
F4D1
F620
F8A1
FB01
FBDF
FB3F
FA91
FAFE
FC0D
FC73
FBD3
FB1A
FB0E
FB45
FAF9
FA5E
FA5A
FB0B
FB6D
FADC
FA12
FA1E
FAE4
FB55
FAF0
FA4A
FA18
FA57
FAA7
FAFF
FB88
FC0E
FC1A
FB9F
FB1C
FAE1
FAAE
FA2E
F968
F86D
F729
F5D7
F525
F542
F52E
F3F7
F291
F39A
F886
FF6D
0487
05D6
04B4
03AB
03BE
0447
0497
04BA
04D7
04C7
047B
043B
042C
0415
03D1
03B3
0400
0445
03D7
02F5
02AA
034F
03EB
03B5
0390
052A
08B9
0C6D
0E44
0DFE
0CF1
0C66
0C92
0CFB
0D3B
0D2F
0CDE
0C86
0C67
0C63
0C1A
0BA1
0BA4
0C76
0D5C
0D5C
0C87
0BE3
0C1C
0CC6
0D19
0CF4
0CB9
0C7F
0C20
0BDC
0C2A
0CBE
0CA0
0BA5
0AE3
0B04
0ADF
08D1
0534
0256
01AE
0239
0258
0250
0365
04CB
0375
FDEC
F705
F32E
F392
F545
F54A
F3DE
F337
F427
F541
F520
F422
F37B
F389
F3D7
F431
F4C0
F55B
F58A
F553
F552
F5D4
F649
F5F3
F4EE
F43C
F4C8
F69C
F8F3
FAD5
FB9F
FB52
FA9D
FA56
FAB5
FB35
FB5B
FB47
FB3D
FB19
FA98
F9FC
F9DE
FA58
FAD6
FADD
FAB0
FAD3
FB2A
FB24
FAB0
FA7D
FAF2
FB90
FBA7
FB52
FB2D
FB64
FB96
FB85
FB6C
FB81
FB87
FB13
F9F5
F843
F644
F4A9
F470
F5BD
F703
F665
F45B
F400
F7CD
FE7C
041D
0629
0595
04CF
04CE
04E6
04C3
0512
0608
0694
05BE
0414
02E2
0288
0270
0268
02E7
03F1
049A
043D
0383
0382
0419
0432
03AE
040D
0689
0A35
0CE0
0D7D
0CDE
0C41
0BF7
0BBF
0BA5
0BF6
0C88
0CC3
0C70
0C18
0C3E
0CA8
0CB2
0C2D
0B8C
0B54
0BB0
0C6A
0D1A
0D69
0D5D
0D40
0D24
0CC1
0BEF
0B11
0AAC
0AB1
0A94
0A52
0AB7
0C1B
0D24
0BE1
0844
049A
0301
032B
0366
0327
0340
03A7
0277
FE25
F80E
F38D
F270
F358
F3F0
F3AD
F394
F412
F45B
F3DC
F338
F353
F414
F4A4
F4A6
F48C
F4C6
F523
F54B
F55E
F5B5
F639
F66C
F609
F551
F4E1
F558
F6EF
F91F
FAD1
FB4C
FAEB
FAA1
FAD9
FB10
FAB9
FA22
FA09
FA82
FADD
FAC7
FAC4
FB4D
FBEF
FBEB
FB50
FAE2
FB07
FB4D
FB2E
FACB
FAA6
FAEB
FB6B
FC05
FC9F
FCBF
FBE2
FA6C
F9A3
FA45
FB7D
FBC8
FA89
F860
F645
F4E1
F4AA
F5C2
F75F
F803
F71E
F655
F829
FD09
0274
0577
057C
0438
035D
0343
0387
03F4
0473
04BE
04AB
048D
04B9
04DC
0469
03A0
0374
0429
04BB
0449
0368
034B
03F3
0430
0392
0375
0578
0949
0CBB
0E09
0D7D
0CA4
0C7B
0CD7
0D1B
0CEC
0C5D
0BD8
0BE4
0CA0
0D76
0DA7
0D11
0C52
0C01
0C1A
0C3C
0C44
0C5A
0C81
0C86
0C5F
0C3E
0C25
0BDB
0B72
0B5E
0BBF
0C14
0BFD
0BE8
0C41
0C3C
0A5C
0685
02CC
0168
022E
0305
02C0
023B
0243
01A7
FEA6
F9BA
F58F
F406
F44E
F46A
F3D1
F38F
F431
F4D4
F496
F3F1
F3F7
F4BC
F565
F569
F510
F4B4
F454
F40D
F450
F53A
F60A
F5D6
F4C0
F403
F4A4
F66D
F866
F9D2
FA84
FA96
FA5F
FA6F
FB0F
FBD0
FBF4
FB54
FA8E
FA4F
FAB0
FB4F
FBD5
FC0F
FBCA
FAFE
FA2D
FA06
FA87
FAEB
FABA
FA6F
FAB2
FB5F
FBBF
FB96
FB53
FB48
FB4B
FB3B
FB77
FC3D
FCE6
FC6A
FAA5
F885
F6D6
F5A1
F4E5
F511
F60D
F6A3
F5F6
F558
F763
FCC7
02CF
05FA
05AF
0460
0429
049A
0449
0343
02D3
0372
0432
0440
03EB
03D7
03F1
03CB
038B
03B4
0430
0457
0408
03E9
0438
0442
03B2
03BC
05D4
0976
0C44
0CA6
0B9C
0B58
0C92
0E00
0E4F
0DAD
0D17
0CD9
0C86
0BFB
0BAE
0BE9
0C58
0C87
0C6B
0C4E
0C69
0CB0
0CF3
0CFE
0CB7
0C3A
0BD4
0BAB
0B82
0B1F
0AD3
0B38
0C31
0CB4
0BCD
09A2
0710
04BC
02F5
022F
02BB
03B8
0317
FF84
FA33
F5F7
F460
F456
F3E9
F2C1
F210
F291
F387
F3F0
F3D3
F3E8
F455
F486
F439
F405
F487
F562
F5A8
F50B
F436
F3FB
F467
F4DE
F4DE
F4A6
F50E
F6C2
F980
FC22
FD7B
FD35
FBF0
FA8C
F993
F936
F999
FAA5
FBBD
FC15
FB93
FAFF
FB0F
FB92
FBD3
FB99
FB4B
FB31
FB11
FAB8
FA7C
FACC
FB6F
FBC0
FB92
FB52
FB35
FAEC
FA7B
FAA7
FBDB
FD01
FC62
F9CB
F704
F5AC
F554
F4A1
F3F9
F5A5
FAD2
0159
059D
0631
04CF
03D3
03CB
03DC
039F
038F
03F3
044B
0437
042A
04AB
0559
055B
0496
03DD
03DF
046C
04E6
0507
04D7
0453
03AA
03A7
053F
085A
0B85
0D45
0D82
0D49
0D5C
0D80
0D30
0C7A
0BE2
0BAA
0BAA
0BB3
0BC6
0BE4
0BE7
0BCA
0BD0
0C20
0C7E
0C95
0C72
0C5D
0C54
0C06
0B73
0B1C
0B67
0BFC
0C2D
0BF1
0BFD
0C9D
0CE4
0B76
081E
0441
01B7
014D
025C
0363
02E0
0006
FB51
F686
F3A9
F36E
F4B3
F5AE
F593
F4F2
F49D
F4A9
F4A9
F478
F461
F489
F4AA
F480
F43C
F434
F455
F441
F3FD
F413
F4D7
F5BE
F5EA
F554
F507
F5FD
F7FE
F9DD
FAC1
FAD4
FAAE
FA89
FA44
F9FC
FA18
FAAE
FB3C
FB4E
FB25
FB63
FC22
FCC8
FCD0
FC71
FC2E
FC09
FB95
FAD1
FA6C
FAEC
FBE9
FC7E
FC5A
FBF8
FBBF
FB7D
FB03
FAC5
FB2F
FB96
FA9B
F804
F578
F4C3
F59D
F623
F5A2
F5FC
F96C
FF5B
0466
05E1
0479
02EB
02CB
0369
038F
033B
0330
0395
03DF
03D0
03D0
0417
0442
040C
03E4
0448
04F3
0540
0517
04D8
0481
03BC
030C
0414
07B8
0C57
0EF0
0E61
0C99
0C17
0D06
0DAB
0D17
0C38
0C2F
0CBC
0CE6
0C93
0C81
0CDC
0CE5
0C2F
0B74
0B8A
0C24
0C4F
0BD4
0B5E
0B6A
0BBB
0BE4
0BD8
0BA7
0B3A
0AB2
0AB2
0B98
0C83
0BE0
093A
05E2
037F
0294
02B0
0359
03D3
02AB
FEBA
F903
F489
F37E
F4EA
F5F4
F543
F420
F41A
F4CF
F4D3
F3F9
F374
F3F9
F4CF
F503
F4BA
F4B9
F514
F528
F4AD
F433
F43B
F47C
F471
F44F
F4CA
F624
F7E4
F966
FA53
FA9A
FA69
FA2C
FA4B
FAB6
FAE6
FA82
F9ED
F9E5
FA9A
FB6C
FBA8
FB40
FAB2
FA7A
FAD1
FB9C
FC5C
FC7E
FBF5
FB5C
FB3E
FB7D
FBA9
FBB2
FBE7
FC3C
FC39
FBC7
FB87
FBBF
FB64
F94B
F646
F4B6
F57F
F698
F5CF
F445
F588
FAFF
01A0
0521
04A4
02FE
02C3
03AB
0433
0434
048C
0526
04F7
03DE
0329
03D3
0516
0577
04B0
03CD
03A8
0414
049D
0517
0537
048B
0392
03FA
06CD
0AAF
0D12
0D1C
0C72
0CE0
0E13
0E74
0D9D
0CD3
0D04
0D8F
0D7E
0D0F
0D10
0D68
0D45
0C80
0BDA
0BBA
0B97
0B0D
0ABA
0B47
0C10
0BC2
0A5B
097E
0A42
0BB0
0C2E
0BB9
0BA8
0C65
0C92
0ACD
077A
0453
029C
026A
0334
0413
0375
FFE6
F9F6
F49A
F291
F38F
F4DD
F4A0
F39A
F36D
F42C
F48E
F418
F3D7
F4AB
F5D4
F602
F541
F4E1
F585
F63F
F5EE
F4D7
F441
F4B7
F55B
F530
F495
F501
F729
F9F2
FB74
FAF8
F9AA
F948
FA3D
FB53
FB38
FA18
F954
F9C5
FAD6
FB7C
FB7B
FB64
FB88
FB8C
FB24
FAA4
FA96
FAE7
FAFF
FA9E
FA2B
FA20
FA88
FB28
FBC5
FC06
FBA2
FAE7
FAAD
FB26
FB2A
F96A
F66E
F471
F4B7
F5D5
F5A4
F4A7
F5EF
FB21
01CB
05CE
05DD
0454
03DB
0483
04CC
0449
040C
04B6
0579
056B
04D3
047C
047E
0468
043A
044D
0477
0431
039A
0388
042B
047E
03C6
033D
0504
0944
0D64
0ED0
0DC1
0C8D
0CA4
0D51
0D56
0CA9
0C1E
0C08
0BFA
0BB1
0B83
0BC4
0C41
0CA3
0CDF
0CF2
0CAB
0C1F
0BEB
0C6B
0CF4
0C8B
0B50
0A96
0B43
0CA5
0D5C
0D16
0CA6
0C82
0BF9
0A4B
07D1
0584
03F2
032F
0354
041C
041E
0188
FC4C
F6E5
F423
F44E
F538
F521
F47C
F481
F508
F4E9
F3F7
F35B
F3D5
F4A4
F4C5
F48A
F4FA
F5F8
F61F
F4D6
F37F
F3D2
F580
F683
F5C0
F472
F495
F688
F8D9
FA1C
FA49
FA34
FA40
FA28
F9D5
F9BE
FA38
FAE9
FB1E
FAB5
FA4F
FA8E
FB40
FB8C
FB02
FA39
FA13
FA9F
FB0F
FAD9
FA6E
FA83
FB09
FB49
FB00
FAC0
FAFD
FB3D
FAD9
FA35
FA3E
FAB7
FA1D
F7CB
F555
F4C2
F5CE
F645
F553
F540
F8BA
FF04
0441
05B8
0487
0389
03C3
0411
03A8
034E
03E1
04D6
050B
047B
0422
0465
048F
0419
039F
03EE
04C5
053F
0501
046F
03E8
0397
03FA
05C1
08C7
0BB2
0D21
0D13
0C9D
0C6F
0C4E
0C0F
0C38
0D1A
0DF7
0DD3
0CCB
0BE8
0BC3
0BFE
0C20
0C4E
0CB6
0CEF
0C7C
0BBE
0BA0
0C3B
0C9E
0C35
0BAE
0BDB
0C56
0C2D
0B7D
0B6F
0C66
0D10
0BDA
08E0
05C9
03EC
0359
0398
0454
04B8
0316
FE75
F846
F3A7
F278
F3B6
F4ED
F4DA
F436
F427
F4BB
F527
F4FE
F492
F456
F454
F45C
F46B
F4A4
F50F
F57A
F5A2
F580
F55D
F575
F599
F576
F53E
F5C9
F7A2
FA0D
FB5F
FAAC
F8E6
F7F6
F8BC
FA58
FB6A
FB89
FB30
FACE
FA77
FA4F
FAA4
FB68
FBFA
FBC8
FB07
FA70
FA5E
FA84
FA88
FA7B
FA8E
FAAA
FA9B
FA6C
FA49
FA31
FA20
FA55
FAFA
FB83
FAEA
F8E4
F687
F537
F503
F4C6
F411
F446
F71D
FC63
01C0
04E6
057B
04D0
0440
0434
0476
04C1
04E2
04C2
0497
04CD
056B
05CD
0561
047B
0400
044F
04D3
04DF
0477
0404
038C
02D4
024C
031E
05DF
098B
0C59
0D68
0D43
0CE1
0C9E
0C61
0C43
0C7F
0CFC
0D4B
0D3D
0D17
0D0A
0CE3
0C7F
0C2B
0C38
0C70
0C68
0C31
0C3F
0C9A
0CA7
0C15
0B88
0BD4
0CB0
0CFE
0C66
0BF0
0C7C
0D4B
0CAB
0A06
0696
0410
033B
03C2
04CA
051B
0353
FEF4
F969
F535
F3AA
F3DD
F435
F452
F4C6
F577
F560
F418
F2BD
F2AA
F3C5
F4BC
F4D5
F4A5
F4E2
F539
F4F6
F456
F456
F547
F645
F651
F58A
F519
F603
F820
FA43
FB36
FAB3
F993
F90E
F9A0
FAAD
FB4A
FB47
FB2B
FB38
FB0A
FA60
F9C3
F9DA
FA7D
FAEF
FAE4
FAD2
FB12
FB50
FB1C
FABD
FAD3
FB4F
FB6E
FADA
FA3B
FA49
FACD
FB0D
FACB
FA3E
F962
F800
F677
F5B6
F602
F64E
F59F
F4E0
F66F
FB4B
0161
054F
05B3
042C
0337
03B1
049B
04CA
043D
03DB
042A
04C0
04D1
0433
0387
0371
03DE
042B
0405
03D0
03F8
042D
03DC
0371
045C
0765
0B4D
0DD0
0DEE
0CCC
0C2D
0C97
0D42
0D71
0D4A
0D3E
0D45
0D0B
0C9A
0C4A
0C36
0C14
0BBA
0B6F
0B98
0C35
0CE0
0D39
0D38
0D15
0CE2
0C7F
0BEE
0B98
0BF4
0CDD
0D63
0C70
09CE
0673
03C9
02A8
02F1
03CC
03E3
01D2
FD2E
F777
F360
F27B
F3BB
F4B5
F445
F371
F3A2
F4B6
F566
F527
F4BF
F4E5
F528
F4C3
F3F6
F3C7
F496
F5AA
F61B
F5CC
F530
F4B3
F49E
F54E
F6FA
F91F
FAAF
FB13
FACB
FAC3
FB4B
FBF6
FC42
FC14
FB98
FB0D
FAB2
FAB3
FB09
FB7C
FBCA
FBC3
FB4B
FA7D
F9D1
F9DF
FAC1
FBBE
FBF4
FB52
FA9B
FA63
FA74
FA71
FA7D
FACD
FADE
F9DD
F7E8
F63F
F5D2
F60C
F5BC
F525
F64A
FA93
0098
050E
05EE
044C
02D3
02EC
03D3
0427
03C2
039F
0445
0500
04D9
03F4
0354
0384
0401
042A
0438
04BC
0576
0565
0444
036E
049B
07D0
0B31
0CFA
0D1E
0CC3
0CAA
0CB0
0C87
0C40
0C12
0C08
0C1F
0C6C
0CE0
0D21
0CE7
0C79
0C71
0CEF
0D6B
0D60
0CE8
0C6A
0C1C
0C0C
0C4D
0CB4
0CC3
0C45
0BC8
0C02
0CB3
0C84
0A5F
06BC
034A
017A
0190
02BE
0383
021A
FDB7
F7DE
F3A9
F2EA
F450
F51E
F457
F360
F397
F465
F461
F381
F31A
F3C3
F479
F449
F3BC
F3E0
F4A7
F52B
F515
F4D6
F495
F407
F384
F458
F72B
FA98
FC47
FB8A
FA0F
F9B1
FA71
FB0F
FAFE
FAC8
FAEF
FB4C
FB95
FBCB
FBED
FBBB
FB1E
FA80
FA69
FACA
FB23
FB40
FB64
FBA9
FBB9
FB6C
FB16
FAEA
FA95
F9F6
F9AE
FA3E
FADE
FA1B
F7DC
F5E5
F5B8
F682
F640
F4F2
F54F
F98D
003C
0563
069E
052B
03D6
03D7
0447
0415
0384
037D
0430
04E1
04E4
044C
03A2
0351
0377
03F3
0487
04ED
04EC
0479
03E6
03F3
056F
086B
0BD1
0E07
0E3D
0D27
0C3D
0C50
0CEC
0D2B
0CCF
0C53
0C27
0C33
0C29
0C0D
0C28
0C8F
0CF0
0CED
0C93
0C4C
0C57
0C81
0C7F
0C62
0C6A
0C86
0C57
0BD5
0B99
0C21
0CE6
0C97
0A64
06F6
03DF
024B
025B
036D
044A
0350
FF6B
F986
F470
F27F
F362
F4C6
F4FA
F45E
F42D
F497
F4CF
F47A
F432
F46E
F4C0
F49B
F43B
F438
F4A9
F536
F59E
F5B4
F526
F40E
F382
F4D2
F7D5
FA88
FB09
F9A9
F885
F90B
FAA8
FBFC
FC6A
FC18
FB30
FA04
F952
F9A0
FA6E
FAC4
FA75
FA33
FA5F
FA7C
FA1F
F9E1
FA9D
FC06
FCD8
FC83
FBC9
FB6B
FB29
FAA4
FA5B
FAC6
FB06
F9BD
F726
F535
F52B
F5E8
F588
F454
F4F1
F935
FFA0
04A8
0643
0575
049F
04F1
05B4
0591
0441
02EB
02E1
0416
052D
050C
040D
0355
036A
03D4
040E
043A
048F
04AF
0439
03E5
0512
07F6
0AFF
0C8E
0CBB
0CCF
0D56
0DA7
0D33
0C75
0C39
0C7C
0C92
0C39
0BE9
0C09
0C66
0CAB
0CE5
0D26
0D20
0C91
0BE6
0BCE
0C53
0CB9
0C5E
0B68
0A89
0A5A
0AF2
0BF8
0CC1
0C88
0ADB
0807
0506
02E9
0255
033F
0489
0423
0078
FA4F
F4B4
F242
F2C1
F3E6
F421
F3E3
F421
F4A5
F497
F428
F474
F5B4
F691
F5E8
F468
F3A7
F419
F4DB
F52F
F547
F56F
F560
F4EC
F4D0
F61F
F8C4
FB39
FC14
FB73
FA9B
FA76
FAD9
FB15
FAC1
FA10
F998
F9C7
FA65
FAD5
FAD5
FACA
FB0C
FB55
FB33
FAD3
FADD
FB65
FB93
FACB
F9BE
F9B6
FACD
FBB6
FB8E
FB04
FB1E
FB78
FAAD
F865
F5FA
F4D6
F4D3
F4D0
F4A4
F5A6
F90D
FE21
02A0
04DF
0525
04EF
0520
0552
04C6
03B3
0344
0420
055F
0576
042A
02FE
0359
04CE
05B7
0546
0454
040C
046A
048E
0441
0473
0605
0898
0AFA
0C77
0D42
0DBE
0DD5
0D49
0C57
0BBB
0C05
0CEA
0D7A
0D23
0C5C
0C34
0D0C
0E0B
0E01
0CBA
0B3B
0A9A
0ADE
0B40
0B49
0B3F
0B72
0BB5
0BBE
0BBF
0C0F
0C71
0C0B
0A41
0753
042F
01DB
0125
0240
041E
046C
013B
FB1F
F53E
F293
F341
F4E8
F557
F474
F387
F36D
F3F4
F491
F506
F538
F51A
F4EE
F516
F571
F55A
F4AC
F42F
F48A
F53B
F550
F4ED
F556
F734
F985
FACE
FAEA
FAE8
FB45
FB5D
FAC0
FA16
FA17
FA71
FA88
FA92
FB1D
FBD1
FBBA
FABB
F9E9
FA2A
FB10
FB88
FB3C
FA9C
F9F9
F980
F9E4
FBA3
FD7E
FD37
FAB9
F901
FA73
FD42
FD4B
F964
F4F7
F3AB
F504
F5BB
F4AD
F476
F7B2
FD7C
02B8
059E
0692
065E
0548
03E8
0363
0432
0559
057E
0483
038D
03A0
0490
0561
0564
04B3
03F6
03E1
0489
052B
04EC
0424
0454
0670
09A1
0C3A
0D7E
0DD8
0DB1
0CF6
0BDD
0B60
0C30
0D8E
0DF0
0CE3
0BAC
0B9C
0C62
0CA5
0C00
0B83
0C0F
0CFE
0CFE
0BE8
0B11
0B95
0CCF
0D12
0BDF
0AAE
0B12
0CA1
0D63
0C34
09D0
075C
04F8
0279
00D4
0170
03B1
046E
00EF
FA3C
F467
F266
F37E
F4F8
F54D
F4EF
F4B6
F4C5
F4D3
F4B7
F467
F3F8
F3C9
F444
F532
F5AF
F52E
F450
F41C
F48E
F4AE
F438
F42C
F557
F720
F889
F99C
FAF2
FC3B
FC68
FB4A
FA1F
FA00
FA7F
FA83
FA15
FA42
FB47
FBF5
FB75
FA9B
FAA5
FB6A
FBBA
FB21
FA5B
FA1C
FA53
FABC
FB58
FBF1
FBC8
FA89
F944
F97B
FB09
FBEF
FAA4
F7F8
F5E7
F53B
F528
F4F1
F4F5
F615
F8B7
FC9C
010B
04CE
0680
05BB
03E3
030D
03D1
04C0
046E
0362
0343
047A
0593
0522
0392
0292
030F
045A
0532
0527
04AA
043B
040C
0463
05CC
0873
0B8D
0DC7
0E61
0DCA
0D0A
0CC1
0CC8
0CBB
0C8A
0C7B
0CAE
0CD1
0C7B
0BC9
0B72
0C10
0D4B
0DEF
0D21
0B7A
0AA5
0BA4
0D8D
0E6F
0D70
0BB4
0AFD
0BC2
0CED
0D28
0BFD
09D1
0745
04F1
0361
02E0
031E
032B
020B
FF66
FBB6
F7F1
F514
F3A6
F381
F409
F4AB
F514
F501
F45E
F39D
F38E
F474
F586
F5C2
F516
F461
F462
F4ED
F55E
F562
F529
F4EB
F4C2
F4F8
F604
F7E6
F9DC
FB09
FB36
FACC
FA6A
FA9B
FB81
FC78
FC8A
FB89
FA68
FA1E
FA89
FAD9
FACA
FACE
FB00
FAC5
F9F4
F9A9
FAD9
FC75
FC5E
FA6C
F909
F9FF
FBF5
FC62
FB1D
FA4E
FB02
FB8A
F9F6
F6F6
F4E5
F48F
F47B
F3C9
F41A
F77D
FD3E
0234
0424
03CB
0350
03B9
0455
0439
038B
033E
03C7
0485
048E
03D9
0358
03CA
04CA
0531
0467
0318
0275
02F2
041F
058F
0769
09BE
0BE7
0D0D
0D34
0D2B
0D73
0DA8
0D3C
0C7E
0C66
0D4D
0E2E
0DAA
0BD9
0A86
0B2E
0D11
0E03
0D1A
0BC8
0BEC
0D6F
0E8F
0E2C
0CF7
0C22
0BDE
0BD7
0C4F
0D53
0D39
09D1
03D6
FF83
0039
043F
065B
0391
FDEC
F95A
F72C
F5D7
F429
F2E8
F315
F42F
F508
F55B
F580
F560
F4C8
F459
F4E0
F5DD
F5DA
F486
F371
F40A
F581
F5CC
F48F
F3B9
F4E3
F74A
F924
FA10
FAFB
FC1D
FC75
FB83
FA66
FA7A
FB8A
FC2B
FBB7
FB02
FAED
FB2B
FAFC
FA86
FA97
FB56
FBE8
FB84
FA60
F970
F986
FAB4
FC35
FCD8
FBF2
FA36
F94B
FA0C
FB3F
FACD
F84E
F591
F462
F4AE
F56F
F6B1
F960
FD54
00D8
02AB
0387
04C1
05FD
059A
0379
01D9
02A2
04C7
05A3
0476
0327
0372
04A0
04D6
03D6
0337
03EA
04C9
044B
02F5
0302
05AE
09AC
0CA3
0D9A
0D5B
0CF2
0C89
0C02
0BCC
0C89
0DE2
0E7B
0D6E
0B8E
0AA5
0B83
0D1B
0DAF
0CA5
0B06
0A5A
0B3F
0CF3
0E03
0D86
0BE4
0A96
0AE3
0CBD
0EAE
0EE4
0C8B
0876
04A6
02E3
0368
04A9
048D
0228
FE55
FAA0
F7BC
F563
F37D
F2A5
F346
F4A7
F574
F50E
F40A
F36A
F3B5
F4A5
F57A
F59E
F52D
F4DA
F525
F5AB
F588
F47E
F37E
F3AA
F4FD
F680
F7BC
F927
FAE6
FC0C
FBCB
FAC3
FA54
FAE1
FB86
FB81
FB21
FB12
FB49
FB2B
FA98
FA3F
FAAF
FB8F
FC03
FBA8
FADD
FA53
FA89
FB58
FBEB
FB87
FA91
FA3C
FAF9
FBB8
FB46
F9CA
F84F
F72D
F5C9
F420
F397
F59B
F9BC
FE06
011E
0336
04BC
053B
0451
02FF
02D9
0408
0511
04C9
03BE
0355
03F0
048A
042A
0335
02EC
03B8
048D
0435
02FD
0285
03FB
06DF
09AD
0B73
0C67
0CFB
0D0B
0C65
0BB6
0C08
0D3B
0DEA
0D32
0BE6
0B77
0C34
0D38
0DA7
0D62
0CA7
0BD2
0B82
0C41
0DAB
0E4F
0D27
0B16
0A36
0B80
0DB2
0EC8
0DEA
0B93
089D
05DD
0421
03A4
03AA
0312
015B
FEB0
FB4E
F779
F410
F261
F2DC
F445
F4EE
F496
F45A
F4CF
F52D
F4C7
F448
F4A7
F581
F59C
F4BA
F3F7
F42E
F4DB
F506
F4A9
F49E
F558
F678
F7AC
F931
FB0E
FC76
FC89
FB7A
FA5D
FA06
FA83
FB69
FC2A
FC28
FB25
F9CC
F963
FA7D
FC25
FCB8
FBAC
FA33
F9D8
FACC
FBDE
FBE2
FADD
F9CE
F9AA
FA84
FB87
FBC7
FB19
FA0E
F90D
F7CE
F5F4
F40D
F38F
F59E
F9DF
FEB2
0276
047A
04F1
0489
041C
043C
04AB
049F
03E3
0355
03DB
0502
0551
0420
029E
0287
040B
0586
055E
03C6
025E
0273
0413
0678
08D9
0AB9
0BDB
0C42
0C36
0C2A
0C70
0CEC
0D24
0CC7
0C26
0BF6
0C7C
0D25
0D21
0C62
0BAB
0B92
0BD0
0BCF
0BB4
0C22
0D0B
0D62
0C88
0B64
0B6B
0CC6
0DF7
0D80
0B52
0888
0626
0483
03A6
0380
037A
0251
FF08
FA19
F55F
F2A4
F244
F334
F424
F48C
F4B3
F4E1
F4D3
F446
F3B6
F3FA
F514
F5E9
F593
F493
F437
F4E6
F5A6
F583
F4E0
F4E4
F5E0
F6FE
F7A5
F85E
F9DE
FBB2
FC94
FBFB
FABF
FA28
FAAC
FBBB
FC71
FC56
FBAB
FB1A
FB21
FB98
FBD2
FB5F
FAA5
FA78
FB07
FB85
FB21
FA29
F9C7
FA9D
FBF7
FC8A
FBDC
FABF
FA56
FAA5
FA67
F878
F564
F343
F3E7
F73D
FB97
FF51
01F4
03D3
0503
0547
04B1
03E4
0373
0377
03CF
047A
0544
057A
0495
0332
02C1
03E2
0563
0586
0417
029F
0278
035D
0456
0557
0728
09E2
0C5F
0D73
0D36
0C9D
0C2A
0BB0
0B3E
0B6C
0C6B
0D64
0D61
0C8D
0BEF
0C21
0CB5
0CDE
0C55
0BA0
0B87
0C40
0D0E
0CE6
0BA5
0A88
0AF4
0CB7
0DF3
0D26
0AE2
08D3
076F
05CD
03C6
029D
02C3
0243
FEEB
F963
F4C0
F304
F344
F38C
F376
F3D8
F4B1
F4E1
F411
F37C
F41A
F514
F50A
F425
F3C5
F484
F59C
F615
F5C1
F513
F499
F4A1
F524
F5F1
F716
F8D6
FB06
FC9E
FC88
FAF6
F99F
FA08
FBC5
FD02
FCC8
FBC6
FAEC
FA54
FA04
FA5F
FB3C
FB9E
FB2E
FAFD
FBC8
FC7A
FBB9
FA3B
FA03
FB4C
FBEE
FA96
F93B
FA79
FD3D
FD6E
F977
F4BF
F350
F4FC
F6C0
F793
F954
FD59
0227
053F
05C9
04D9
03D5
0370
03C4
0497
0547
0520
043F
0391
03AA
042A
0489
04C5
04CA
042E
0320
02B4
0368
043B
042E
040F
0596
08F5
0C5C
0DFF
0DD5
0D12
0C8F
0C54
0C59
0CC4
0D4A
0D23
0C2A
0B5D
0BA2
0C8C
0D00
0C99
0BD7
0B59
0B6A
0C01
0CA6
0CBE
0C44
0BEC
0C24
0C82
0C87
0C69
0C70
0BE5
09A7
0603
031D
029F
0360
0267
FE6A
F92E
F530
F32D
F289
F2E3
F405
F511
F525
F489
F448
F4A9
F4E5
F478
F3E9
F3FA
F493
F501
F50A
F51B
F563
F570
F4F5
F46B
F479
F540
F69F
F878
FA51
FB47
FB23
FADE
FB68
FC54
FC74
FB86
FA94
FA93
FB49
FBAF
FB3A
FA5B
F9FA
FA9B
FBED
FCDC
FC59
FAA3
F999
FAB8
FCD1
FCFA
FA67
F80C
F91D
FCAD
FE7C
FC26
F7FD
F5D9
F653
F6C1
F5A4
F532
F86C
FEBE
042E
05B4
042F
02A9
02C5
03C4
0464
047F
0494
04AA
0469
03F6
03E2
044D
049D
044D
03A9
036A
03CF
0457
045D
03C8
0326
0363
053C
087C
0BAC
0D25
0CB8
0BEC
0C28
0D34
0DDC
0D9A
0D03
0CBD
0CC2
0CC3
0CB7
0CC0
0CC5
0C9E
0C78
0CAB
0D0F
0D1A
0CBA
0C77
0C91
0C85
0C01
0B9B
0BFC
0CD5
0D1F
0C27
09EE
070A
0482
0340
02E4
0192
FDB7
F82F
F3E9
F2F5
F455
F56D
F526
F49E
F4CC
F509
F47B
F3A3
F371
F3CD
F40E
F430
F47F
F4A4
F430
F3B0
F423
F566
F61B
F582
F4AE
F52E
F700
F8BC
F9A7
FA62
FB66
FC11
FBD9
FB43
FAE2
FA78
F9FB
FA42
FB87
FC49
FB2B
F95A
F967
FBAE
FD68
FC24
F926
F7F9
F9F3
FC93
FCDE
FAFD
F987
FA15
FBCE
FCF0
FCA7
FB4C
F9AC
F81C
F645
F427
F333
F571
FAEC
00D7
0414
043B
036B
037F
044D
04AC
0445
03BC
0384
0387
03DB
04B9
0589
0521
037E
0251
02E9
0475
0524
0461
030E
022C
0245
03B0
0656
0943
0B38
0BE8
0C26
0CBD
0D7A
0DA3
0D0E
0C4A
0BD2
0BC0
0C40
0D6B
0E7E
0E2A
0C5F
0ABB
0AA1
0B9F
0C76
0CC3
0CD6
0CAF
0C30
0BBE
0BD5
0C38
0C61
0C69
0CAF
0C97
0AC4
0731
041F
0376
03C3
019F
FC5B
F74B
F56D
F5BA
F545
F38E
F298
F377
F4D5
F51F
F481
F412
F41B
F423
F425
F49B
F560
F58A
F4E0
F45D
F4B6
F53B
F509
F49D
F52E
F6E5
F8B7
F9E2
FA9C
FB5C
FC11
FC3F
FB8E
FA34
F90D
F91F
FAAF
FCB8
FD95
FC87
FA96
F9AA
FAA0
FC64
FD28
FC48
FACA
FA27
FAD4
FBF1
FC38
FB59
FA57
FA54
FB09
FAFE
F956
F6CA
F4C1
F432
F5B7
F9AE
FF5D
0470
067F
055A
0338
025A
02FA
03D8
0433
045C
047E
0417
0314
0283
033E
047D
04A0
0355
0205
0217
035A
046B
0464
0402
04FA
080D
0BDE
0E19
0DCF
0C40
0B45
0B6F
0C0E
0C94
0D2A
0DDE
0DFE
0CFB
0B8C
0B0B
0BB5
0C72
0C8A
0C75
0CA4
0CA3
0C1E
0BBA
0C02
0C5E
0C1B
0BC8
0C48
0CDA
0B80
07E3
0477
0380
03CA
01FA
FD21
F813
F5A1
F532
F482
F33D
F2FC
F442
F582
F564
F47D
F41B
F45D
F46E
F423
F439
F4E1
F534
F4A0
F3FB
F442
F500
F4F4
F42A
F441
F64C
F947
FB2D
FB3A
FA79
FA44
FACB
FB53
FB69
FB4E
FB45
FB22
FAC0
FA80
FAD3
FB84
FBEE
FBE6
FBD5
FBE0
FB90
FAB3
FA12
FA9C
FC0B
FD04
FCB8
FBD6
FB83
FBBA
FB4E
F975
F6CC
F4BE
F47E
F6AA
FB10
0042
040C
052F
0485
03F1
0455
050B
051E
0472
03A5
033C
033A
0360
0385
03A0
03BA
03E7
0427
0444
0407
039A
0356
0348
0382
04BA
079B
0B3B
0D5D
0CFD
0BC3
0BFC
0DA5
0E9D
0D97
0BC5
0B1E
0BE1
0CB5
0CC1
0C72
0C39
0BD4
0B47
0B4F
0C0F
0C6A
0BA0
0ABA
0B29
0C88
0D10
0C2F
0B4A
0B78
0BA7
0A29
0751
050D
03D5
01B8
FD3D
F7F1
F4B8
F446
F4B6
F466
F3BE
F3CD
F463
F486
F424
F41C
F4B2
F50B
F49D
F437
F4C1
F5A6
F590
F47F
F400
F4EF
F60E
F5B6
F460
F44A
F687
F97C
FADD
FA5B
F985
F97F
F9E8
FA09
FA0D
FA81
FB39
FB7D
FB25
FAD7
FAFA
FB30
FB18
FAF9
FB36
FB7F
FB51
FADB
FACE
FB48
FB93
FB29
FA7A
FA72
FB49
FC03
FB38
F87F
F52B
F3AA
F5D7
FB4D
0158
04F6
054C
0400
032B
036F
042E
04BC
04DE
0495
0416
03CF
03F1
0427
0413
03E9
0428
04B1
04C6
0418
0369
0383
040C
043A
048A
0664
09CD
0CB5
0D73
0CD7
0CC2
0D72
0D8C
0C8B
0BB3
0C1F
0D10
0D1B
0C51
0C05
0C97
0CEB
0C54
0BAA
0BBB
0BF2
0B9D
0B6E
0C59
0D87
0D2B
0B68
0AA2
0C1B
0D97
0BF5
0790
03FE
0322
0273
FE8F
F81F
F33D
F26F
F41A
F537
F4E6
F45D
F466
F47D
F44E
F47A
F557
F5F9
F578
F472
F438
F4D9
F51E
F47F
F3F6
F477
F561
F55C
F462
F40E
F596
F839
FA2C
FAA6
FA5F
FA50
FAAB
FB09
FB22
FB08
FAF7
FB06
FB06
FAB8
FA2E
F9D7
FA09
FA93
FAEA
FAC6
FA73
FA6B
FAC4
FB3D
FBB0
FC0B
FC02
FB66
FACA
FAE1
FB11
F9AD
F664
F3C4
F51A
FAAF
011A
04A7
04D0
03DB
03B0
042A
0468
0455
0450
044A
0418
0401
0429
040E
0353
02AD
0310
0425
048A
03C5
030B
0377
0453
0448
03D8
0513
0877
0BC6
0CD7
0C5D
0C82
0DAF
0E48
0D76
0C78
0CA3
0D58
0D0C
0BC2
0B14
0BD6
0CF3
0D32
0CD5
0CB5
0CBF
0C74
0C2A
0C85
0D06
0C7B
0B22
0AE7
0CAE
0E59
0D03
08DE
052D
03E3
02DA
FECE
F826
F2F4
F222
F43C
F5AE
F50A
F3EB
F413
F529
F5BC
F568
F4FE
F500
F50B
F4C6
F484
F4A1
F4D3
F49A
F414
F3DB
F421
F46A
F461
F48E
F5C0
F7E0
F9C7
FA7A
FA2E
F9E0
FA1E
FA87
FA85
FA3A
FA56
FB18
FBD3
FBBA
FAEE
FA4D
FA5A
FAB3
FAD1
FACA
FB00
FB58
FB59
FB0C
FB2B
FBFB
FC96
FC09
FAE3
FA8B
FAF7
FA49
F78D
F4EF
F5DF
FB07
0120
0461
0448
0349
0366
044D
04CD
04AB
0464
0412
0394
0339
035F
0399
032B
024E
021B
02FC
03F4
0406
03A8
03E8
0485
044F
0380
042B
077C
0B9F
0DBC
0D5B
0C86
0CBE
0D51
0D06
0C3F
0C46
0D28
0D88
0CAE
0B8C
0B3E
0B99
0BF4
0C60
0D25
0DB6
0D59
0C7B
0C43
0CD0
0CFC
0C39
0BA8
0C67
0D7A
0CAA
098D
062B
0413
0211
FE1C
F8A2
F471
F35D
F446
F4D8
F43E
F37A
F393
F455
F4F9
F53A
F554
F560
F540
F506
F4E9
F4E4
F4C0
F483
F46B
F48E
F4B6
F49D
F44F
F44D
F546
F759
F995
FAA2
FA23
F937
F93E
FA46
FB12
FACA
FA15
FA1A
FAD1
FB2E
FACC
FA76
FABC
FB02
FAA3
FA26
FA6E
FB2F
FB49
FA9B
FA62
FB4F
FC45
FBE8
FAD4
FAC1
FB88
FAC4
F75E
F42D
F549
FB29
01D1
0523
04DA
03B6
03C3
04A0
0513
04E9
04BB
04B2
0487
0445
043E
0465
0450
03FB
03E0
042C
0460
040D
0386
0364
0396
038D
0367
043F
06D8
0A50
0CD1
0D7F
0D2E
0D1F
0D8A
0DBA
0D3D
0C7D
0C1D
0C3C
0C83
0CA8
0C9A
0C64
0C22
0C05
0C1C
0C2C
0BF9
0BB2
0BCC
0C4B
0C96
0C44
0BD8
0C1C
0CD5
0CBC
0AFB
0824
0527
01E7
FD9D
F88B
F47C
F2FB
F3A0
F49F
F4DC
F4B3
F4C2
F4D8
F48F
F43C
F477
F501
F505
F466
F419
F4CD
F5D2
F5E7
F4E6
F400
F426
F4D4
F4EC
F468
F483
F628
F8B9
FAA2
FAF4
FA2E
F990
F9C2
FA5B
FA9D
FA6D
FA47
FA66
FA79
FA40
FA06
FA3E
FACB
FB1B
FAEC
FA9F
FA94
FAA3
FA89
FA89
FAEE
FB39
FAB9
F9F2
FA42
FB90
FB8B
F88F
F4C2
F4B6
FA40
01DF
063F
05D6
03BE
0347
045D
04F1
0462
03EE
0466
050B
04F2
045C
0428
047D
04C2
0492
042B
03EB
03EC
0437
04C5
0520
04AD
03CB
0402
065E
09F4
0CB6
0D91
0D2C
0CA9
0C6B
0C42
0C35
0C79
0CE7
0CFB
0C8C
0C00
0BA5
0B5F
0B2E
0B6E
0C2D
0CB6
0C76
0BE8
0BF8
0CA2
0CE4
0C3D
0B8E
0BEF
0D11
0D7B
0C4B
09E9
06D1
029C
FD06
F761
F3E3
F35E
F465
F4F8
F48E
F40E
F42D
F493
F4AD
F499
F4CC
F523
F501
F44B
F3C8
F432
F53B
F5DB
F585
F4C3
F47C
F4D8
F528
F4E6
F486
F50F
F6E1
F922
FA7C
FA78
F9DA
F9BA
FA58
FB0A
FB31
FAF0
FAD6
FB0F
FB47
FB30
FAF1
FADA
FAF5
FB08
FAFA
FAE6
FAD8
FABD
FA97
FA89
FA8E
FA72
FA46
FA6D
FAE8
FACE
F939
F6F2
F67F
F9B4
FF62
042F
05E8
055D
04AE
04AB
0496
0400
03A4
0430
0505
04F0
03D8
02EB
0318
03F2
045E
03EE
032C
02E0
0368
046E
0502
0450
02BD
020D
03D1
07A7
0B6F
0D5B
0D7B
0D19
0D00
0CF8
0CB7
0C7A
0C6D
0C40
0BC5
0B69
0B98
0C14
0C68
0CA9
0D24
0DA0
0D8A
0CEA
0C78
0C90
0CA5
0C46
0C1D
0CEF
0DE0
0D04
09F5
068E
044B
0216
FDED
F833
F3C5
F2A4
F3B5
F47C
F41D
F3AF
F3FC
F465
F43C
F3F7
F44B
F4E7
F50B
F4CE
F4E1
F552
F583
F542
F504
F4FE
F4BA
F41B
F425
F5E8
F8DA
FB11
FB65
FA97
FA04
FA08
FA47
FABB
FB8F
FC50
FC3A
FB5F
FAC4
FB10
FBB4
FBC4
FB3D
FAE3
FB05
FB21
FADB
FA88
FA79
FA60
FA0C
FA19
FB02
FBD9
FAE0
F7CF
F4D3
F4C4
F876
FDFF
028E
049D
0484
0395
030A
035A
0415
0459
03CC
0311
030C
03D5
04A1
04B3
041D
038A
037F
03F1
0467
0460
03BC
02F9
030D
04B3
079E
0A85
0C33
0C86
0C4B
0C50
0CBC
0D2D
0D43
0CFB
0CAD
0CAA
0CE3
0CF8
0CAE
0C40
0C18
0C40
0C4C
0BF5
0B8E
0B88
0BB4
0B8C
0B2E
0B69
0C72
0D20
0C1C
0991
06EC
04C2
01D7
FD00
F769
F3E1
F3A6
F4F7
F54B
F442
F380
F419
F53D
F5A4
F542
F4EF
F4F2
F4CD
F459
F426
F47E
F4E1
F4DE
F4D1
F520
F55C
F4FA
F4AC
F5DF
F8AE
FB2F
FB8D
FA4F
F9A7
FAA4
FC06
FC33
FB44
FA7F
FA6F
FA8F
FA73
FA56
FA7B
FAB0
FABF
FADB
FB2F
FB71
FB4D
FB08
FB1B
FB4B
FB0A
FAB3
FB49
FC73
FBF8
F87F
F446
F39A
F838
FF2C
03E7
04C6
03CF
0375
03FA
0439
03D3
0372
0386
03BD
03B3
036E
031D
02DC
02E1
0367
0440
04D5
04C9
0469
0433
042B
0423
049B
0687
09E5
0D18
0E5A
0D9E
0C6B
0C09
0C5B
0C97
0C82
0C82
0CC6
0CE3
0C7D
0BF9
0C1A
0CF2
0D9E
0D4A
0C3F
0B9D
0C04
0CD5
0CF3
0C34
0B96
0BD4
0C37
0B5E
0902
0618
032B
FF84
FAAA
F5F6
F39A
F40A
F551
F558
F443
F3BA
F464
F523
F4F1
F453
F456
F4F2
F548
F518
F4F7
F535
F566
F52F
F4E4
F4E8
F4F5
F4AC
F496
F5D0
F870
FB01
FC0E
FBAE
FB11
FAF2
FB1F
FB37
FB39
FB4C
FB78
FBBC
FC0D
FC27
FBA7
FAA2
F9CE
F9BF
FA1D
FA33
FA16
FA7D
FB53
FB70
FA66
F9A4
FAAA
FC6E
FBFA
F837
F429
F43E
F984
0078
04C0
0542
0418
0378
03B7
0417
043F
0462
0481
0445
039C
030D
0339
0421
0519
0563
04DE
0420
03EA
0467
04E7
04A5
03EA
0420
065A
09F1
0CEA
0DDA
0D1F
0C2B
0BF1
0C3E
0C76
0C75
0C6E
0C56
0BE6
0B36
0AEE
0B8B
0CA9
0D49
0CF4
0C3D
0C12
0C8F
0CD5
0C39
0B39
0AEC
0B94
0C2F
0B98
09B4
0715
03CF
FF59
F9DA
F4FE
F2B8
F338
F4A7
F529
F496
F401
F41A
F48C
F4DA
F505
F538
F540
F4DA
F442
F40A
F457
F4C1
F500
F535
F564
F532
F498
F468
F594
F7EF
FA38
FB5F
FB82
FB74
FBB1
FC0F
FC3E
FC21
FBAC
FAFF
FA9E
FB05
FBD8
FC16
FB67
FAA1
FA99
FAF3
FAD7
FA61
FA70
FB0C
FB02
F9D3
F906
FA3E
FC4F
FC02
F86E
F505
F605
FB89
017B
0443
0410
0358
036D
03B9
0396
0379
03E0
0460
045B
0405
03EC
040C
0406
03E4
03ED
0404
03DE
03BA
041A
04B8
049B
03B3
03A5
0617
0A52
0DA2
0E52
0D5C
0CAB
0CAF
0C92
0C1E
0C13
0CBD
0D49
0D03
0C66
0C65
0CF0
0D06
0C33
0B4D
0B50
0C1D
0CC5
0CBE
0C42
0BBF
0B7B
0B95
0BE9
0BE1
0AB2
07D4
033C
FD79
F7D8
F40E
F317
F429
F528
F4AC
F368
F30D
F408
F510
F50F
F48A
F491
F521
F562
F510
F4BE
F4C4
F4CD
F49E
F4A2
F533
F5C1
F588
F4F7
F578
F796
FA15
FB71
FB8A
FB58
FB6A
FB8C
FB8A
FB8C
FBA4
FB9F
FB79
FB7F
FBC6
FBDE
FB6D
FADE
FACA
FAF7
FAB2
FA20
FA2E
FAF4
FB41
FA88
FA19
FB3A
FCA0
FB92
F7E9
F563
F7B4
FDF4
036B
04DA
0393
02D0
0395
047A
0473
040F
03FC
03DA
0319
0228
01F6
02A6
0373
03C8
03C7
03B7
0395
0386
03E7
0480
0467
0375
032E
0541
0939
0CA2
0DA6
0CDA
0C20
0C4D
0CB3
0C97
0C3B
0C26
0C41
0C37
0C2C
0C6E
0CC6
0CC1
0C76
0C6D
0CC1
0CF0
0CA5
0C3E
0C38
0C70
0C64
0C19
0C17
0C55
0BA1
08A3
0344
FCE7
F769
F41B
F339
F3DE
F49B
F493
F40A
F3C8
F402
F43E
F431
F443
F4E6
F5C1
F610
F5B7
F564
F57E
F5A6
F583
F563
F58C
F584
F4CA
F404
F49D
F6F8
F9B4
FB1A
FAF3
FA7B
FAA9
FB41
FB9C
FBA4
FB9B
FB8A
FB66
FB5F
FB8F
FBA5
FB61
FB0A
FB0B
FB36
FB05
FA8A
FA73
FAEA
FB21
FA99
FA43
FB3B
FC89
FBCD
F8C5
F6BE
F91D
FF0C
0423
0554
03E9
031B
03FB
04E5
0476
036B
0328
03AF
0408
03E6
03CA
03DF
03B5
031F
029F
02AE
0334
03D8
0468
04A7
042F
032F
02F7
04F4
08D0
0C49
0D6E
0C98
0B9F
0BA0
0C2F
0C77
0C57
0C24
0C0D
0C07
0C1A
0C53
0C8A
0C83
0C5C
0C69
0CA0
0C8B
0C0E
0BB3
0BDC
0C11
0BBB
0B35
0B6D
0C4D
0C12
08BF
0242
FAED
F5AA
F3BC
F424
F4F0
F4ED
F444
F3D0
F40D
F4AF
F519
F513
F4CC
F469
F3FF
F3E8
F487
F585
F5E0
F52B
F45B
F4A4
F5BE
F617
F4FB
F3E5
F4DA
F7C2
FA63
FB15
FA86
FA57
FAEC
FB68
FB4A
FAFF
FAF4
FAF7
FAD2
FAE0
FB7C
FC3C
FC65
FBEA
FB68
FB1E
FAC2
FA74
FAD4
FBC4
FC06
FAF8
F9D3
FA22
FB45
FB00
F8DC
F7AD
FA71
0047
0502
05E1
0457
0383
0449
0518
04CB
040E
03E8
042F
0419
038F
0335
0364
03D0
0425
045A
044D
03D3
0353
0395
047E
04CA
03D8
0319
04AB
0899
0C78
0E05
0D6F
0C8B
0C6D
0C99
0C6F
0C3B
0C76
0CD2
0CB5
0C31
0BD7
0BD0
0BD7
0BEC
0C47
0CB6
0CA2
0BFF
0B9E
0C0D
0C99
0C35
0B3A
0B39
0C80
0CB4
08F7
0153
F931
F431
F313
F3DF
F46C
F436
F3F1
F415
F45D
F471
F46F
F4A2
F4F9
F515
F4D0
F476
F462
F47E
F45B
F3E3
F3A9
F435
F518
F553
F4BD
F47A
F5A5
F7DA
F99A
FA14
F9F7
FA4F
FB1C
FB89
FB41
FAE3
FB03
FB66
FB90
FB7F
FB6C
FB43
FAD2
FA60
FA71
FAF9
FB51
FB13
FAA5
FAA1
FB0A
FB79
FBD8
FC3D
FC33
FB1D
F996
F992
FC46
006B
036C
042A
03CB
03D7
0453
044E
039F
0324
0368
03E8
040A
03FC
0419
0427
03C8
034F
035B
03E4
044E
0468
048A
04A6
0401
0295
0215
0469
090F
0D1A
0E4C
0D56
0C73
0C8D
0CD5
0CAB
0C97
0D18
0D8C
0D1A
0C1E
0BC1
0C41
0CAA
0C5C
0BEE
0C09
0C4D
0C20
0BD5
0C15
0C75
0BE9
0AC5
0ADD
0CBE
0DAA
09FD
01B0
F92B
F4CA
F494
F545
F4BD
F3ED
F469
F5C4
F648
F57B
F4A6
F4E8
F5C8
F62C
F5EC
F5B8
F5D9
F5E5
F5A2
F571
F5AF
F614
F61C
F5A9
F50C
F48B
F45E
F4FD
F6D8
F997
FBF8
FCF4
FCC6
FC86
FCCB
FD28
FD03
FC79
FC28
FC52
FC9C
FC98
FC52
FC23
FC3A
FC7D
FCB8
FCC4
FC9B
FC64
FC64
FCA5
FCD0
FC96
FC2E
FC23
FC8E
FCCF
FC67
FBF6
FCE1
FFB3
0330
055F
0577
0475
03D5
0410
048D
04AD
0478
0445
0425
03EA
03A2
03A3
0410
0491
04B0
045E
03F1
03B7
03B9
03EF
045D
04ED
0543
0525
0508
05E5
082B
0B00
0CE9
0D38
0C92
0C03
0BE9
0C07
0C37
0C9A
0D12
0D23
0CA0
0C1A
0C2B
0C8D
0C81
0BFA
0BBC
0C1A
0C68
0C15
0BC2
0C54
0D45
0D16
0BA7
0AF5
0C51
0D7D
0A66
021F
F8D9
F3BF
F3BC
F568
F59B
F485
F409
F4A3
F52A
F505
F4FA
F5A1
F644
F601
F53D
F4FE
F579
F60D
F671
F6E0
F736
F6CF
F590
F46D
F43E
F491
F47D
F45F
F5A9
F8A5
FB81
FC5F
FB95
FB10
FBCD
FCFE
FD7C
FD2F
FCB0
FC50
FC07
FBFE
FC68
FCF0
FCF9
FC93
FC6B
FC9F
FC6A
FB7D
FACE
FB49
FC4C
FC84
FBEF
FBE8
FCF0
FD9D
FCAA
FB52
FC49
0029
044D
05D1
04BD
035E
0336
03D0
043D
0466
0487
046C
03D5
0340
036A
0420
045B
03B8
031D
0375
0466
04E2
04A7
0466
0491
04BE
0461
03AB
037D
04A0
0722
0A41
0CD9
0E09
0DCC
0CF9
0C7D
0C7F
0C7B
0C30
0BF6
0C11
0C3C
0C22
0BE5
0BC8
0BC1
0BB4
0BCE
0C2B
0C5F
0BF3
0B43
0B3B
0BDB
0BE2
0AB9
09FB
0B86
0DE4
0C93
050F
FA97
F361
F24C
F4AA
F635
F5B7
F4F1
F52F
F5B4
F588
F51B
F54B
F5DA
F5E5
F55A
F4E8
F4D8
F4D6
F4CD
F50E
F589
F5A4
F534
F4F5
F579
F605
F56B
F40C
F3DF
F611
F969
FBB2
FC2C
FBCC
FB95
FBAC
FBDA
FC13
FC3E
FC12
FB93
FB5A
FBDE
FCB5
FD0D
FCD5
FCBE
FCF7
FCE4
FC50
FC08
FC9A
FD32
FCB5
FB86
FB15
FBBB
FC2B
FB80
FAFA
FC9F
0065
03E1
050F
0462
0396
0365
0366
0360
039F
0405
03E6
0324
02B3
0365
04B2
0544
04B0
03F6
0417
04D5
0532
04D6
0453
0456
04F0
0593
0591
04D7
0469
05A9
08BC
0BF7
0D6B
0CFF
0C6D
0D00
0E01
0DEB
0CAA
0BB9
0BFF
0CA9
0C9B
0BFE
0BB4
0BE4
0C0A
0BF8
0BEB
0BC4
0B1B
0A4B
0A6C
0BB1
0C9E
0BF3
0AE1
0B91
0D54
0C1B
052B
FB3D
F42F
F2E1
F4CB
F5CF
F4D0
F3AF
F3CE
F470
F473
F421
F463
F526
F597
F578
F543
F52D
F4F1
F490
F479
F4BF
F4DA
F471
F3FD
F416
F46D
F432
F387
F3C3
F5DB
F90A
FB98
FCA4
FC99
FC3A
FBEC
FBD6
FC15
FC92
FCF6
FCF9
FCAB
FC4E
FC11
FC01
FC22
FC4B
FC0F
FB3B
FA5D
FA49
FAED
FB49
FAEB
FABC
FBB3
FD34
FDA9
FCC0
FC2F
FDBA
00EB
0387
0421
0379
0320
038E
041F
045F
0480
04B8
04D4
04A0
0443
0408
03FA
03E5
03AF
038E
03D1
0485
054F
05B1
057E
0525
0546
05C0
0582
03F7
0279
0367
0755
0BE7
0E2A
0DB5
0CA2
0CB1
0D66
0D5D
0C7E
0BF0
0C32
0C7C
0C2B
0BC3
0BF2
0C69
0C7B
0C41
0C41
0C4B
0BBD
0AD5
0AAF
0B8D
0C15
0B3C
0A3A
0B07
0CD8
0BD4
0572
FC29
F54F
F397
F4DB
F572
F446
F2EB
F2C0
F355
F3AC
F3B7
F3F0
F438
F407
F37B
F34B
F3C7
F471
F4CC
F4F9
F553
F5C8
F5F6
F5C3
F57C
F555
F524
F4D0
F4CC
F5C4
F7C4
F9F9
FB56
FB78
FAE5
FA89
FAE1
FBA4
FC37
FC65
FC66
FC4F
FBEF
FB56
FB1B
FBAA
FC81
FC97
FBB3
FADD
FB0E
FBD6
FBF3
FB2B
FAB7
FB6E
FC6C
FC42
FB36
FB3F
FDAB
0168
0422
04B9
0418
03C3
0436
04D7
050B
04CA
0470
0454
048C
04D1
04BB
0445
03E9
0404
0462
0497
04A4
04D0
04FD
04A1
03B4
0325
03BE
04D2
0503
0468
04ED
07DE
0BD8
0E1C
0DAB
0C25
0B85
0BF1
0C4E
0C25
0C0E
0C57
0C74
0C06
0B92
0BA5
0BE7
0BCB
0B9A
0BE5
0C54
0BF0
0AC7
0A2B
0AD6
0B9B
0B0C
09E1
0A2A
0BD0
0B71
0614
FD45
F5F8
F364
F427
F4D0
F404
F31B
F357
F41C
F43A
F3C6
F3B2
F430
F484
F44D
F415
F44D
F490
F459
F405
F470
F5A4
F698
F67B
F5C4
F57E
F5D5
F5F2
F563
F502
F601
F852
FA8E
FB79
FB44
FB10
FB6D
FBD4
FBAC
FB49
FB77
FC3F
FCCB
FC8B
FBF0
FBAD
FBAC
FB58
FAB9
FAA0
FB70
FC4C
FC22
FB33
FAC3
FB40
FB9E
FB12
FA9E
FC0B
FF7F
02FC
0489
0438
039A
03BE
0459
04C6
04F3
0505
04D0
0438
03AA
03A5
0409
0460
049B
050B
05A0
05C8
0549
04B7
04AD
04DF
049E
0408
03EB
0446
0417
0318
02E7
0546
098D
0CF0
0D7E
0C19
0AFF
0B18
0B83
0B6B
0B1E
0B23
0B41
0B14
0AE0
0B0B
0B4D
0B29
0AEA
0B51
0C3D
0CA1
0C10
0B81
0BD0
0C38
0B7B
0A46
0AB6
0CCE
0CF5
0799
FDEA
F54B
F1DB
F2BC
F434
F459
F432
F4E9
F5B6
F548
F3F8
F34B
F3C0
F460
F467
F445
F498
F500
F4B9
F3EF
F39E
F420
F496
F42A
F352
F335
F406
F4C7
F4CD
F4D9
F633
F8FA
FBCD
FD39
FD24
FC94
FC53
FC34
FBCD
FB58
FB72
FC22
FCAE
FC8F
FC1D
FC07
FC50
FC53
FBC5
FB31
FB21
FB4F
FB2A
FAFA
FB8E
FCBC
FD1E
FBFA
FACC
FBF1
FFB5
03A7
053E
0484
038E
03AF
043E
041F
037D
033D
0383
03A6
036A
036C
041D
04FE
0540
04BE
0410
03B4
03AB
03C8
03FD
0428
041C
0400
043F
04C8
04E6
0456
0417
057B
0867
0B2D
0C4C
0BF4
0B7B
0BA3
0C00
0BFF
0BBE
0BB0
0BE4
0C1F
0C45
0C42
0BE0
0B2F
0AC1
0B0E
0BB0
0BDE
0B92
0B9B
0C32
0C43
0AF1
0966
09BC
0BBB
0BEE
0737
FEC2
F740
F428
F4A4
F57C
F4FF
F41D
F423
F4C4
F4D7
F426
F38D
F3A5
F41C
F46A
F48A
F4AE
F4C4
F48A
F40B
F3AF
F3CB
F447
F4CA
F51B
F544
F553
F542
F51D
F52D
F5E0
F76A
F964
FAF2
FB71
FB21
FAD7
FB0A
FB63
FB6A
FB3D
FB5C
FBD4
FC19
FBBD
FB08
FA96
FA94
FABF
FAF6
FB60
FBEC
FC29
FBEB
FBA2
FBC1
FC18
FC52
FCCE
FE69
0127
03AB
047E
03B6
02D6
0304
03E9
0485
048B
0470
047C
0468
0400
039A
03B1
0440
04BC
04AB
041D
0392
037F
03E3
0445
0424
038C
0331
039E
045A
0457
0371
0302
047B
079A
0A8E
0BD9
0BAA
0B2E
0B08
0AF1
0AAD
0A97
0B0F
0BD0
0C41
0C26
0BB4
0B2A
0ABE
0ABD
0B51
0C15
0C5F
0C11
0BB7
0BA0
0B3F
0A1F
0923
09D3
0BF0
0C88
0893
0084
F864
F415
F3D9
F4EE
F501
F44D
F452
F562
F644
F5EA
F4BE
F400
F442
F4FA
F55C
F53B
F4FB
F4E4
F4DA
F4B1
F48B
F4AB
F50A
F548
F51B
F49F
F42F
F408
F427
F496
F58C
F72A
F915
FA97
FB3A
FB34
FB17
FB26
FB2C
FAE3
FA74
FA58
FACD
FB78
FBC7
FB98
FB5E
FB8C
FBEB
FBD4
FB17
FA60
FA81
FB6D
FC35
FC23
FB8A
FB35
FB52
FB85
FBFE
FDBA
0124
04E3
06C3
0605
0435
0361
03E5
047A
042C
037A
035F
03E0
043B
0410
03C7
03CC
0408
0441
0480
04B9
0474
036C
0256
0261
03A0
04A7
0438
02ED
0278
0366
046A
0446
03AE
048B
077A
0ADB
0C9D
0C75
0BC0
0B9C
0BD6
0BC5
0B6D
0B5D
0BB9
0BF5
0B9C
0AE9
0A82
0AC1
0B7A
0C3B
0C90
0C32
0B50
0A9A
0AA0
0B0A
0AD3
09AE
08CB
0994
0B74
0B8C
0756
FF84
F7C7
F37B
F2E7
F3D6
F464
F485
F4F8
F598
F57F
F47B
F391
F3C8
F4D9
F58A
F530
F462
F41C
F48C
F517
F54E
F56E
F5D2
F63E
F61E
F560
F4B7
F4CD
F563
F58A
F4E4
F454
F536
F7CB
FAB4
FC33
FBEC
FB23
FB34
FC19
FCB2
FC53
FB89
FB35
FB59
FB40
FAC4
FAAA
FB82
FC97
FCB1
FBBD
FB04
FB79
FC70
FC99
FBE9
FB9C
FC3E
FCB1
FBF2
FB45
FD4C
028F
07F0
0996
0704
0375
021F
02FE
03CC
034C
027E
02C3
03E7
04A8
0477
03E2
0386
0364
0362
03B6
0461
04CA
0472
03D5
03EE
04BE
0510
0417
02B3
0261
0334
03AB
02D7
01E6
02E6
0646
0A31
0C86
0CD2
0C2C
0B9C
0B4B
0B13
0B14
0B81
0C19
0C5A
0C0C
0B72
0AEF
0AB4
0AC1
0AEE
0AEB
0A73
09C5
0994
0A3E
0B17
0B10
0A1F
0995
0A8E
0C1B
0B99
072E
FFD1
F8A1
F43C
F2F1
F34B
F3E2
F446
F491
F4B9
F499
F454
F44F
F4B7
F53F
F57F
F56E
F560
F593
F5E2
F5FB
F5B9
F54A
F4E7
F49A
F44E
F419
F44F
F518
F5EE
F5DE
F492
F328
F38A
F68A
FAB9
FD7D
FD89
FBFE
FAFE
FB58
FC0F
FBFF
FB58
FB18
FB84
FBE3
FBA6
FB38
FB33
FB55
FAEF
FA30
FA36
FB83
FD0B
FD6D
FCD1
FCA2
FD57
FD91
FC3D
FAF2
FCCE
0283
0890
0A73
0783
0385
0255
03D9
04FC
03F3
0236
021B
03AB
04D5
044C
02FC
027C
0304
038F
0396
0398
0400
045F
0437
03F7
0469
055F
05B3
04D1
0393
032E
039A
03CD
0370
03A2
0594
08CB
0B68
0C1D
0B64
0AA5
0AA4
0B0F
0B4F
0B54
0B5B
0B63
0B2E
0AB3
0A55
0A79
0B07
0B70
0B34
0A60
099D
0998
0A56
0B1A
0B30
0ABE
0AA2
0B43
0B9B
09CE
04F2
FE39
F82B
F4B3
F3E4
F46E
F4EF
F4C9
F424
F38E
F39B
F481
F5CB
F69A
F66E
F5A5
F500
F4D3
F4CA
F494
F46F
F4C5
F56D
F5AD
F50F
F3F0
F31B
F30D
F3AD
F480
F4F4
F4B3
F41C
F452
F654
F9AC
FC6A
FCFE
FBEB
FB19
FB7C
FC1F
FBC7
FAD3
FAA3
FB85
FC47
FC0B
FB9A
FC1E
FD23
FD17
FBB2
FA9D
FB22
FC3B
FC1B
FAF9
FAD8
FC5E
FD70
FC39
FA97
FC96
032D
0A03
0BC5
080D
0391
0299
04A1
0613
0514
0334
02B2
038E
0420
03B0
032D
037F
043A
047A
0450
047D
050D
0516
041A
0304
031C
044A
050E
0460
0301
0273
02FF
0388
0352
033C
04BA
07D9
0AF6
0C7A
0C68
0BE8
0BB4
0B8A
0B09
0A85
0A8F
0B1C
0B87
0B66
0AFC
0AD1
0B14
0B73
0B88
0B3F
0AE7
0AE1
0B2B
0B47
0ABC
09D5
0998
0A7E
0B42
0992
0461
FD51
F76E
F489
F419
F477
F49E
F483
F446
F3D8
F356
F32B
F37B
F3D7
F3D4
F3B3
F3FE
F4A8
F509
F4C0
F43A
F419
F468
F4AF
F4A3
F476
F46F
F49D
F4FA
F581
F5F1
F5CE
F51C
F4D3
F60D
F8A5
FB1E
FC2D
FC09
FBDE
FC39
FC96
FC7C
FC5A
FCC5
FD5A
FD17
FBDC
FACF
FAE9
FBA3
FBB6
FAED
FA64
FAE0
FBA9
FBB4
FB58
FBE0
FD44
FD9F
FBD6
FA29
FC7E
03A0
0B35
0DA8
09E8
0458
01E3
0324
04F8
04F0
03B4
0319
035F
0367
02E2
02CD
03B6
04A9
0481
03A6
037B
044F
04D8
0410
02CC
02AC
03F0
0531
0538
0467
03E3
03F9
03F5
0378
0352
04A3
0775
0A80
0C54
0C83
0BBF
0B0B
0ADD
0AED
0AC9
0A81
0A9B
0B54
0C29
0C69
0C12
0BC7
0BD6
0BBA
0AED
09FE
0A07
0B0F
0BAC
0AC5
0947
092C
0AC5
0BC1
0973
03BF
FD3B
F885
F619
F4D4
F3DD
F345
F33B
F375
F3A3
F3F2
F497
F532
F51F
F46A
F3EB
F442
F507
F558
F4FC
F496
F4AB
F4FE
F508
F4CB
F4BF
F515
F56C
F56C
F542
F54B
F578
F57E
F591
F67F
F8A6
FB22
FC71
FBFF
FABB
FA04
FA4D
FB13
FBD3
FC8F
FD45
FD81
FCE7
FBF0
FB7E
FBC5
FC05
FB9F
FAEE
FAA9
FAC7
FAB5
FA87
FB19
FC8C
FD68
FC72
FB29
FD06
0360
0AC9
0DDB
0AC3
0525
0207
02B5
046C
047C
033D
0297
0307
0353
02CC
0264
0315
0432
0448
033D
0297
036C
04E6
0568
04A8
03E6
0412
0499
0456
0332
023E
0238
02AD
02D0
02D6
03E9
06A0
09F6
0C22
0C5B
0B8D
0B36
0BCB
0C7D
0C6B
0BB3
0B1D
0AFE
0AE6
0A75
0A06
0A2C
0AC2
0AFA
0A88
0A32
0ACC
0BE7
0C21
0AFE
09DF
0A7B
0C67
0CE0
097D
02D3
FC02
F7BB
F621
F597
F4FD
F488
F495
F4AC
F42A
F369
F372
F488
F59B
F5A0
F4E6
F49A
F520
F5A3
F55B
F4B0
F497
F529
F585
F51A
F457
F3EA
F3E3
F407
F479
F563
F634
F609
F514
F4E7
F6AE
F987
FB68
FB89
FB29
FB9E
FC8F
FCC6
FC22
FBC5
FC52
FD04
FCE5
FC37
FBEE
FC2B
FC12
FB42
FA7B
FA7D
FAEC
FB0C
FB18
FBE1
FD1E
FD4E
FBE2
FAD4
FD0D
02E6
0910
0B86
095C
054D
02B3
028D
037F
03FE
03D3
03A6
03B5
0392
02FB
0274
02A7
0373
03FF
03D5
0370
0380
03EA
0402
03A0
0382
0439
0520
04FD
03AB
0273
027D
0365
03F0
03E7
0482
06C9
0A12
0C81
0CF5
0C0F
0B3E
0B35
0B86
0B83
0B16
0AB9
0AD4
0B5A
0BDF
0C0E
0BF6
0BD3
0BAE
0B5B
0ADB
0A80
0A89
0ABA
0AB3
0A8C
0ACA
0B65
0B2D
08B3
03EB
FE82
FA5E
F801
F6A5
F592
F4D0
F49C
F4B7
F4A6
F457
F427
F43F
F448
F3EE
F377
F37C
F42A
F4FC
F53F
F4C7
F405
F39D
F3E0
F495
F531
F551
F517
F4FB
F545
F5A6
F583
F4BD
F424
F4E3
F73F
FA11
FBC7
FBE5
FB65
FB7A
FC33
FCA2
FC43
FBC0
FC00
FCDE
FD59
FCF9
FC60
FC47
FC7E
FC6C
FC14
FC03
FC50
FC65
FBF4
FB7E
FB61
FB0E
FA1D
F9FD
FD1B
03A6
0A16
0C34
0962
050E
02D0
0304
0399
0340
02A9
02D9
0386
03BF
0365
0326
0353
038E
0389
0376
038C
03A0
036E
0313
02ED
031F
0374
03AA
03A2
0358
02ED
02BE
0305
0354
02FB
023B
028A
0503
08CC
0BAE
0C66
0BC4
0B65
0BC1
0C00
0B86
0AD0
0AAE
0B22
0B89
0B7B
0B1C
0AB4
0A77
0AA1
0B45
0BFF
0C2D
0BB5
0B43
0B85
0C48
0CC5
0CB5
0C88
0C4D
0AF1
0746
01B6
FC5E
F923
F7F7
F747
F5F8
F47F
F3F8
F48B
F529
F4EB
F429
F3F8
F4AE
F575
F557
F463
F38C
F389
F429
F4C8
F509
F4F3
F492
F3FB
F394
F3DC
F4BD
F572
F55F
F4D5
F497
F4CF
F4EF
F4AB
F4A2
F5BB
F7F9
FA54
FBC6
FC38
FC3E
FC46
FC46
FC1C
FBEA
FBF2
FC54
FCE3
FD42
FD30
FCC4
FC44
FBCF
FB63
FB2E
FB7C
FC38
FCB5
FC65
FBBF
FBCD
FC9A
FCC5
FB7C
FA91
FD26
03B8
0A7C
0CD7
0A15
05D4
03C3
0411
0473
0397
0261
020E
0279
02CA
02DC
031A
0383
03AB
038B
037F
0389
033A
0288
0228
02A4
038C
03F9
03BF
037B
0387
0392
036D
0385
03FF
041E
034A
0260
0313
05D7
0927
0B1E
0B64
0B15
0B2B
0B88
0BA0
0B5A
0AF9
0AB1
0A9B
0AD0
0B26
0B34
0AF0
0AF3
0B9D
0C4C
0C0D
0B0B
0A87
0B20
0BCB
0B50
0A53
0AB0
0C90
0D3A
09E8
0337
FCCB
F973
F89F
F7E5
F62D
F488
F430
F4C5
F4FB
F462
F3D5
F423
F502
F57D
F51B
F447
F3C4
F3F6
F4AF
F56E
F5B4
F540
F43F
F33B
F2CA
F30E
F39E
F40F
F476
F522
F5E9
F614
F547
F43A
F439
F5D9
F856
FA64
FB63
FBAF
FBDC
FC11
FC2A
FC1E
FC00
FBD9
FBB6
FBB6
FBE9
FC2F
FC62
FC7D
FC7B
FC46
FBFC
FC09
FCAE
FD70
FD7E
FCCE
FC54
FC92
FC87
FB2C
F9E5
FC03
02BE
0A9E
0E45
0BD9
06AA
0355
0333
0438
045F
03C8
0377
0392
039E
038D
0399
0385
0303
0280
02BA
0383
03D0
0330
0288
02CD
0390
03A9
02F9
0296
0309
0389
036D
0357
0405
04BE
0439
02DD
02DD
058F
0991
0C3E
0C99
0BDE
0B7B
0B7D
0B59
0B27
0B53
0BAB
0BA2
0B40
0B0D
0B28
0B26
0AE3
0AD4
0B3A
0BA2
0B96
0B67
0B9A
0BCB
0B10
09A8
0932
0A62
0B4B
0918
0382
FD75
F9F0
F8F6
F83D
F65A
F44A
F3B9
F4AB
F594
F567
F4B5
F4A0
F54B
F5CA
F55A
F449
F391
F3C0
F47A
F4ED
F4B8
F434
F3F7
F445
F4E2
F55D
F56C
F520
F4D1
F4D3
F51F
F555
F51E
F4A9
F4A0
F5A2
F79C
F9C4
FB36
FB9A
FB42
FAD1
FABF
FB0A
FB4F
FB3F
FB02
FB0E
FB9A
FC6C
FD30
FDAF
FDB3
FD0E
FC09
FB72
FBC9
FC7C
FC7B
FBC3
FB9E
FCB2
FD85
FC51
FA47
FB4A
015E
0948
0D53
0B43
0665
0363
036A
043E
0412
0375
0378
03C3
038B
032E
038E
0460
0476
0396
02DE
0317
039E
037E
02F7
0305
03BC
042A
03E6
03A1
03DB
03FF
0397
0366
0439
0551
0528
03DC
0382
05A0
0919
0B73
0BB7
0B1A
0AFA
0B48
0B54
0B1C
0B0B
0B0F
0AE2
0AC4
0B1D
0B9D
0B97
0B23
0B18
0BA4
0BCC
0ADF
09D0
0A14
0B58
0BBD
0A9A
09A7
0A61
0B4F
0969
040C
FE18
FAA3
F9A2
F8B5
F694
F46F
F3DC
F49C
F530
F4E6
F466
F461
F4AF
F4D6
F4C7
F4B3
F492
F444
F403
F438
F4DB
F54E
F519
F498
F490
F528
F59D
F532
F42B
F392
F408
F50F
F59D
F55A
F510
F5DE
F7FA
FA77
FC20
FC7C
FBF9
FB62
FB42
FBA4
FC28
FC61
FC38
FBF9
FBFB
FC47
FC9A
FCA8
FC4F
FBB2
FB2F
FB2F
FBC1
FC5C
FC51
FBB2
FB6A
FBFA
FC7A
FBC8
FAD1
FC7B
024C
09B0
0DC6
0C32
0769
03DC
036E
0476
04AE
03CD
02F4
02C8
02FF
0337
035A
0356
0325
0318
0375
03E4
03BF
0316
02D0
0363
03FC
039D
02BD
02C7
03F5
04D9
047A
03BE
03D6
0439
0393
024C
02A2
05BD
09C9
0BEF
0BA1
0AC8
0AF7
0BC3
0C29
0C35
0C65
0C67
0BAE
0AB7
0A85
0B0B
0B31
0A93
0A2C
0AB5
0B55
0AE1
09D8
09CA
0ACE
0B2F
0A38
09A8
0B01
0C6F
0A5B
0422
FD67
F9F6
F988
F8D7
F637
F36C
F2C2
F3E1
F4B2
F45F
F405
F495
F57A
F5A9
F529
F4D3
F505
F54A
F542
F536
F584
F5F1
F5F1
F56F
F4E4
F4AD
F4BB
F4DE
F519
F578
F5D2
F5E0
F589
F50A
F4DC
F57C
F720
F979
FBAA
FCB5
FC42
FB05
FA34
FA72
FB51
FBF1
FBEF
FBA3
FB83
FB9A
FBB8
FBCB
FBE2
FBEB
FBCA
FBA6
FBD8
FC57
FC97
FC53
FC18
FC7A
FCE8
FC50
FB47
FC70
01A3
08E1
0D65
0C4D
079E
03F5
03B0
0530
05B4
048F
0312
025A
0265
02CB
035D
03CE
03B2
0313
02A3
02DE
035D
036D
031F
031A
037C
03AA
036C
0360
03E3
044A
03F3
036A
03AA
046A
045D
0350
0307
0530
08FC
0BC2
0C1C
0B46
0B27
0BE4
0C47
0BC4
0B13
0AF0
0B32
0B4F
0B23
0AE8
0AC8
0ACD
0AF8
0B1E
0AE4
0A4E
0A1F
0AF3
0C0D
0BF3
0A8F
09BB
0AC0
0C08
0A7B
0535
FED6
FAA3
F917
F814
F5FF
F39E
F2A5
F367
F4A6
F53C
F515
F4BE
F4A1
F4CE
F50F
F4FF
F46D
F3BE
F3AC
F474
F56A
F5B3
F540
F4C9
F4CF
F50A
F500
F4CB
F4DC
F53F
F591
F590
F566
F553
F577
F60E
F772
F990
FB85
FC3D
FB9D
FAC4
FACD
FBA0
FC3F
FC2E
FBFB
FC50
FCF1
FD1A
FCA1
FC2C
FC33
FC59
FC0F
FB8D
FB98
FC3D
FC99
FC20
FB99
FC01
FCCC
FC7B
FB33
FBAE
0057
07C1
0D25
0D01
0894
0442
02F9
0406
0512
0501
0453
03B9
0360
0355
03A8
0415
042A
03ED
03DE
042C
0448
03BF
030A
0301
039C
0403
03E3
03D8
042B
0425
0344
0264
02B5
03DB
0445
0385
033B
050A
0843
0AAC
0B48
0B2C
0B6F
0BA7
0B24
0A8E
0B02
0C26
0C6A
0B3D
09DC
0995
0A1C
0A4E
09FE
09F5
0A65
0A8E
0A2D
0A24
0AF3
0BA5
0B44
0A96
0B13
0C35
0B53
06D0
0074
FBA1
F992
F88F
F6CE
F4CE
F41F
F4DB
F57E
F4FC
F3E4
F34B
F376
F3F0
F456
F494
F499
F44D
F3F1
F401
F494
F52B
F555
F539
F537
F549
F51A
F4AC
F460
F475
F4BD
F4E4
F4BE
F45E
F413
F47C
F630
F8FC
FB9A
FCA6
FC1B
FB63
FBB8
FCB5
FD07
FC3D
FB55
FB5E
FC22
FC9D
FC71
FC33
FC59
FC78
FC0B
FB7D
FBBA
FCBF
FD5D
FCD3
FBF9
FC0F
FCBC
FC56
FA9F
FA39
FE1F
05AF
0C4C
0DA6
09F3
054A
0327
0384
0442
0436
03E2
03E3
03EC
0394
0339
0379
0428
0483
0447
040A
0448
04B1
04AD
0443
03F2
03F4
0416
043C
0488
04E4
04D6
041E
0338
02EF
034E
037D
02D8
020B
02A2
056C
0967
0C6E
0D10
0BC2
0A5A
0A42
0B3E
0BFF
0BCC
0B19
0AAA
0A8D
0A5F
0A29
0A5C
0AF3
0B36
0AB9
0A2E
0A8B
0B97
0C16
0B73
0A89
0A55
0A9D
0A9E
0A75
0AD5
0B3F
09BE
0525
FF0E
FA85
F8C5
F82F
F6C9
F4C5
F3C9
F466
F55E
F56D
F4C1
F447
F432
F3F4
F361
F31B
F3A3
F48A
F4F4
F4A8
F428
F3F1
F405
F429
F44C
F486
F4EC
F56E
F5C5
F59B
F4F3
F45A
F476
F537
F5B9
F54D
F48A
F4E0
F6EE
F9A5
FB60
FB9B
FB30
FB0E
FB43
FB5E
FB58
FB94
FC2C
FCA8
FC9D
FC49
FC3E
FCA7
FD15
FD13
FCA6
FC2C
FBED
FBE1
FBD8
FBB5
FB97
FBC2
FC51
FCD9
FC9D
FB94
FB2A
FD7F
032D
09D7
0D9D
0C7F
083E
0489
0379
0434
04D2
04B5
048D
04B3
048C
03AD
02CD
02E2
03C6
046E
046D
0468
04DB
0534
04B6
03C2
0369
03DD
042C
03BC
033D
039A
0476
0497
03BC
0305
033E
03B0
036D
0318
044A
0746
0A3C
0B5D
0AE2
0A6C
0AD1
0B6C
0B8F
0B8F
0BF0
0C50
0C02
0B4C
0B22
0BA0
0BB9
0AC7
09AB
09B3
0AC6
0B81
0B36
0AD4
0B56
0C1E
0BCF
0A8A
0A1D
0B7C
0CDD
0B55
062D
FFD6
FB4A
F925
F7D1
F611
F468
F3E0
F44E
F491
F42C
F3DD
F45E
F539
F554
F475
F393
F39C
F457
F4D1
F49B
F43B
F451
F4D1
F525
F4F5
F476
F426
F451
F4D2
F533
F513
F49A
F473
F50C
F5EC
F616
F54A
F4AD
F5AB
F84B
FAF2
FC0D
FB9F
FAE9
FAD8
FB3D
FB75
FB54
FB2D
FB3C
FB6B
FB97
FBCC
FC10
FC40
FC36
FBFE
FBBC
FB8C
FB81
FBA3
FBD4
FBE7
FBFE
FC69
FCFF
FCDF
FB9A
FA92
FC6C
0241
0993
0DF3
0D1E
090B
0589
0461
0470
040C
0339
030D
03C6
0468
042F
0387
034A
0390
03C2
03A3
0394
03D3
0409
03D5
0370
035F
03B1
03E6
03BA
0390
03E3
0479
0494
03F4
0337
0301
031F
02F0
02A3
0368
060D
09A4
0C18
0C49
0B2D
0A90
0B10
0BCF
0BF9
0BD5
0C15
0CA5
0CD7
0C72
0BFA
0BD0
0B99
0B04
0A90
0AF8
0BF2
0C56
0BA9
0AC0
0A77
0A75
09F8
0964
09E9
0B59
0B73
082E
0263
FD1E
FA4F
F914
F7A7
F5E1
F4F2
F53D
F5A5
F52E
F447
F3E8
F41F
F42F
F3E6
F3D6
F433
F453
F3CD
F35B
F3E1
F503
F588
F509
F472
F4A7
F554
F597
F55A
F54C
F5A8
F5D8
F587
F53B
F564
F57C
F4E8
F452
F535
F7DD
FAB3
FBF0
FB91
FB09
FB4B
FBE2
FC13
FBF2
FBFD
FC2D
FC22
FBF6
FC1F
FC99
FCC6
FC55
FBC4
FBB7
FC1B
FC63
FC5E
FC50
FC4B
FC1B
FBEE
FC53
FD24
FD45
FC59
FC3A
FF82
0614
0C16
0D5A
09A2
04C3
0282
0327
045A
047A
03F9
03DE
042D
0441
03FD
03E2
0423
044A
03F5
0379
0377
0404
0494
04A8
0442
03AE
0329
02DA
02E6
0348
03B2
03C5
0376
0321
0319
0332
0303
02BC
035C
05B6
0935
0C0A
0CD8
0C0D
0B41
0B58
0BAD
0B53
0A93
0A82
0B5F
0C1E
0BE5
0B2D
0AF3
0B43
0B58
0AEF
0AB2
0B09
0B50
0AE1
0A48
0A85
0B47
0B2B
0A03
0989
0AD6
0C10
0A11
045A
FE0C
FA61
F92D
F7E4
F569
F355
F353
F4AA
F55B
F4C1
F3EF
F3D0
F41E
F447
F456
F47F
F47F
F416
F3C6
F449
F55A
F5D6
F544
F481
F46E
F4C6
F4D1
F4AF
F50B
F5C8
F607
F58E
F54A
F5D3
F640
F55B
F3D3
F3EC
F6AF
FA55
FC4A
FC1A
FB6C
FB8F
FC15
FC05
FB70
FB30
FB9C
FC39
FCA5
FD00
FD52
FD30
FC6A
FB95
FB64
FBC9
FC33
FC68
FC96
FCAF
FC68
FBEC
FBE6
FC64
FC5C
FB39
FAA5
FD75
041E
0B15
0DCB
0B3E
06BC
0421
0423
04BC
0451
035F
0320
03AA
0416
0402
03F4
0457
04BD
0482
03BF
0326
0322
0372
03A6
03B0
03C1
03D6
03BF
0389
038E
03F2
0451
043C
03E1
03D6
043A
0467
03E4
0371
047E
0766
0A98
0C1D
0BBC
0B06
0B38
0BD3
0BB3
0AE0
0A78
0AF8
0B84
0B4A
0ACD
0B0C
0BC9
0BBE
0A9A
09A6
09F3
0ACC
0AD8
0A39
0A44
0B4B
0BDE
0AF8
09CB
0A21
0B5C
0A99
063C
002A
FB8E
F950
F7E2
F611
F487
F443
F4CE
F4EC
F473
F45A
F4FF
F582
F533
F4AB
F4CF
F55F
F56A
F4DC
F4A3
F52F
F5BB
F576
F4C5
F4BA
F58B
F647
F621
F562
F4C8
F494
F4AB
F51C
F5DF
F655
F5CF
F4B3
F473
F5FD
F899
FAAB
FB7A
FBA7
FC00
FC75
FC80
FC16
FBAF
FB97
FBB3
FBE7
FC40
FCAB
FCD4
FC8D
FC0B
FBAA
FB84
FB88
FBCB
FC4F
FCAA
FC5C
FBAE
FB93
FC4C
FCA9
FBA0
FA7A
FC57
029C
0A5F
0E7E
0CA1
0797
0430
045B
05F9
0631
04BB
0375
0386
0417
03D8
02E0
0262
02F5
03DB
0422
03D4
03B6
042D
04C6
04E2
046D
03DF
03A4
03C5
03FD
03FC
03A5
0328
02F6
034D
03C9
03B8
030C
02DE
0481
07E8
0B45
0CA7
0BEC
0ACD
0AD7
0BC2
0C1B
0B53
0A75
0AA9
0BAE
0C37
0BB0
0AE4
0AC8
0B27
0B12
0A53
09B3
09D4
0A65
0ABC
0AC3
0ABF
0AB0
0A7E
0A9D
0B97
0CAB
0BA9
072B
00B5
FB8E
F953
F878
F6B6
F404
F24D
F29E
F3D9
F476
F479
F4E9
F5E9
F670
F5E1
F4FB
F4B0
F4D8
F4B8
F454
F45E
F509
F5A6
F59A
F527
F4F2
F523
F561
F56E
F550
F501
F47E
F436
F4B8
F5C3
F63E
F5AB
F51D
F602
F84D
FA73
FB53
FB62
FBB3
FC62
FCAE
FC4A
FBD7
FBE1
FC22
FC2A
FC1A
FC40
FC5D
FC01
FB67
FB3C
FBA1
FBF3
FBC2
FB70
FB8A
FBE8
FC0A
FBFF
FC29
FC35
FB60
FA4D
FB7B
00A7
07F3
0CE4
0CB5
08FA
058E
047A
04B2
0476
03AD
0366
03E2
0444
03F5
0377
037F
03ED
040F
03AF
0353
0380
0419
04A2
04D3
04AB
0434
0383
02FB
0316
03C9
0457
041D
035E
0301
036D
03F7
03C1
0314
0365
05B6
0933
0BDF
0C94
0BF3
0B51
0B29
0B13
0AE3
0B1E
0C0C
0CE9
0CB1
0B89
0AAE
0AE4
0B89
0B9E
0B2A
0B07
0B7B
0BD5
0B8C
0B11
0B07
0B24
0ABE
0A29
0A8F
0BEF
0C3B
0959
03C7
FE44
FAC9
F8C0
F696
F445
F33D
F40E
F560
F5A9
F4FC
F476
F471
F444
F39E
F324
F363
F3EC
F413
F410
F4A8
F5C1
F63D
F581
F46D
F43A
F4EB
F58D
F5A0
F58E
F5B9
F5E2
F5B4
F56E
F579
F5A9
F586
F54A
F5F1
F7F6
FA88
FC60
FD0C
FD0A
FCE8
FCCF
FCB5
FC7B
FBF5
FB27
FA8D
FAC1
FBAB
FC6A
FC51
FBBB
FB83
FBCD
FBFF
FBE6
FBFC
FC58
FC40
FB67
FACE
FB6F
FC75
FC12
FA62
FA42
FE4A
055F
0B77
0DB6
0CCA
0AFA
093B
072B
04F3
03A6
03B6
043D
043D
03CF
03A6
03D5
03DC
03AE
03CD
044D
0475
03E4
0357
03AB
048A
04D7
043F
0397
03A2
041C
0447
03FB
03B7
03C4
03D3
0381
02FA
02B5
02D7
0321
034F
0361
03AF
04BE
06C9
0930
0AD0
0B2D
0AFE
0B43
0BFD
0C43
0BA5
0AD6
0AC4
0B64
0BE7
0BF5
0BF8
0C24
0C0F
0B82
0B0B
0B23
0B5D
0B19
0AB9
0B28
0C3F
0C9C
0B93
0A77
0AD1
0BA7
09F4
0469
FDAC
F9C6
F9CB
FB0A
FA67
F794
F4A9
F36F
F3D3
F4AB
F51B
F506
F4B2
F47A
F496
F4D2
F4B0
F417
F3A1
F3E0
F492
F4EE
F4C3
F4B1
F533
F5D3
F5BA
F4E7
F44B
F4A7
F5A5
F656
F647
F5CA
F55E
F530
F530
F53B
F534
F51F
F549
F631
F801
FA41
FC16
FCF8
FD04
FCAB
FC49
FC07
FBF1
FBF5
FBEA
FBC8
FBBC
FBE8
FC2B
FC4C
FC44
FC39
FC2D
FBFC
FBAB
FB89
FBC4
FC08
FBE4
FB77
FB3D
FB44
FB13
FAC6
FBA6
FF00
045C
0982
0C7E
0D2B
0C86
0B06
0879
055E
0335
02F7
03CB
0412
0368
02D6
032C
03EE
043A
0414
0424
0470
043A
0340
0261
0283
0362
03F7
03D3
036F
034E
0364
037A
039F
03E5
0408
03AF
0308
02B0
02E5
0333
0327
0305
038C
052C
07A4
0A31
0BE7
0C3C
0B96
0B0D
0B56
0C01
0C19
0B7B
0B07
0B6C
0C29
0C41
0BB0
0B5F
0BBB
0C17
0BC5
0B23
0AF5
0B50
0BB8
0BEF
0C02
0BC7
0B1B
0A98
0B1B
0C04
0ADB
05F1
FF23
FA99
FA3A
FB92
FAFF
F7FE
F515
F423
F459
F422
F38A
F3C6
F508
F617
F611
F585
F54C
F53E
F4C1
F405
F3C6
F418
F450
F40F
F3BD
F3C4
F3FA
F40A
F417
F47E
F52A
F593
F57C
F548
F55C
F59F
F5C8
F5D5
F5D4
F5A1
F558
F5A6
F724
F96B
FB44
FBEA
FBB3
FB79
FB91
FBB8
FBB5
FBB2
FBD1
FBD2
FB83
FB2C
FB54
FC25
FD36
FDE3
FDB6
FCC9
FBDE
FBC3
FC6B
FCF4
FCC3
FC4C
FC48
FC61
FB86
F9D2
F978
FCCB
035F
09FA
0DAA
0E24
0CD7
0AAD
07AB
045D
023A
0231
0377
0463
0435
037E
0305
02E5
02E0
02F4
032D
0358
0357
036D
03D4
043B
0432
03F0
0413
04B1
050C
0491
03AF
034D
0397
03D4
037C
02FF
0308
0374
0381
02DA
0223
026C
0450
0769
0A81
0C53
0C88
0BF6
0BC1
0C2C
0C82
0C32
0BAF
0BD0
0C88
0CE7
0C6B
0BB0
0B7D
0BAD
0B9D
0B41
0B26
0B62
0B55
0AB0
0A1C
0A4B
0ACE
0AB0
0A1B
0A44
0B45
0AFE
0741
00E9
FB94
F9F5
FB01
FB66
F94C
F5EE
F39F
F32D
F3AA
F422
F48E
F53B
F5F4
F63A
F5EB
F567
F511
F4EE
F4C0
F468
F410
F3FF
F440
F482
F45A
F3CF
F388
F427
F562
F622
F5B6
F4AF
F437
F4B5
F580
F5DE
F5E2
F608
F65E
F689
F6A1
F760
F931
FB5E
FCA7
FC91
FBBD
FB17
FAF7
FB21
FB4A
FB60
FB6A
FB69
FB6C
FB93
FBE8
FC49
FC8C
FCAB
FCB7
FCC6
FCE2
FCF5
FCD1
FC6C
FC20
FC46
FC87
FC15
FAF0
FAB4
FD61
031D
0988
0DB3
0E95
0D39
0AEE
0821
0521
02EB
026E
034F
0438
0456
03FE
03E3
042A
0488
04D3
0502
04D2
040E
031A
02BB
0319
0388
0392
039B
0416
049C
0473
03C7
038B
041C
04AC
0459
036A
02EC
033C
0397
0341
0298
02A8
0416
06B3
09AA
0BD6
0C5C
0B7E
0A8D
0A99
0B61
0BEE
0BED
0BEF
0C47
0C6B
0BDC
0B12
0AD4
0AE5
0A69
0987
0988
0AD2
0C02
0BD8
0B09
0B0A
0BAF
0B7C
0A51
0A05
0B64
0BDC
080B
0080
FA04
F858
FA16
FAFA
F916
F633
F4A1
F481
F4A0
F494
F4DB
F585
F5CE
F547
F476
F40D
F40D
F422
F448
F48C
F4A6
F466
F428
F448
F47E
F44E
F3E1
F3CD
F429
F473
F470
F499
F541
F5D9
F5A6
F4FF
F4EA
F57B
F5A0
F4FD
F4F0
F6D9
FA10
FC80
FD0E
FC7A
FBEF
FBA8
FB59
FB24
FB63
FBD1
FBC3
FB49
FB3C
FBF0
FCAF
FCE2
FCF0
FD4E
FD82
FCF6
FC36
FC59
FD3D
FD84
FC97
FBAD
FC0A
FCE6
FC85
FB43
FBFB
0095
074B
0C6B
0E19
0D43
0B61
08DA
05E0
0392
0319
0419
04F9
04D6
044E
042F
0434
03BA
0310
031A
03F1
04A3
047D
03D8
0380
03AC
03F6
03F8
03AD
0340
02DA
02BE
0332
0413
04BF
04B5
0426
03A1
036E
035B
032B
02EF
0315
043C
06AE
09D6
0C56
0D1D
0C68
0B7D
0B44
0B66
0B25
0A9D
0A93
0B0F
0B22
0A59
09A6
0A26
0B78
0C26
0BA7
0B07
0B4C
0C01
0C0C
0B74
0B42
0BB6
0BD8
0B3E
0B05
0BF1
0C50
0953
02C3
FC1E
F91D
F9C2
FAB7
F96A
F693
F47E
F402
F41B
F3DA
F385
F3BA
F464
F4EA
F502
F4D3
F499
F46D
F466
F491
F4BF
F4B2
F480
F47E
F4B3
F4C5
F4A2
F4BF
F54F
F5C4
F581
F4D5
F4A0
F51F
F5A3
F5A1
F572
F59F
F5E4
F5B6
F589
F6A3
F93D
FBBD
FC6F
FB71
FA4A
F9FC
FA5A
FB01
FBFF
FD2C
FDBA
FD1E
FC18
FBF9
FCEB
FDB7
FD7B
FCC4
FC71
FC69
FC18
FB9C
FB92
FBF3
FC16
FBC8
FB92
FBAE
FB8A
FB10
FBD6
FFB0
0600
0B8F
0DAB
0CA3
0A84
086B
0627
03E4
02BA
032F
043D
048E
041D
03F4
046F
04C8
0468
03DB
03E2
0446
0456
0407
03E3
0406
03FD
03A0
0364
039C
03E5
03A8
02F4
0270
0277
02B1
02BB
02BF
0319
03AC
03F4
03BD
0379
03F5
05C2
0898
0B3A
0C60
0C00
0B5B
0B84
0C36
0C74
0C08
0BBE
0C14
0C65
0BFB
0B55
0B89
0C75
0CB9
0BC7
0AD0
0AF9
0BA3
0B72
0A7E
0A26
0AD7
0B5E
0AF3
0AB5
0BCD
0CB8
0A4E
03FB
FD55
FA57
FADF
FB57
F955
F61E
F45E
F4C2
F5B4
F5CA
F542
F512
F567
F59E
F541
F46E
F38F
F313
F348
F40A
F4B3
F4C6
F484
F480
F4D0
F501
F4D8
F4B6
F50E
F5C1
F646
F658
F621
F5D3
F57D
F558
F5B5
F65A
F672
F5A6
F4F3
F5D6
F885
FB7D
FCF0
FC79
FB40
FAA6
FB0F
FBD7
FC35
FBEE
FB6C
FB48
FBA6
FC08
FBE4
FB63
FB40
FBC0
FC4E
FC46
FBE1
FBD1
FC27
FC3A
FBB7
FB40
FB80
FC0C
FBEF
FB6B
FC45
FFDC
0554
0A32
0CB2
0CE5
0BB8
09A5
06DD
041B
028A
02A1
038C
041A
03F6
03AF
03B9
03DB
03A8
032B
02E3
032B
03E2
048B
04B4
043B
0359
028D
0253
02C8
0380
03DD
03AA
033C
0306
0315
0318
02EB
02D3
0319
037F
0377
0302
031F
04E4
0824
0B4B
0CC6
0C7F
0BB9
0B94
0C10
0C81
0C96
0C88
0C7B
0C3E
0BC3
0B6B
0B7A
0B9E
0B5B
0ADE
0ADE
0B99
0C5B
0C5D
0BC7
0B5F
0B5D
0B3E
0AE5
0B1E
0C60
0D5B
0BBB
06AA
001B
FB37
F998
FA58
FB73
FB81
FA26
F7B3
F503
F344
F321
F403
F495
F42F
F37B
F383
F462
F53B
F55A
F50A
F517
F5BB
F657
F627
F51F
F415
F40E
F534
F685
F6BD
F5B9
F49D
F481
F543
F5E9
F5F3
F5C9
F5D4
F5D0
F557
F4C6
F4E0
F599
F60E
F5EB
F61B
F787
F9AC
FB24
FB5C
FB13
FB20
FB70
FB88
FB7E
FBC9
FC51
FC6C
FBE4
FB60
FB6A
FBAA
FB85
FB0F
FAD1
FB00
FB63
FBD9
FC53
FC73
FBDA
FAF9
FADD
FBC3
FC6C
FBD8
FB57
FD8B
02F6
08BB
0BB3
0BF2
0C06
0D24
0DA4
0B9F
07DE
0505
0462
04BE
047D
03B1
036B
03D8
041D
03C8
0359
0353
0372
0343
02F8
0328
03EF
04B2
04D8
0478
041E
0414
041B
03DC
0354
02D7
02C0
0323
03AD
03F6
03EC
03E3
0427
0490
04B3
0449
0375
02D4
0349
0561
089F
0B8D
0CE3
0CAE
0C29
0C48
0CB9
0C96
0BC4
0B1D
0B3A
0BC1
0C1D
0C38
0C2D
0BCA
0AF7
0A45
0A61
0B0A
0B47
0ACD
0A8A
0B43
0C36
0C19
0B2C
0B16
0C36
0C50
08E8
0281
FC71
F983
F99E
FAC0
FB48
FAC4
F949
F725
F545
F4BC
F570
F5ED
F529
F3EE
F3C2
F4D0
F5BE
F58A
F4BC
F470
F4D0
F516
F4D3
F481
F4BB
F561
F5DE
F5E4
F58F
F505
F46B
F40E
F42C
F49A
F4ED
F4F0
F4CB
F4A5
F47F
F466
F488
F4E6
F51D
F4E4
F4BC
F5A9
F7FE
FABE
FC7D
FCC2
FC35
FBB7
FB9D
FBBA
FBD1
FBCC
FBB1
FB95
FB8E
FB93
FB7E
FB59
FB7A
FC14
FCC8
FCF9
FCA4
FC6C
FCA3
FCC6
FC4C
FBA4
FBA8
FC31
FC27
FB6C
FC07
0028
0709
0CE1
0EA7
0D35
0BE2
0C5E
0D00
0B6B
07CB
0492
0379
03D5
041B
03F0
040D
04A7
04F5
0471
03B0
0390
03FF
0422
039F
031D
0357
0420
049D
0462
03D9
03AF
040D
0483
048C
0405
034C
02FE
036A
0439
04B3
047D
03F9
03C2
03CE
0383
02BA
026A
03C7
06CF
0A10
0C00
0C5C
0C03
0BC7
0BBB
0BA6
0B8E
0B93
0B88
0B26
0A9B
0A78
0AE3
0B3A
0AEA
0A5E
0A8B
0B90
0C45
0BA3
0A34
098E
0A5F
0B93
0BD7
0B50
0B26
0B6C
0A68
0684
008C
FB53
F916
F99E
FAF7
FB79
FAB9
F917
F711
F541
F453
F47D
F52D
F59A
F591
F578
F59C
F5D6
F5ED
F5F2
F60A
F617
F5D1
F535
F4A6
F483
F4CB
F538
F587
F58A
F532
F4B0
F46B
F498
F50A
F573
F5BC
F5E5
F5C5
F540
F4AB
F495
F4FB
F521
F498
F43A
F56C
F83D
FAEB
FBBE
FAE7
FA04
FA1D
FABB
FAFE
FAE5
FB11
FBB3
FC43
FC4A
FBED
FB93
FB67
FB67
FBA0
FBFA
FC28
FC0A
FBE5
FBF4
FC0D
FC05
FC2B
FCC1
FD2B
FC7A
FB38
FBDF
006B
0781
0D26
0EC0
0D9D
0CC5
0D16
0CB5
0A25
0694
046B
045C
04E0
0472
0350
02B3
0302
0399
03E2
03E4
03CE
038F
0337
0331
03D4
04CD
055D
0517
0446
038A
0347
0374
03D0
0407
03E8
039B
0393
040A
0499
04A6
0438
0402
046B
04CF
0435
02D1
024C
041D
07C7
0B1C
0C6C
0C07
0B64
0B40
0B36
0AF0
0AE8
0B95
0C60
0C44
0B4B
0AB8
0B5D
0C6F
0C8F
0B9A
0AB3
0A7C
0A59
09C1
0969
0A47
0BCF
0C5E
0B7A
0AA4
0B30
0BF1
0A23
04CC
FE4D
FA15
F960
FA9E
FB92
FB29
F98A
F759
F557
F435
F423
F491
F4C4
F49D
F48C
F4C2
F4E1
F4A4
F462
F48C
F4FB
F524
F4E7
F4A9
F4A3
F48D
F41C
F393
F37C
F3F2
F482
F4C6
F4D7
F4FC
F533
F545
F524
F4FC
F4EC
F4F6
F51C
F557
F57E
F574
F580
F63F
F806
FA55
FC1F
FCBE
FC87
FC5A
FCB6
FD58
FD9A
FD24
FC4A
FBC8
FC11
FCCC
FD20
FC9A
FBB4
FB49
FB9E
FC38
FC8A
FC94
FC95
FC88
FC4A
FC1E
FC6C
FCDF
FC7D
FB38
FAF5
FE01
0434
0A5C
0D29
0C8B
0B5F
0BDA
0D0C
0C70
0948
0598
03BB
03EA
0483
0449
038D
0343
039C
03FE
03F4
03A3
0362
034D
035E
03A5
041E
0488
0494
0448
03FB
03EB
0401
03FB
03BC
034C
02CC
0282
02C1
0388
0448
0464
03FF
03EF
049C
053B
04C6
03A0
039C
05EC
0973
0BC7
0BD4
0ACF
0A7C
0B10
0B75
0B28
0AE8
0B69
0C3C
0C8F
0C6E
0C80
0CC9
0C94
0BBC
0B3F
0BE1
0CD6
0CA5
0B4E
0A6D
0B08
0C22
0C45
0BBC
0BFF
0D0F
0C98
0889
01E6
FC1F
F9AD
FA10
FB1A
FB4B
FA6E
F8C0
F690
F493
F3A2
F3D4
F44C
F449
F402
F429
F4CD
F541
F513
F493
F444
F434
F437
F45E
F4BA
F4F0
F48A
F3BA
F34D
F3C2
F4AC
F53A
F51D
F4B5
F473
F46D
F484
F4A9
F4C9
F4CF
F4D7
F519
F575
F56F
F4F7
F4E5
F626
F87E
FA80
FB14
FA93
FA3A
FAAC
FB7A
FC07
FC47
FC70
FC70
FC2C
FBF3
FC2B
FCBD
FD27
FD1D
FCD0
FC83
FC46
FC21
FC3E
FC95
FCB7
FC57
FBDB
FBD8
FC0B
FBAD
FB16
FC36
007D
069C
0B54
0CBA
0C06
0BAA
0C4B
0C5C
0A97
07C6
05BA
0521
052E
04FC
0486
043E
044D
0481
049C
0470
03DA
02F3
022E
0202
0267
02D9
02FD
02F4
02F8
02F9
02DA
02D0
0324
03A5
03C8
0368
030C
0346
03F4
046B
0452
040B
0416
0446
03FD
0337
0305
04A5
0817
0BC7
0DD3
0DB8
0C9F
0BF4
0BF7
0BE8
0B5B
0AC5
0AB5
0B0A
0B53
0B92
0C0E
0C93
0C87
0BE5
0B91
0C15
0C9D
0BFB
0A89
09F1
0AD4
0BBE
0B43
0A47
0AC0
0C6B
0C2E
07A7
0072
FAD2
F935
FA3D
FB24
FAD4
F9D8
F882
F687
F431
F2A7
F289
F323
F369
F355
F3A5
F484
F53A
F53C
F4E1
F4B6
F4BE
F4C3
F4E2
F539
F571
F530
F4D6
F50A
F5B0
F5E0
F520
F42B
F40A
F4BD
F553
F53A
F4CD
F48E
F484
F4A8
F533
F5FC
F624
F544
F482
F594
F88B
FB6E
FC5E
FB9E
FAF0
FB4A
FC03
FC36
FC02
FBF8
FC17
FC0B
FBF6
FC30
FC8D
FC88
FC25
FC08
FC89
FD30
FD5B
FD10
FCC4
FCAA
FCAE
FCEF
FD76
FD8D
FC74
FB23
FC35
0112
07A9
0C2D
0D03
0C0B
0BC3
0C3D
0BB2
0963
06A6
0503
0483
046E
04A7
055E
05F8
057F
041F
0325
034E
03CF
0382
0290
022B
02D4
03BA
03E9
0381
0335
033A
034A
035E
03AF
0419
0429
03DC
03C2
0427
047C
0415
033E
02FD
03AE
045E
0409
0317
0320
0523
0871
0B5C
0CB3
0C90
0BE5
0B87
0B90
0B9E
0B74
0B40
0B57
0BC3
0C3F
0C8C
0CA7
0C95
0C2F
0B60
0A88
0A30
0A63
0AA7
0ABA
0AD2
0B0A
0B10
0ADA
0B20
0C57
0D2D
0B26
0578
FEC1
FAD6
FACC
FC29
FC33
FAF8
FA4B
FAA4
FA76
F888
F5BA
F3E6
F3AA
F41F
F467
F48F
F4DA
F503
F4BF
F462
F466
F4AD
F4CD
F4BA
F4AF
F4A5
F46F
F440
F481
F513
F54A
F4DA
F46B
F4AE
F538
F506
F409
F35E
F3AB
F43C
F445
F423
F49D
F56E
F5A5
F52C
F4EF
F559
F59C
F517
F4C2
F620
F8FA
FB51
FBE3
FB9C
FBF2
FCC9
FCFA
FC43
FB88
FB6E
FBA7
FBC9
FBF0
FC3C
FC48
FBC5
FB46
FBAF
FCE7
FDD3
FDCC
FD43
FCBD
FC2A
FBA7
FBED
FD03
FD87
FC78
FB75
FD9E
03BB
0A8B
0DEB
0D2E
0B5B
0B4A
0CD5
0E15
0DFE
0CB5
0A6B
0752
0475
0339
03B5
046C
0419
0328
02E6
03A1
0455
042D
0392
0367
03C7
041A
03FF
0398
0330
030B
0365
042D
04C2
0488
03BA
034A
03C9
04A8
04E1
0428
033D
02F0
0347
03B5
03E6
03FE
0431
0475
0490
0459
03F5
0400
052E
078E
0A36
0BEB
0C3C
0BCD
0B89
0BB8
0BFF
0C10
0C0A
0C1B
0C23
0BEE
0B98
0B70
0B87
0B97
0B71
0B32
0B03
0AD7
0AA2
0A9D
0AFA
0B6A
0B5E
0AF3
0B10
0C15
0C89
0A0F
0426
FD86
F9DC
FA15
FBB4
FBF8
FADA
FA3F
FAE7
FB49
F9C1
F6D5
F49A
F433
F4CC
F511
F4D0
F4AE
F4E2
F4F8
F49A
F3FE
F393
F396
F3FF
F492
F4F4
F4FF
F4DC
F4C6
F4B2
F46E
F413
F40D
F480
F4E3
F4AB
F427
F421
F4AA
F4F1
F492
F43B
F496
F537
F55D
F52D
F55C
F5D8
F5C3
F4F4
F4B5
F64A
F91C
FB41
FBCF
FBAB
FBF0
FC7B
FCA7
FC8A
FC96
FCAA
FC5C
FBE3
FBD5
FC1F
FC0B
FB67
FAF8
FB5F
FC2C
FC8C
FC90
FCE5
FD6D
FD4B
FC76
FC0A
FC75
FC90
FBA5
FB65
FE54
0465
0A7B
0D94
0DA2
0CB8
0C57
0C71
0CA2
0CE5
0CC8
0B29
07BC
0423
0270
02EE
041C
0496
0444
03CC
03B0
040B
04A3
0501
04C5
0420
03BB
03F3
0450
0424
039B
0386
0415
0478
041E
038C
0380
03CF
03D5
0386
035D
036D
0350
02F1
02D1
034C
0409
0484
04C2
04FE
04F4
044E
03C8
04E5
07EE
0B0B
0C2C
0B63
0A8C
0AEC
0BFB
0C92
0C71
0C2B
0C23
0C2C
0C14
0BFB
0BF4
0BC8
0B68
0B33
0B71
0BC4
0B9F
0B22
0AFA
0B52
0B76
0AD7
0A13
0A64
0BD2
0C4D
0959
02F6
FC63
F938
F9D6
FB5A
FB38
F9FC
F9D8
FB30
FBD0
F9CE
F635
F3D3
F3DA
F4CE
F4E1
F42A
F3EA
F483
F526
F52E
F4D2
F490
F48B
F49E
F49D
F45E
F3D4
F341
F31C
F38B
F41B
F450
F454
F4B2
F564
F5C2
F586
F52D
F526
F530
F509
F4FB
F53C
F554
F4DC
F45D
F49D
F548
F539
F452
F430
F654
F9F9
FCC5
FD7A
FCFB
FC7B
FBF7
FB1E
FA84
FADA
FBAD
FC07
FBDE
FBEA
FC46
FC3E
FBA7
FB61
FC15
FD11
FD31
FC92
FC4F
FCAC
FCD4
FC80
FC7F
FCEA
FC7B
FAEB
FAB2
FE95
05BA
0BE8
0E00
0CFB
0BE0
0C01
0C62
0C3D
0C2D
0C72
0BBE
0906
0578
0363
0380
0489
0523
0521
04F7
04E5
04F5
0527
054B
04FC
041F
0331
02CB
02E1
02F0
02E2
0329
03DB
0462
046B
046C
04BB
04E0
0462
03BA
03B0
0425
0454
03FC
039D
038B
0378
033E
035F
042F
04D7
044E
033C
03B4
068C
09FE
0BB3
0B6D
0ABB
0ABA
0B29
0B86
0BDB
0C38
0C43
0BCC
0B63
0BA3
0C25
0BFC
0B31
0AF3
0BD2
0CBA
0C60
0B20
0A73
0AD4
0B3A
0AD2
0A4C
0AD0
0BE5
0B3D
070A
005D
FABB
F8E4
FA3F
FBC8
FB64
F9ED
F9A8
FB21
FC45
FAE2
F76F
F48D
F3ED
F4A1
F4D6
F433
F3CD
F443
F4E7
F4D6
F421
F39A
F3D3
F4A2
F578
F5E0
F5B6
F51F
F473
F408
F3DD
F3B4
F37E
F382
F3F1
F499
F524
F570
F57D
F551
F52C
F55D
F5C9
F5E9
F58A
F539
F579
F5E1
F59E
F4C6
F4A9
F65D
F953
FBD4
FCCA
FC82
FBC6
FB00
FA7C
FA9F
FB55
FBDD
FBC2
FB8A
FBD8
FC6E
FCA3
FC7A
FC88
FCD1
FCAA
FBE6
FB74
FC1A
FD29
FD6F
FD15
FD43
FDD0
FD33
FB6B
FB65
FFBC
06F6
0CAB
0E50
0D66
0CB6
0CE3
0CCC
0C21
0BD9
0C0C
0B24
0825
0492
02D1
035A
0492
0508
04B3
0433
03F1
040B
0475
04D7
04C7
044C
03F7
041E
0451
03FC
035C
0346
03D2
0427
03C1
0336
0327
0351
0338
031E
0374
03E1
03BE
0343
0355
0429
04D2
0495
03FD
03F5
043C
03DF
0319
039A
0640
09A5
0BBA
0C20
0C0B
0C5B
0CDA
0D26
0D41
0D19
0C5A
0B2C
0A89
0B2B
0C5A
0CA3
0BB8
0ADC
0B12
0BB8
0BA2
0AE0
0A75
0AAB
0AB2
0A14
099D
0A39
0B32
0A50
0611
FFA6
FA51
F880
F9A8
FB2A
FB2C
FA52
FA72
FBFE
FD33
FC25
F91B
F63A
F504
F4EE
F4B0
F416
F3DD
F452
F4E2
F4F9
F4A6
F448
F40F
F404
F43A
F49C
F4C4
F460
F3C8
F3B4
F44D
F4EE
F50D
F4ED
F515
F577
F59B
F557
F4F2
F4A1
F460
F432
F438
F479
F4CD
F512
F549
F55F
F518
F47C
F442
F54C
F797
FA02
FB6B
FBC2
FBBE
FBDC
FC07
FC03
FBD1
FBA6
FBBA
FC11
FC63
FC6A
FC4E
FC91
FD55
FDF1
FD9E
FC80
FBA9
FBD2
FC8B
FCFD
FD20
FD62
FD72
FC99
FBA5
FD0F
0229
08C8
0D17
0D93
0C44
0BC6
0C55
0C80
0BD9
0B78
0BBB
0B1E
0843
0442
01C8
020A
03A7
0490
0432
0382
037C
0418
04A2
04A9
045F
0438
044E
0458
040F
03A0
0380
03DA
0434
0401
0366
0310
033A
0365
033F
032C
0392
0419
0433
0405
0431
04C4
0507
048B
03E4
03D7
0438
0444
0408
0497
0684
08FE
0AD4
0BCE
0C5D
0C8E
0C20
0B6C
0B50
0C02
0CA5
0C7E
0C04
0C1F
0CA0
0C72
0B56
0A74
0AB9
0B7C
0B91
0B1C
0B41
0C2F
0CAE
0BFA
0B17
0B52
0BD9
0A17
04E1
FE67
FA36
F9A5
FAEF
FBA9
FB3B
FABC
FB15
FBEE
FC3D
FB48
F913
F642
F3CD
F28D
F2A0
F34F
F3C8
F3E1
F3FB
F44B
F494
F498
F478
F46B
F45B
F412
F3C5
F3F6
F4C3
F58B
F594
F4CC
F3BB
F2F6
F2D0
F368
F495
F5C2
F633
F5B1
F4CB
F447
F464
F4DA
F566
F5ED
F620
F582
F42D
F326
F393
F5A5
F882
FB0A
FC7E
FCAE
FBF9
FB3C
FB42
FC04
FCA8
FC7E
FBD8
FB85
FBAD
FBDA
FC01
FCA8
FDC9
FE5E
FDB5
FC96
FC42
FCA5
FC90
FBC1
FB85
FCA6
FDC2
FD13
FBAD
FD1A
0300
0A61
0E8A
0E1F
0BEC
0B09
0BB3
0C60
0C8B
0CEA
0D6B
0C8B
096C
0594
0384
03E9
0517
053B
044A
0388
03BE
0478
04BA
0417
02F8
0215
01DD
0244
02F0
037A
03A6
037B
032B
02F4
0308
0379
041D
049B
04AF
0466
040C
03EB
041F
047B
0499
042E
035A
028E
0225
023D
0302
04C6
0782
0A54
0BFB
0C0F
0B77
0B5A
0BCC
0C08
0BCC
0BBC
0C43
0CC6
0C8E
0BF9
0BF1
0C6C
0C58
0B48
0A67
0AEC
0C39
0C90
0BA9
0B33
0C1A
0C6E
0954
02C8
FC42
F938
F9D4
FB91
FC58
FC14
FB8E
FB08
FA6F
F9F2
F99C
F8D8
F727
F523
F3FD
F410
F48C
F4B2
F4BD
F534
F5D7
F5E7
F556
F4E7
F502
F514
F49A
F40B
F42D
F4E7
F567
F537
F497
F3DE
F32E
F2C7
F317
F41C
F50F
F540
F50A
F551
F612
F645
F563
F437
F3B2
F3CF
F435
F54E
F7B5
FACB
FCE8
FD33
FC8C
FC44
FC7E
FC83
FC32
FC1D
FC47
FBF8
FB1D
FABE
FB5B
FBEF
FB87
FAEC
FB88
FD14
FDC2
FCE4
FBED
FC21
FC82
FBA0
FAD8
FD73
0414
0ADD
0DA3
0CB0
0BA0
0C63
0D70
0CF7
0BC8
0BC0
0C8B
0BCB
0883
04BC
0310
03A5
0494
049A
0423
03F1
03FA
03DA
0394
0376
0399
03D6
040F
043A
0437
03E9
0382
0370
03DA
0465
04AE
04BA
04C3
04C1
0488
0432
040C
041C
040D
03A3
031C
02F9
0369
03EE
03D3
0327
0309
04A2
07B6
0A9C
0BE0
0BBB
0B8F
0C0E
0C76
0BEB
0AE7
0AA0
0B30
0B71
0AD4
0A56
0AFC
0C29
0C76
0BBD
0B37
0B76
0B77
0A6B
0979
0A5D
0C5B
0C1D
0770
003F
FAD5
F987
FAF8
FC69
FC97
FC0B
FB9A
FB75
FB72
FB57
FAAF
F8F5
F661
F42C
F375
F40E
F4C8
F4DD
F49B
F4AF
F531
F59E
F58C
F516
F4A3
F478
F489
F4A5
F4A4
F48B
F489
F4C4
F51D
F54B
F53D
F52B
F530
F51C
F4D6
F4C4
F55E
F667
F6EC
F65C
F550
F4D9
F52A
F589
F5A1
F632
F802
FA90
FC74
FCF1
FC9C
FC59
FC3A
FBDE
FB6E
FB8C
FC47
FCDD
FCC8
FC61
FC38
FC4A
FC58
FC7B
FCCC
FCDB
FC2E
FB36
FAF1
FB5C
FB4C
FA88
FB3E
FFC6
06F5
0C69
0D48
0B65
0A91
0BD9
0D0F
0CA1
0BC9
0C22
0CB0
0B10
072C
03D8
034E
0486
050E
043A
034E
0326
0352
0358
037D
03E8
0400
0360
02C9
0348
0498
054B
04C2
03FF
0420
04CD
04F8
0482
042F
044D
045B
0416
03EF
0435
045E
03CE
02E5
02A9
033A
0374
0281
0160
020B
0519
08DD
0B20
0B56
0AD6
0B0B
0BEA
0C51
0BB4
0ADB
0ABB
0B1B
0B09
0A79
0A79
0B9B
0CE6
0D0D
0C35
0B9C
0BAA
0B58
0A15
093D
0A54
0C1D
0B26
05E0
FF03
FACA
FA79
FBB6
FBF5
FB27
FAC9
FB6B
FC1D
FBD7
FA8C
F8C3
F6EC
F575
F4D3
F4EB
F4F2
F46A
F3DB
F411
F4F4
F5AE
F5CB
F591
F557
F51B
F4CA
F48C
F47D
F45D
F407
F3EC
F491
F59E
F615
F5A8
F52D
F55A
F5C5
F5BE
F578
F598
F5EE
F59D
F488
F3CF
F455
F578
F5F8
F5F1
F6E4
F98F
FCA4
FE3A
FDED
FCE7
FC47
FC36
FC64
FC93
FC99
FC60
FC2F
FC83
FD5C
FDF5
FDAD
FCE4
FC7A
FC7F
FC3B
FB8C
FB41
FB9C
FB7A
FA1F
F94F
FBFB
028A
097D
0CE0
0C6F
0B43
0B97
0C76
0C0E
0AD7
0ACF
0C27
0C72
09B7
053D
0239
0232
03B1
047B
03FD
0322
02A9
0289
02A7
0324
03DF
0453
044E
0449
0497
04B8
0402
02DB
0285
037C
04A7
04AB
03B2
0330
03E9
04FF
0526
044A
037F
0383
03FA
0422
03D2
0360
0302
02DB
0377
0590
08E8
0BE4
0CE8
0C05
0AED
0B0F
0C1E
0CC0
0C4D
0B65
0AD6
0AA2
0A65
0A41
0A9A
0B2A
0B16
0A33
097E
09D6
0AB1
0AED
0AA6
0B33
0CDF
0D75
0A4A
03A4
FD0F
F9DB
F9FF
FAE7
FAB4
F9C6
F965
F9F3
FAC3
FB03
FA4D
F8AB
F69E
F514
F4B8
F528
F555
F4DF
F47F
F4CF
F548
F50D
F448
F402
F4A8
F56D
F55D
F48E
F3EF
F41B
F4D2
F57F
F5D4
F5C6
F561
F4E5
F4AA
F4B3
F4B0
F49F
F4ED
F5A4
F603
F57C
F4B2
F4D3
F5EE
F6B5
F642
F584
F63C
F8AC
FB31
FC37
FBDE
FB4F
FB2D
FB51
FB93
FBFD
FC71
FCBF
FD02
FD73
FDE0
FDCD
FD44
FCF8
FD3B
FD55
FC9D
FBD2
FC34
FD4F
FD28
FB5A
FABC
FE67
058A
0BBD
0DCE
0CE1
0C2C
0CC0
0D1B
0C66
0C19
0D7C
0F03
0DC9
095B
0488
023B
028C
0371
037C
0303
02E6
0332
0367
0367
0383
03DA
042B
0456
0483
04B9
04B8
045E
03EE
03CC
03FE
0428
03F8
0383
0325
031A
0349
0379
0393
03B6
040B
0492
0509
050E
0474
038E
0324
0401
0655
094E
0B7C
0BF4
0B31
0A93
0AE9
0BAB
0BD2
0B29
0A72
0A5C
0ABE
0B14
0B3D
0B50
0B09
0A1D
090A
08CE
097C
09E4
094D
08DE
0A34
0C8A
0C90
07E9
0054
FA52
F89C
F9D8
FB00
FAD9
FA65
FAAE
FB62
FB9C
FAFD
F9A5
F7BF
F5A8
F429
F3EC
F49C
F526
F4FD
F4A0
F4B6
F520
F55A
F551
F555
F57D
F59B
F5A4
F5B1
F5A7
F559
F4FC
F517
F5BD
F62A
F599
F45C
F394
F3D7
F4AB
F568
F5E7
F616
F5B2
F4F4
F4D3
F5D0
F6E3
F69A
F53B
F4E4
F703
FA6B
FCA4
FCD5
FC52
FC69
FCC0
FC7A
FBCB
FB90
FBF6
FC78
FCD3
FD1C
FD1C
FC82
FBC0
FBDE
FD00
FDDF
FD6F
FC7D
FC7F
FD1E
FC9F
FB1C
FB9A
0076
07BB
0CDD
0DBE
0C85
0C2E
0CEC
0D01
0C0D
0BA4
0C84
0CF0
0AE5
06F9
03C5
02DE
037E
041F
0442
0451
0482
0484
0411
035E
02E2
02E1
0342
03B2
03C7
0355
02B1
027A
02E5
0379
03A2
035B
030C
02FB
032E
038B
03E5
0405
03ED
03EC
043A
048F
0464
03A1
02CE
0284
02F4
0426
0648
092B
0B9F
0C3F
0B2F
0A42
0AE1
0C4E
0CAD
0B6F
09F2
09AD
0A96
0B9B
0C21
0C46
0C1B
0B6A
0A75
0A02
0A43
0A73
0A1E
0A13
0B25
0C3E
0ADD
05E6
FF56
FA8B
F918
F9C9
FA97
FACB
FAF1
FB78
FBFF
FBD5
FA91
F85A
F5EF
F45B
F424
F4C3
F534
F511
F4E1
F52F
F5AE
F5AE
F524
F4C9
F50F
F588
F591
F532
F4E8
F4E9
F501
F505
F4FD
F4E7
F4B7
F493
F4C9
F54F
F5A5
F576
F525
F539
F584
F563
F4EC
F4FE
F5DF
F68C
F625
F576
F624
F870
FAB8
FB7E
FB37
FB5C
FC31
FC8F
FBD4
FAF4
FB18
FC14
FCF3
FD58
FD85
FD6F
FCC6
FBDF
FB97
FC12
FC5E
FBE0
FB6A
FC06
FD1E
FD42
FCD4
FE5A
032D
0917
0C94
0CE2
0C5C
0CE5
0DA8
0D0A
0B8E
0B27
0C1A
0C2A
099B
05B4
033E
032A
03F2
03F5
0344
02EB
0356
03FB
043B
0405
03B1
0386
0387
039E
03C3
040F
04A0
054F
058A
04E6
03D5
0357
03B9
043F
0435
03DF
03CA
03CE
0363
02B2
0285
030C
036D
0320
0325
0504
08A1
0BEF
0D2F
0CA8
0BC6
0B43
0AF5
0AD8
0B38
0BE9
0C1F
0B6F
0A75
0A15
0A73
0AF8
0B40
0B6A
0B8D
0B72
0B1A
0AE5
0AE9
0ABA
0A41
0A36
0AF1
0B22
08B5
033B
FCF5
F8F1
F858
F9C2
FAE8
FA90
F8ED
F6E9
F56A
F4D8
F4DB
F4BC
F453
F434
F4BE
F55E
F540
F47D
F404
F469
F540
F5CA
F5E1
F5DE
F5E8
F5D8
F5BA
F5D4
F615
F60A
F5AC
F58F
F5EB
F618
F57D
F497
F460
F4EA
F555
F528
F4FC
F57A
F650
F6F2
F7D7
F9DA
FC69
FD9F
FCBB
FB66
FB8C
FCB8
FCE8
FB8B
FA5B
FAC7
FBDF
FBCA
FA8C
F9FD
FB09
FC6E
FCB1
FC15
FBB6
FBAC
FB50
FAC3
FAD3
FB6A
FB7E
FB2D
FCA0
0181
0816
0C6F
0CD8
0BB8
0C3C
0E36
0EAC
0BE9
078C
045B
0346
033C
0325
0304
033C
03AB
03E8
03EE
03FC
0412
0401
03CC
03A4
039B
03B1
03FA
0471
04CF
04CE
0483
0421
0394
02B7
01E4
01D3
02A7
0369
0325
0248
0225
0307
03AD
0341
02F7
04BC
0886
0BF8
0CE9
0BA4
0A35
0A03
0AB4
0B42
0B58
0B46
0B4E
0B6D
0B97
0BB4
0B8A
0B18
0AC8
0AF4
0B5E
0B79
0B21
0AA8
0A41
09DC
09B9
0A87
0C38
0D0E
0AB4
04D3
FDFE
F985
F88E
F9AF
FAD8
FB02
FA17
F844
F5E9
F3E1
F325
F3DA
F50A
F583
F4F9
F428
F3FE
F4BA
F5C4
F63B
F5C5
F4F1
F4B0
F543
F601
F625
F5AD
F529
F4FB
F516
F54D
F59B
F5E6
F5E6
F582
F51C
F531
F5B1
F614
F611
F5D1
F57E
F52D
F566
F702
F9F3
FCAE
FD8F
FCBB
FBE1
FC1C
FCBF
FCB8
FC49
FC77
FD15
FCD0
FB5F
FA64
FB35
FCBE
FCDA
FB4C
FA07
FA65
FB6E
FBA0
FB49
FBC8
FCEC
FCED
FB8B
FB89
FF9E
06A2
0C4B
0DD3
0C96
0BC3
0C7D
0D15
0BA2
0850
04EB
02F5
029E
032A
03B5
03C4
0383
0370
0396
0375
02D2
024E
029B
0374
03DF
0383
0319
035C
03FE
0432
03F6
0406
048A
04B1
03F8
0313
02EC
0351
036B
0325
033F
03E6
042B
0377
02D0
03E8
06E2
09F7
0B82
0BA0
0B6C
0B5B
0B19
0A98
0A4F
0A65
0A69
0A0F
09C9
0A29
0B01
0B93
0B8C
0B57
0B65
0BAF
0BFF
0C3B
0C14
0B26
09DC
0995
0B06
0C88
0B12
0579
FE34
F949
F88A
FA5D
FBF3
FBDC
FA49
F7E9
F576
F3F9
F437
F5A0
F687
F5DC
F461
F3BC
F489
F5D4
F66C
F61D
F57B
F4FA
F4BC
F4DF
F561
F5D2
F5B3
F538
F534
F60E
F70E
F721
F61A
F4DA
F437
F438
F47F
F502
F5DD
F697
F660
F51F
F3F6
F452
F67E
F953
FB5C
FC12
FC04
FBF6
FC2B
FC7F
FCDC
FD45
FD91
FD62
FC9A
FBBB
FB86
FC16
FC9E
FC51
FB65
FAC0
FABD
FADB
FAC7
FB16
FC4E
FD98
FD63
FBC4
FB56
FEBC
0556
0B5D
0DBC
0D04
0C1B
0C8A
0D06
0B89
07F6
0443
025F
0290
03AF
0473
0465
03DE
037E
038B
03B2
037E
0307
02E5
0352
03CD
03D2
0396
039D
03CF
0396
02D9
0260
02D6
03CB
0432
03B9
030B
02C3
02CC
02FC
038A
045D
048A
0370
022A
02EC
0688
0B1D
0DD1
0DA3
0C07
0AE6
0AB7
0AC8
0A9F
0A6A
0A78
0ADB
0B7A
0C14
0C3A
0BB8
0AEE
0A81
0A95
0AB7
0A93
0A61
0A58
0A22
097F
092A
0A23
0BAE
0B21
06A0
FFAA
FA17
F861
F9A0
FB28
FB56
FA50
F8BB
F6E2
F52F
F46D
F4E0
F5AA
F5C4
F53B
F4EC
F51B
F52A
F4B4
F44F
F4B0
F58A
F5DD
F558
F4CB
F501
F5A7
F5DA
F56A
F50E
F559
F60A
F67D
F671
F629
F5FD
F60F
F652
F69F
F6AF
F631
F53D
F492
F51E
F716
F992
FB37
FB5C
FA9F
FA4A
FB08
FC43
FCE3
FC96
FC0D
FBF8
FC31
FC27
FBD6
FBD3
FC5A
FCD1
FC90
FBD7
FB6B
FB85
FBB0
FBC8
FC42
FD20
FD5A
FC4D
FB74
FD78
02FF
093E
0CA1
0CA1
0BE4
0C89
0D7D
0C4D
08BA
0536
03D8
041A
0426
0379
0328
03C7
0458
03BB
026B
01E7
02B4
03C8
040B
03AD
0391
03E6
03F5
0347
0269
023F
02DD
0370
0351
02C6
0298
030E
0397
037F
02CE
024A
0285
0322
0353
0313
0382
05B2
093B
0C50
0D68
0CA1
0B64
0ADE
0B10
0B5C
0B76
0B8A
0BBF
0BEB
0BD8
0B80
0B0A
0A98
0A32
09E0
09CF
0A39
0B07
0B9A
0B43
0A28
0986
0A75
0C32
0C1C
082A
0176
FBAB
F998
FABC
FC5A
FC75
FB13
F913
F6DA
F48D
F2DB
F28F
F371
F459
F486
F463
F4AC
F54F
F5BD
F5D2
F5D7
F5D3
F573
F4C3
F468
F4DB
F5C1
F665
F69C
F6CF
F71C
F709
F64C
F564
F505
F53B
F591
F5C3
F5EA
F5FA
F5AC
F4F5
F461
F4AD
F622
F859
FA8B
FC0F
FCAB
FCA0
FC7E
FC9F
FCCD
FCA2
FC2C
FBE5
FBEF
FBE9
FBA2
FB71
FB93
FBA9
FB55
FB05
FB62
FC1E
FC2B
FB64
FB1E
FC40
FD7A
FCDC
FB35
FC2C
01D5
096C
0DF7
0DCD
0BFD
0BFC
0D69
0D2F
0A02
0616
0435
0484
0507
0481
03A6
039C
0468
0521
051A
0470
03BC
036B
0366
0346
02DA
0274
0286
0314
038E
037E
0314
02DA
02EB
02DE
028B
0250
0269
0291
029F
02F2
03C2
0461
03FD
0310
0355
05CE
0954
0BAD
0BF1
0B39
0AE6
0B0C
0AF3
0A76
0A2D
0A6D
0AE3
0B2B
0B3C
0B3E
0B33
0B16
0B01
0B0D
0B34
0B6F
0BCE
0C29
0BEE
0ADF
09DB
0A1A
0B37
0ACF
06ED
00A3
FB65
F9B3
FAE1
FC57
FC49
FAC6
F89F
F657
F45D
F361
F3B6
F4A0
F4F6
F470
F3D9
F3F3
F4A4
F557
F5BB
F5E7
F5F1
F5D9
F5C2
F5E5
F621
F5FE
F55F
F4E8
F547
F63A
F6B2
F61A
F512
F4AF
F52B
F5BC
F5B2
F557
F56D
F5FA
F628
F583
F4F1
F5E6
F89E
FB85
FCC0
FC1C
FB26
FB4F
FC62
FD1C
FCE9
FC75
FC83
FCD6
FCAA
FBDA
FB0B
FABB
FAB7
FAB9
FAFD
FBCD
FCAE
FCD3
FC51
FC39
FD0F
FDC5
FD22
FBF6
FCE6
0177
07C6
0C22
0CD3
0B96
0B1E
0BD6
0BD8
09C3
0692
0468
0415
0484
0452
036B
02BE
02EC
03A2
042A
0432
03EC
03A9
0397
03AE
03D6
03F4
03F6
03D5
03A8
03A0
03D8
0426
042C
03BC
032A
0306
0378
03F9
03F5
038C
0364
03AE
03D8
037D
0349
046F
0735
0A5E
0C40
0C45
0B46
0A83
0A98
0B4A
0BF9
0C1E
0BAD
0B26
0B12
0B56
0B3F
0A7F
09B9
09CD
0AC0
0BB6
0BFE
0BB7
0B59
0B0B
0ABF
0AA8
0AD2
0A58
07D4
0311
FDD2
FA68
F9A6
FA86
FB67
FB2D
F984
F6DD
F46C
F381
F44B
F57A
F5A6
F4F6
F4BB
F56F
F604
F58D
F4A0
F468
F4E7
F527
F4DF
F4E3
F5AF
F662
F5E6
F491
F3CC
F429
F4B2
F476
F3D7
F3CC
F481
F55C
F5FA
F64D
F611
F517
F42C
F4DF
F7C1
FB44
FD16
FC96
FB5A
FB2C
FC25
FD02
FCDC
FBED
FB0D
FAEF
FBAB
FC90
FCA7
FBCE
FB1E
FBB3
FD18
FD9C
FC7E
FB15
FB12
FC19
FC53
FB81
FC21
0071
070D
0C07
0D3A
0C67
0C6E
0D89
0D4E
0A3F
05F9
0364
0361
043D
042A
0340
02D1
036B
043D
044C
0398
02EA
02C9
0306
0343
0376
03C9
0430
0475
048D
0492
0473
0406
037B
0365
0401
04A9
0484
03A8
031C
0377
03F5
038F
02B7
033F
0615
09CB
0BFE
0BE9
0AFD
0AEB
0BC4
0C60
0C1A
0B78
0B3D
0B73
0BAB
0BBB
0BC9
0BC2
0B61
0AC4
0A86
0AF6
0B86
0B6E
0AD0
0AAC
0B6F
0BCD
09AA
046D
FE1B
F9C7
F8E1
FA44
FBB8
FBD4
FA70
F805
F550
F362
F323
F458
F587
F56B
F465
F3E7
F479
F512
F4AC
F3C5
F3A4
F47A
F51A
F49F
F3A7
F37F
F46D
F561
F549
F44E
F37F
F3A3
F48F
F57B
F5C2
F571
F541
F5BB
F66B
F65E
F59C
F594
F780
FAA1
FCD3
FCE2
FBCE
FB68
FC20
FCDD
FCB4
FC01
FB90
FB90
FBBE
FBF9
FC28
FC03
FB8E
FB70
FC1D
FD01
FD2B
FCBE
FCC8
FD6F
FD48
FB89
FA46
FCC8
0347
09DE
0CAF
0C12
0B65
0C56
0D18
0B56
0781
042C
02F5
0334
0396
03C7
0419
0479
0496
048F
04B3
04D1
048A
0416
0419
04A3
050A
04CE
043B
03F2
0412
043A
042E
041A
041D
0414
03FA
0418
047D
04B8
0461
03A8
0317
0326
0437
067C
0960
0B7A
0BC6
0ADD
0A5E
0AF6
0B9F
0B4B
0A96
0AE4
0C1E
0C9C
0BA1
0A90
0ADA
0BC4
0B90
0A3E
09AC
0AC1
0C01
0BC0
0AB8
0AEE
0C41
0BC7
0750
0067
FAD5
F8CB
F97A
FAE2
FBA4
FB19
F90D
F625
F3F3
F3A8
F4B4
F56B
F4FE
F435
F3FB
F428
F41C
F3F1
F424
F488
F471
F3E3
F3B4
F449
F4E5
F4BA
F426
F429
F4C8
F502
F470
F415
F4E1
F632
F6AC
F625
F5C6
F628
F66D
F5CB
F52C
F640
F90E
FBA1
FC5E
FBD9
FBAA
FC2A
FC58
FBAE
FAFC
FB25
FBD9
FC2F
FC0F
FC2C
FCB7
FCFE
FC8A
FBDC
FBA2
FBC9
FBEF
FC2A
FC9A
FC9C
FB98
FAAE
FC6F
01D9
084F
0BD9
0B86
0A3F
0AD6
0C70
0C08
08B1
04DA
0335
03B9
045F
0401
0360
0382
0433
0495
046A
0425
0416
041F
041F
040A
03CC
0375
0363
03DD
0487
04B0
0440
03E4
0421
0487
044D
0388
0328
0398
0418
03DC
0348
0381
0519
0791
0A00
0BA9
0C2D
0BAB
0AD0
0A67
0AA6
0B1A
0B66
0BC9
0C78
0CDE
0C34
0ADD
0A33
0AC8
0BA6
0BCF
0B97
0BBE
0BE2
0B1A
09E4
0A0D
0BFC
0D16
0A3B
03AD
FD41
FA4F
FA92
FB80
FB7C
FAA0
F940
F74C
F531
F40D
F45A
F51B
F513
F45A
F407
F472
F4CB
F489
F452
F4D2
F585
F577
F4B0
F411
F409
F446
F48A
F503
F59B
F5A9
F4E5
F41A
F437
F4DA
F4C9
F3E1
F375
F452
F562
F54C
F4B2
F57E
F829
FAE3
FBE4
FB9C
FBCA
FCEF
FDCE
FD6D
FC69
FBE0
FBE4
FBD7
FBA8
FBC1
FC0D
FC03
FBAE
FBCA
FC85
FCEA
FC3A
FB3C
FB3C
FBFA
FBDA
FAA7
FAE3
FF08
05F4
0B7F
0CEB
0BAD
0B1C
0C24
0C7F
0A1E
0610
034E
032F
0433
043D
031E
025D
0304
045D
04ED
043B
0335
02FF
03B6
0486
04B0
0438
03A6
036D
03A0
040C
046A
0470
0406
0375
0340
039D
0427
044B
03FA
039E
0370
0358
0388
04C6
077C
0AAF
0C8E
0C58
0B3C
0AF6
0BCB
0C87
0C54
0BBE
0B9D
0BCC
0B9A
0B15
0B02
0B98
0C16
0BE6
0B87
0BA2
0BC2
0AF4
09A1
098C
0B59
0CE2
0B25
05AC
FF3C
FB15
FA28
FB25
FC54
FCA9
FB8F
F8FF
F601
F437
F438
F4DC
F4C1
F3FF
F3B7
F440
F4BF
F48D
F437
F480
F518
F50E
F454
F3E9
F456
F4EB
F4E9
F4B2
F516
F5EB
F641
F5CD
F54A
F53B
F524
F47B
F3C9
F408
F50F
F59F
F54C
F564
F735
FA1E
FC23
FC44
FB69
FAF7
FB40
FBA1
FBAB
FB8E
FB94
FBD5
FC59
FD03
FD4A
FCAB
FB95
FB3F
FC17
FCEF
FC84
FB52
FAF5
FBBD
FC21
FB44
FB14
FE68
0510
0B2D
0D42
0C04
0AF4
0BC7
0C91
0AC3
06B9
034A
026F
036E
0461
047C
0439
03FB
0399
0313
02EE
0373
0420
044D
040A
03F7
044F
0490
043D
0398
034B
0390
0405
0447
0456
044B
0411
03AA
0375
03D0
046A
046A
0388
02D6
03F7
0740
0AFC
0CEC
0C6F
0AFB
0A61
0AF5
0BAD
0BC4
0B98
0BCB
0C1D
0BCD
0AE8
0A6F
0AF1
0BA6
0B7D
0AAC
0A6D
0B2F
0BE5
0B95
0AF1
0B52
0C4A
0B53
06AE
FFDF
FA83
F8CB
F9C2
FAFD
FB1C
FA4C
F909
F76A
F5A3
F469
F441
F4CF
F540
F536
F4E9
F49C
F45A
F439
F457
F493
F494
F44A
F42B
F49E
F552
F58F
F529
F4C3
F4E9
F563
F5A3
F58C
F562
F53F
F509
F4DD
F4F9
F531
F4EE
F42B
F412
F5EF
F970
FC8E
FD92
FCC9
FBE1
FBE9
FC74
FC95
FC1E
FBA1
FBA1
FC1C
FCB0
FCE2
FC5B
FB4F
FA91
FAD4
FBBC
FC22
FB94
FAFA
FB3E
FBCE
FB7A
FAC8
FC49
0198
089A
0D0C
0D13
0B29
0ACF
0C32
0C51
093F
04CE
026A
0318
04C5
0527
043A
036F
0373
03AD
038A
034B
0360
03A6
03BA
03A3
03BD
041B
0467
0463
043A
0428
0424
0401
03C5
0383
032C
02C6
02C0
0391
04EC
05BB
054C
0456
0481
06AF
09DF
0C17
0C59
0B7B
0AFD
0B58
0BD1
0BB8
0B62
0B89
0C18
0C26
0B57
0AA2
0B17
0C3E
0C91
0B9F
0AB8
0B07
0BCC
0B83
0A5D
0A42
0BC9
0C65
08F0
01CF
FB26
F899
F9D5
FBDB
FC87
FBC6
FA1A
F7A9
F501
F37B
F3CD
F4DC
F4EE
F3E8
F351
F40C
F526
F562
F4F0
F4BC
F4D5
F491
F405
F420
F51F
F5F3
F5A7
F4D3
F4C7
F5AC
F65C
F620
F59B
F58D
F5B7
F58D
F550
F583
F5C9
F567
F4C9
F56A
F7E0
FAC5
FC40
FC27
FBDD
FC34
FC89
FC26
FB91
FBAA
FC48
FC87
FC2A
FBBF
FB9B
FB73
FB1B
FAE4
FB0A
FB3B
FB34
FB60
FC1B
FCA7
FC00
FAF1
FC22
0103
0762
0B5A
0B91
0A76
0AEC
0CAF
0CF2
0A16
05C5
02FF
02DF
03F4
0473
0413
03B1
03CE
040A
03DA
0359
031D
0381
0439
04A6
0477
03DE
034F
0325
0365
03B0
037F
02B9
0202
022C
033A
0438
0454
03DC
03CF
0469
04BA
041A
0385
04C3
0819
0B94
0D18
0C9B
0BC7
0BC9
0C46
0C68
0C33
0C3A
0C7F
0C56
0B70
0A74
0A33
0A9C
0AFE
0B1D
0B66
0C0D
0C6D
0BD7
0ABC
0A7E
0B98
0C4D
09DE
03B4
FCD2
F947
FA08
FBFA
FB78
F831
F4E5
F3CD
F458
F4B2
F473
F49C
F578
F5DB
F4FB
F3C7
F3A3
F47F
F527
F50F
F4DC
F525
F59B
F59F
F526
F48C
F3F6
F370
F36D
F461
F5CA
F681
F62D
F5A1
F56C
F518
F475
F4B6
F70A
FA89
FCC2
FC87
FB3D
FADF
FB8D
FBE9
FB67
FAE1
FAF3
FAFE
FA83
FA3C
FAED
FC05
FC75
FC47
FC4C
FC99
FC71
FBC9
FB99
FC32
FC5A
FB30
FA68
FCEB
0306
097D
0D25
0DF3
0D89
0C17
08B0
041D
0134
01A8
03CD
04A2
0374
0242
02AB
03F4
048D
0453
0443
04A9
04D4
0461
03D3
03CE
0456
04F0
0515
0488
038D
02E1
0318
03E4
044F
03EB
0376
03C4
0462
0436
038A
0443
075E
0B20
0CD9
0C14
0ADF
0B15
0C57
0D10
0CA4
0BDB
0B76
0B4F
0B0D
0AEC
0B44
0BC6
0BDC
0B93
0B7A
0BA5
0B7B
0AAB
09ED
0A5C
0BF8
0CEC
0AD1
0518
FE37
F9CF
F958
FAD7
FB17
F8F8
F625
F4AA
F4A6
F4CE
F48F
F48F
F513
F53B
F46E
F388
F3C0
F4DC
F582
F512
F460
F463
F4FF
F57A
F598
F5AE
F5CA
F59B
F528
F4F7
F52F
F550
F51E
F511
F555
F541
F482
F427
F582
F843
FA9C
FB6A
FB5C
FBA5
FC3B
FC47
FBCC
FBB4
FC37
FC6B
FBE9
FB94
FC04
FC61
FBC2
FAE0
FB12
FC16
FC5A
FB7D
FB11
FC15
FCFE
FBD6
F9D9
FAE5
00B8
0858
0D59
0E6D
0D68
0BD6
098C
067A
03F8
035A
0424
04A5
0417
033B
02F9
0345
03B0
0422
047E
0444
035C
02A2
02E2
03BB
042E
03FF
03CB
03F5
0436
044E
0466
0495
047C
03E7
0361
0386
03EA
03BA
0379
04EA
088B
0C44
0D99
0C9B
0B78
0B82
0BE1
0B67
0A85
0A8F
0BAC
0C80
0C11
0B02
0A78
0A8F
0A99
0A78
0AC1
0B9F
0C4C
0C01
0B05
0A7F
0B16
0BB3
0A08
04EB
FE40
F9C7
F983
FB87
FBF8
F93E
F586
F3DA
F487
F547
F4A1
F392
F38F
F444
F45C
F3B0
F36C
F432
F543
F5AC
F570
F532
F534
F546
F562
F5B6
F609
F5DB
F53E
F4E3
F50E
F533
F503
F50B
F5A1
F611
F5A0
F509
F5CE
F824
FA7F
FB71
FB4D
FB51
FBBE
FBC5
FB32
FAF3
FB97
FC60
FC74
FC19
FBF9
FBF8
FBB1
FB81
FBFC
FCA2
FC51
FB26
FACA
FC0B
FD44
FC77
FAC3
FBD5
015C
087E
0CF8
0DA8
0C9B
0B80
09E1
070C
0401
0284
02E5
03D4
0434
0432
0460
04A0
0487
0436
0418
042F
043E
0448
045E
0438
03A1
0307
030E
03A7
041E
0415
03EA
03FD
040F
03C1
0364
038E
0401
03F0
039F
04A5
07D4
0B8E
0D47
0C6A
0AD6
0A89
0B8D
0C82
0C82
0BEA
0B81
0B7F
0BA5
0BC2
0BCB
0BAC
0B66
0B30
0B32
0B38
0AED
0A44
0991
095F
0A0F
0B07
0A62
0669
FFF8
FA9D
F958
FB3C
FC42
F9DA
F5BF
F390
F43F
F55D
F4CB
F36A
F33E
F466
F540
F4EF
F431
F3D8
F3B9
F382
F3A2
F495
F5D5
F656
F5F8
F597
F59B
F568
F4AB
F427
F491
F561
F5A9
F56F
F54E
F541
F4D8
F488
F5A3
F888
FBA4
FCFD
FC6B
FB79
FB35
FB33
FAE5
FABE
FB45
FBF8
FC04
FB8A
FB3A
FB35
FB23
FB23
FBB1
FC8D
FCC9
FC3E
FC10
FCF5
FD9F
FC6B
FA79
FB60
00DC
082C
0CF5
0DDD
0CE4
0BDF
0A6E
07BF
04C3
0352
03BF
0488
047E
041E
0457
04EC
04F3
044D
03B6
039A
03B5
03BC
03C3
03DE
03E7
03D3
03DB
0434
04B6
04FA
04BC
040E
033F
02C0
02F5
03AD
03FC
0349
0289
03A8
0727
0B05
0CBF
0C07
0AC9
0AB3
0B90
0C32
0C27
0BF4
0BF7
0BE9
0B99
0B71
0BC3
0C10
0B9E
0A90
09D9
0A13
0ACC
0B18
0AB3
0A64
0B0C
0C18
0B42
06A3
FF53
F94B
F7D1
FA0D
FBD8
FA27
F623
F35B
F37D
F4E5
F54F
F48D
F3FD
F451
F4FF
F567
F574
F540
F4D6
F486
F4BF
F561
F5A3
F520
F491
F4D5
F589
F578
F483
F3FC
F4B4
F5C0
F5ED
F58E
F5BE
F66A
F669
F58C
F55D
F729
FA11
FBF8
FC0B
FB6B
FB4A
FB7F
FB71
FB59
FBB8
FC41
FC3F
FBB8
FB54
FB51
FB5F
FB62
FBAA
FC37
FC7D
FC47
FC3D
FCCE
FD0E
FBDA
FA34
FB0B
FFDC
0681
0B64
0D27
0D15
0C7B
0B14
086C
0582
03FC
0426
04B1
048C
040C
03F7
043F
0456
0438
0447
046F
043B
03AC
034C
0374
03D8
040E
0409
0404
0414
0421
0420
0410
03DB
0378
0338
0370
03CB
03A2
032B
03C7
065D
09DE
0C1F
0C28
0B1F
0ABD
0B66
0C1F
0C0B
0B68
0B02
0B2E
0BA4
0C05
0C30
0C0F
0B92
0AE2
0A6A
0A7F
0B07
0B74
0B49
0ABE
0AAA
0B3D
0AF2
07B2
0173
FB3F
F8A0
F9F2
FBE1
FAFF
F756
F3E2
F2DF
F3B7
F485
F48C
F45A
F464
F484
F498
F4C6
F4F9
F4D5
F460
F433
F4B0
F556
F564
F4EA
F4AB
F4E8
F504
F4A6
F463
F4DB
F5BD
F643
F646
F617
F5B3
F4E2
F42E
F4D0
F740
FA46
FC20
FC59
FBF7
FBD5
FBBB
FB4D
FAF6
FB36
FBB8
FBD0
FB8D
FB8F
FC01
FC5E
FC57
FC33
FC2C
FC04
FBB0
FBD3
FCBF
FD53
FC24
FA11
FA53
FEFD
0621
0B9D
0D65
0CE1
0C1E
0B26
08DA
0598
036E
0398
04EB
0567
049F
03BF
03AB
0408
042B
0414
042C
0482
04B7
048D
043C
0425
046A
04CD
04EA
0488
03CB
0327
0300
033D
0378
0396
03D6
0432
042B
03B2
03D7
05DD
096F
0C62
0CD3
0B44
0A0B
0A99
0BFA
0C5B
0B70
0AA6
0B06
0BDF
0BF1
0B37
0AC7
0B1D
0B67
0AE0
0A13
0A17
0AD4
0B17
0A7D
0A43
0B4A
0BE8
091A
025D
FB32
F7E0
F8FF
FB2A
FAF5
F84E
F5A5
F4A5
F4CA
F4CF
F466
F409
F3F5
F401
F41B
F44F
F46F
F448
F41E
F46D
F531
F5CA
F5CD
F58A
F577
F563
F4D2
F3F9
F3B5
F455
F520
F564
F566
F5A2
F5C3
F51C
F414
F42F
F64D
F96C
FBB0
FC57
FC2A
FC17
FC2F
FC25
FC08
FC09
FBFC
FBB8
FB90
FBD6
FC2B
FBEF
FB52
FB42
FC06
FCAD
FC54
FB96
FBB3
FC8E
FCA2
FB87
FB5C
FE9A
04D8
0ADC
0DE2
0DF5
0CBE
0B0C
088D
0579
033A
02DF
03B6
0439
03EB
0394
03CA
0429
041F
03E3
0411
04AF
0519
04EC
047D
0445
0437
0409
03D7
0407
049A
04F7
049E
03CA
0336
034C
03BE
03E3
0374
02F7
0373
058F
08CD
0B9B
0C92
0BC6
0AB4
0AB9
0BB7
0C8D
0C93
0C3C
0C24
0C1E
0BA4
0AE3
0A9E
0B09
0B60
0B0C
0A92
0ABD
0B45
0B1C
0A42
0A34
0BB1
0CB3
09FA
0312
FBBD
F872
F9BD
FBF3
FB72
F83D
F51F
F411
F479
F4BC
F45C
F405
F426
F461
F459
F449
F499
F535
F5A9
F5B4
F575
F51B
F4B1
F44D
F428
F465
F4D4
F520
F522
F4F2
F4B8
F48C
F47E
F49B
F4E1
F560
F65D
F813
FA3B
FBFC
FC9E
FC48
FBD5
FBDF
FC31
FC48
FC18
FBF9
FBFB
FBC7
FB48
FB07
FB6D
FC03
FBF2
FB4C
FB21
FBF4
FCB8
FC16
FAAB
FB0A
FEF1
0502
09FC
0C17
0C54
0C5A
0C05
09FF
0646
02F5
020E
033C
0466
0437
0344
02CE
031C
038D
03B5
03BC
03D0
03D7
03C9
03E0
0437
047D
0462
0414
03F9
0406
03D2
035D
033F
03BD
041B
0373
022B
01F0
03EC
075E
0A4D
0B87
0B91
0B9C
0C0C
0C4F
0BF0
0B4B
0B0E
0B62
0BD6
0BF7
0BC2
0B7B
0B5E
0B7F
0BD3
0C1C
0BF7
0B40
0A8A
0AB6
0BAD
0BAE
08A4
0299
FC6F
F980
FA61
FC4C
FBFF
F8F2
F56A
F3BA
F405
F4D1
F507
F4CE
F4B4
F4C7
F4BD
F49B
F4BC
F547
F5E8
F635
F616
F5B9
F543
F4BB
F437
F3EC
F400
F461
F4CB
F4FA
F4E9
F4D7
F4F3
F514
F4F3
F4CD
F581
F7B0
FAB6
FCEE
FD45
FC56
FB9F
FBC7
FC17
FBCC
FB48
FB7B
FC6C
FD1E
FCEC
FC5B
FC28
FC14
FB5C
FA42
FA2E
FBB7
FD45
FCC3
FAA3
FA39
FE3A
055F
0B63
0D72
0CA5
0BDA
0BDC
0AE3
07AF
03D2
0205
02D3
041E
03F6
02D9
0289
0383
0493
04A2
0408
03B0
03BD
03A9
0359
0335
0356
0346
02E8
02DA
0383
043F
0430
0395
037D
0433
04B5
042E
036D
0415
0694
0985
0B56
0BCD
0BA9
0B6F
0B29
0AF9
0B1E
0B72
0B7A
0B2C
0B0D
0B53
0B66
0AC4
0A13
0A74
0BC2
0C68
0B86
0A73
0B15
0CE9
0CD5
0883
0158
FB5F
F95D
FA6F
FB91
FAD1
F89B
F66A
F510
F46D
F42F
F447
F4A5
F4FE
F502
F4C4
F4AB
F4F2
F553
F54F
F4D0
F44C
F446
F4C9
F56C
F5D4
F600
F61B
F613
F5A4
F4CB
F408
F3F3
F48C
F524
F511
F493
F4C2
F686
F975
FBFA
FCD1
FC3A
FB8A
FB96
FBF9
FBF8
FB9F
FB8B
FBD6
FBE7
FB81
FB57
FBFA
FCBC
FC75
FB66
FB2E
FC72
FD7F
FC73
FA64
FAF1
0016
075D
0C42
0D09
0BFC
0BD7
0C48
0B04
077B
03F2
02CA
03CD
04D7
0499
03B8
035F
03AB
03E9
03DA
03E1
0432
0466
042D
03D3
03D6
0423
0435
03DE
0398
03D2
043E
0420
0356
02AA
02DF
03AC
0415
03CC
03D1
055D
085A
0B39
0C78
0C0F
0B40
0B21
0BB0
0C38
0C40
0BE3
0B76
0B23
0AE0
0A93
0A48
0A43
0AB9
0B65
0B9A
0B0C
0A68
0AA8
0B85
0B02
0751
0131
FBC7
F9B0
FA78
FB6C
FA94
F85C
F663
F578
F527
F4DC
F49E
F4A2
F4BB
F498
F458
F463
F4C7
F518
F4F8
F488
F436
F441
F493
F4F0
F52D
F551
F57E
F5C4
F5F1
F5B1
F505
F472
F482
F4FD
F514
F486
F44C
F5A9
F882
FB32
FC35
FBB6
FB27
FB76
FC29
FC58
FBF1
FB98
FB95
FB85
FB3E
FB4D
FC19
FCF4
FCCF
FBC7
FB42
FC0C
FCF5
FC52
FAC2
FB4D
0002
0707
0C28
0D4B
0C4E
0C0C
0C99
0B9B
080D
041D
02A2
03A7
04A6
03F3
0291
025B
0378
0483
04B0
048B
04A9
04B4
0444
03EB
0479
0585
05A6
0457
02DD
02BA
03C3
0485
0446
03C3
03D7
0424
03BB
02C3
02B0
04AF
0831
0B5A
0CBE
0C6F
0B91
0B3D
0BB6
0C71
0CB6
0C4E
0BAB
0B4E
0B38
0B0A
0AAC
0A86
0AE2
0B56
0B37
0AA1
0A93
0B98
0C80
0B0D
0639
FFA9
FA83
F8C4
F9BA
FB09
FAED
F965
F778
F5E6
F4CB
F428
F426
F4AF
F52D
F515
F492
F45E
F4D6
F578
F589
F4F9
F46F
F465
F4A5
F4B3
F47E
F45D
F497
F517
F590
F5C0
F598
F552
F54D
F5A1
F5DF
F595
F522
F5B8
F805
FB08
FCCF
FC96
FB96
FB68
FC22
FC92
FC0C
FB39
FAF1
FB23
FB4A
FB7E
FC36
FD13
FD07
FBE8
FB11
FB9A
FCA7
FC92
FBAB
FC94
0114
0764
0BC2
0C8E
0BC2
0BEC
0CC8
0BF2
0872
0453
0249
02A8
0389
036A
02B8
02AC
0375
0437
0463
0442
0430
0403
038B
032F
037C
043C
0498
0436
03C5
0409
04BB
04D7
0405
0320
031D
03BA
03E0
032F
02BD
03F7
06F6
0A45
0C3F
0C71
0BB2
0B20
0B37
0BAC
0BF7
0BDE
0B9D
0B89
0BAB
0BBA
0B92
0B6F
0B92
0BAC
0B27
0A1A
0994
0A5C
0B75
0A85
0633
FFFF
FB2D
F9CB
FAFE
FC43
FBEE
FA24
F7E2
F5CE
F431
F363
F3AA
F4A8
F57A
F592
F530
F4E5
F4E2
F4F2
F4F5
F500
F512
F501
F4CE
F4C5
F510
F562
F558
F50D
F4FA
F535
F547
F4EC
F498
F4DB
F579
F5A9
F55E
F5AA
F785
FA65
FCA4
FD44
FCD1
FC6F
FC81
FCA3
FC98
FC8A
FC7D
FC24
FB8B
FB53
FBD9
FC6D
FC21
FB44
FB34
FC61
FD51
FC8C
FB3B
FC8F
01F5
08C2
0CB8
0C9A
0B2F
0B75
0CE4
0C86
0920
04F8
0308
038E
044E
03C1
02BC
02B7
0397
040D
039A
0329
0382
041D
0402
034A
02F9
0373
03E8
038E
02D4
02C1
037A
0405
03AD
02F4
02DD
0387
0405
03A6
0304
0391
0607
0982
0C33
0CEE
0C25
0B54
0B72
0C0F
0C18
0B58
0AB7
0AEC
0B70
0B40
0A6C
0A27
0B17
0C32
0C14
0B12
0AF6
0C5B
0D2C
0AAF
04CD
FE84
FAF6
FA9E
FB9A
FC15
FB9B
FA75
F8B7
F687
F4A4
F3EA
F445
F4B3
F475
F3D9
F3AC
F427
F4C6
F50B
F504
F50C
F53D
F564
F568
F56C
F588
F597
F568
F50E
F4C8
F4B1
F4A0
F462
F407
F3D3
F3E4
F41D
F482
F57B
F769
F9F7
FC12
FCD7
FC69
FBBE
FBA2
FC13
FC92
FCC3
FC9C
FC39
FBC9
FB97
FBC0
FBE9
FBAD
FB4C
FB81
FC47
FC81
FB81
FABB
FCDF
02B4
0980
0D66
0D67
0C1B
0C3C
0D5F
0CDE
098C
0556
0309
0345
044F
0477
03E2
03BC
0462
04FE
04C8
040F
03B0
03EC
042E
03ED
0369
034E
03C1
0422
03DC
0337
0303
0378
03F6
03E8
039B
03C2
046B
04E6
04D6
04E9
062A
08A8
0B2F
0C6F
0C31
0B4C
0AA4
0A7D
0A96
0AA4
0AA6
0AD2
0B38
0B8A
0B6E
0B05
0AD9
0B2E
0BA1
0BBF
0BAF
0BD2
0BA0
099D
0510
FF82
FBB6
FAE0
FB9D
FBD8
FAFC
F9C0
F87B
F6C7
F4BC
F376
F3C6
F4F0
F573
F4E1
F42E
F41C
F453
F445
F445
F4E4
F5D3
F634
F5E0
F591
F5B7
F5CD
F53F
F467
F410
F446
F45D
F422
F43F
F4FE
F582
F4E6
F3D0
F3FC
F637
F963
FBBD
FC93
FC78
FC2C
FBEC
FBCC
FC19
FCF3
FDD7
FE06
FD68
FCAA
FC74
FCD1
FD65
FDF6
FE6C
FE76
FDA1
FC2B
FB9B
FDDD
0332
0939
0CBC
0CC0
0B5F
0B46
0CA9
0D4D
0B76
080D
057D
04E4
053E
0533
04BD
04A0
04FB
0530
04E2
046E
0451
0497
04F8
052E
0507
047C
03E3
03DC
04A4
0594
05BB
04FE
0420
03AF
0377
034C
0393
0478
0526
04BC
03D3
0440
06E2
0A51
0C46
0C0E
0AF9
0A85
0AD9
0B4C
0B89
0B9E
0B73
0AF5
0A7E
0A88
0AF0
0B29
0B06
0AE5
0AF5
0AE1
0A8B
0A8A
0B3E
0B95
09BA
055C
0085
FD96
FCE8
FD0E
FCEC
FC96
FC3B
FB3F
F911
F65B
F4A4
F49C
F55E
F5A1
F538
F503
F595
F67E
F6EA
F696
F606
F5E4
F64B
F6BA
F6BE
F68D
F6A6
F6FC
F6DF
F5FE
F518
F52E
F625
F6CB
F665
F5AB
F5BA
F665
F67A
F5CF
F5F7
F848
FBCA
FE19
FE28
FD4B
FD3F
FE04
FE40
FD5E
FC63
FC76
FD54
FDC8
FD54
FCAD
FC91
FCCD
FCC9
FC84
FC92
FD0B
FD2B
FC6A
FBD7
FD9A
028C
08A7
0C95
0CF8
0B9D
0B1F
0BE9
0C24
0A67
0797
05B0
0558
0576
04F9
0427
03D4
0414
0455
044B
0423
0409
0400
0420
0482
04E9
04E0
0461
0400
0434
04B5
04EC
04CA
049D
0442
0358
0260
0299
0431
0578
04D9
032B
02F4
055F
08DF
0B25
0BB4
0BB1
0BDB
0BCF
0B59
0B28
0B9C
0BEF
0B61
0A7B
0A45
0AB4
0AE5
0AA5
0AA7
0B17
0B19
0A4D
09E6
0AFF
0C3E
0AB1
0589
FF9B
FC4B
FBF1
FC65
FC49
FC23
FC4A
FB89
F8D2
F551
F38C
F46A
F629
F6AC
F5E0
F539
F576
F5FC
F612
F5DF
F5EF
F65A
F6BB
F6B4
F649
F5CE
F59C
F5CA
F626
F661
F664
F65B
F66E
F67F
F663
F641
F666
F6B2
F6B7
F694
F72E
F91C
FB94
FD0A
FCDD
FBF8
FBAC
FC44
FCFF
FD2F
FCF6
FCD8
FCEF
FCEB
FCA7
FC62
FC52
FC59
FC3F
FC27
FC7B
FD45
FDC1
FD19
FBE5
FC72
0098
0721
0C3F
0D4C
0B90
0A8B
0BB5
0CE7
0B6E
07AC
0492
03EA
0475
042E
0313
02AE
0392
0491
047F
03B0
034E
03D1
04A4
050F
04F3
049D
0449
0414
0405
03FF
03E2
03DF
043A
049C
0439
02FC
01FB
0234
0336
03C4
03A5
0418
062B
0933
0B6E
0BED
0B50
0AA5
0A57
0A60
0AC6
0B5C
0B9D
0B50
0AE9
0AD3
0AC4
0A5C
0A0A
0A81
0B68
0B7C
0A6F
09BA
0A98
0BA8
0A05
04F4
FF41
FC24
FBD3
FC30
FBFD
FBD2
FC0F
FB85
F921
F5F8
F469
F531
F693
F6A6
F5A2
F514
F594
F633
F60A
F561
F525
F5B5
F69B
F711
F6BB
F5EF
F569
F5A2
F655
F6C8
F6A3
F65D
F693
F719
F72F
F69B
F606
F5FC
F629
F627
F690
F860
FB4D
FD88
FD9F
FC3A
FB58
FBFD
FD31
FD7E
FCC9
FC29
FC3F
FC88
FC6C
FC31
FC6A
FCDB
FCAD
FBC5
FB3A
FBE9
FCFE
FCD7
FB8D
FBBF
FFCC
0684
0BC3
0CBB
0AE0
09D1
0AF8
0C35
0AF1
0766
0425
02F9
035C
03DE
0403
0425
0463
0470
0438
03F2
03BF
03A5
03C4
0425
0459
03E0
030B
02E8
03DE
04DC
04A1
0391
033B
040D
04A1
03EB
02E9
031F
0428
0434
02ED
0269
0496
0893
0B9D
0C4B
0BB3
0B58
0B4C
0AE9
0A5A
0A4A
0A9F
0AA8
0A4C
0A2C
0A89
0ADC
0ABF
0A96
0AC9
0AEE
0A7F
0A10
0AAD
0BD2
0B28
0727
0141
FC89
FA99
FA9C
FB12
FB60
FB5F
FA86
F86C
F5D2
F43B
F444
F4F9
F539
F512
F54B
F603
F682
F647
F5A3
F532
F53B
F59C
F610
F655
F638
F5C8
F560
F560
F5CA
F648
F697
F6AE
F68C
F633
F5DE
F5ED
F651
F676
F621
F61F
F788
FA47
FCDF
FDE1
FD64
FCB1
FCB4
FD1F
FD2B
FCB9
FC57
FC64
FCA9
FCD8
FCFA
FD28
FD27
FCAA
FBEF
FBB4
FC40
FCC5
FC37
FB0D
FB83
FF71
05CE
0B27
0CE6
0BD5
0AD8
0B7A
0C68
0B7B
0877
052D
033C
02A9
02B8
0324
03E1
0458
03DE
02C0
022C
02C0
03C6
0423
03B5
0355
039B
0429
0448
03D9
035E
035E
03ED
04AB
04FD
0493
03E1
03B9
0439
0476
03B0
029D
02EA
0557
08C2
0B4F
0C3F
0C2A
0BC9
0B41
0AAE
0A7F
0AD5
0B24
0AFA
0AB0
0ABE
0AD5
0A5C
09A1
09AE
0AAD
0B59
0AC1
09E8
0A7B
0BE5
0B2E
067F
FFD3
FB14
FA09
FB25
FC1B
FC41
FBFF
FB22
F8FC
F5FB
F3D5
F39E
F47B
F4DB
F476
F443
F4D5
F590
F5AF
F552
F527
F571
F5D8
F612
F646
F69D
F6D4
F689
F5D0
F531
F518
F561
F590
F54F
F4C3
F46F
F4AD
F53B
F586
F574
F5C9
F751
F9C6
FBD6
FC82
FC32
FC1F
FCC8
FD71
FD55
FCC3
FC9D
FCFB
FD08
FC4F
FB88
FB9D
FC4C
FC78
FBCE
FB55
FBE4
FCAE
FC3F
FAF2
FB56
FF6D
05EB
0B1A
0CA7
0BC4
0B46
0C44
0D3D
0C4E
095D
05EE
0382
02A2
0313
0432
0516
04F7
03F1
02EE
029D
02BD
02BA
02A5
02F5
03A2
0405
03C8
036D
0396
0420
0479
0492
04D8
053E
0511
0421
0355
037D
0413
03E9
02FB
02C2
0472
0771
0A00
0B15
0B0B
0AB7
0A7F
0A7A
0AB5
0AFC
0AE6
0A85
0A91
0B5A
0C0C
0BAA
0A8F
0A13
0A9C
0AF1
0A09
08DC
092A
0AA4
0A8A
06DF
00F6
FC14
FA07
FA0C
FAA5
FB2A
FB5E
FA96
F864
F5AC
F40C
F403
F473
F44E
F3EF
F446
F53B
F5CF
F590
F519
F50E
F53F
F537
F50C
F535
F5AE
F5E5
F597
F539
F548
F598
F5A4
F559
F519
F528
F56F
F5C2
F601
F604
F5CB
F5DC
F700
F94B
FBA5
FCBD
FC87
FC37
FCB8
FD8E
FDA7
FCDB
FC08
FBDA
FC1A
FC4E
FC79
FCCF
FD03
FC98
FBD3
FBB1
FC81
FD1E
FC4D
FACC
FB2C
FF25
0565
0A8B
0C59
0B94
0AB3
0B23
0C20
0BF2
09DC
06B6
040C
02E3
032B
03F8
044C
03D4
0311
02C7
032C
03BE
03E6
03A7
038C
03F5
049B
04E0
046A
0384
02D3
02D8
038A
045F
04B2
0451
03AD
0371
03D0
0452
0466
0415
040E
04FC
06E3
0912
0AAD
0B41
0B08
0AB1
0AD6
0B72
0BDE
0B7C
0A77
09AD
09D4
0ABB
0B95
0BD0
0B78
0ADB
0A2B
099F
09A5
0A76
0B56
0ABA
0791
0287
FDB9
FB06
FAA8
FB63
FBD1
FB5A
FA28
F896
F6EC
F57F
F4B0
F4A0
F4FB
F53D
F522
F4CE
F48D
F485
F4A8
F4DA
F503
F50C
F4E6
F4A3
F47A
F499
F4F8
F567
F5BD
F5F0
F5FA
F5CB
F567
F503
F4D7
F4DB
F4C0
F44B
F3C7
F3FC
F58E
F843
FAF5
FC67
FC54
FBAE
FBB1
FCA7
FDA7
FDAD
FCB6
FBB7
FB78
FBE0
FC5F
FCAE
FCD5
FCBA
FC1E
FB29
FA87
FAA9
FB37
FBB9
FCB0
FF56
03E9
08C3
0BAF
0C19
0B74
0B60
0BE3
0BA9
09C4
06B9
03E3
0247
0211
02BF
0382
03A8
0327
02A6
02C9
0377
0402
0401
03BF
03B3
03DC
03DB
038F
0349
0351
0390
03D1
040F
044E
0458
03F3
034D
02DC
02E6
0336
0367
0357
0353
03F5
05C6
08B5
0BBF
0D5C
0CCA
0AF4
09A3
09AD
0A55
0A9B
0A8C
0ADB
0B7A
0B83
0A8F
0973
0929
0980
09AA
09C2
0AB8
0C5A
0C7C
0914
02DC
FD05
FA1E
F9F3
FA9E
FAE5
FB04
FB82
FC40
FCC5
FCBD
FBD0
F99D
F683
F3F3
F345
F433
F529
F520
F4A4
F4C6
F58B
F608
F5CA
F563
F56E
F5B3
F5B5
F58B
F59F
F5E1
F5DD
F57E
F542
F579
F5D1
F5D5
F58F
F54C
F50C
F4AB
F477
F4E0
F589
F579
F4AA
F4B4
F711
FAFA
FDDE
FE24
FCBA
FBA7
FBAC
FBFD
FBE5
FBAD
FBBD
FBD7
FBBB
FBD6
FC90
FD62
FD66
FCAF
FC31
FC50
FC69
FC40
FD25
008D
05BD
0A08
0BAF
0B97
0B95
0BE9
0B88
0A58
09AD
0A3F
0AC3
0974
0680
03F9
0352
03E2
0432
03E5
039E
03A4
038B
032B
02FE
0357
03BA
037D
02A6
01E0
01A5
01E9
028C
0395
04C4
0563
0500
0405
0338
02D9
02A5
0299
031B
0430
04F5
0468
02B7
016F
022F
0525
08E8
0BAB
0C8C
0BF4
0B01
0A83
0A75
0A5E
0A18
09E8
09F5
09FF
09EC
0A1C
0AD6
0B8D
0B59
0A49
09A1
0A2F
0ABD
090A
0486
FF4E
FC12
FB6B
FBD9
FBE3
FB6D
FB1E
FB3B
FB81
FB97
FB1F
F9A3
F72A
F4D7
F421
F524
F647
F606
F4AD
F3B6
F3E1
F499
F520
F573
F5D1
F5FC
F58E
F4CD
F476
F4A9
F4C5
F481
F476
F528
F60E
F638
F59C
F514
F537
F5C8
F64B
F68A
F654
F558
F3F4
F3A6
F5C3
F989
FC73
FCF1
FC0D
FBD4
FCC0
FD9D
FD8A
FD07
FCCF
FCB5
FC40
FBCE
FC1A
FCF8
FD78
FD6B
FDA3
FE3C
FDFC
FC61
FB7B
FE21
0428
09D1
0BB1
0A4D
08F3
0987
0AEB
0B80
0B85
0C09
0C92
0B78
0860
0512
0367
034E
0374
0335
030D
0356
0391
034C
02F3
0322
03A5
03C9
037D
0364
03C7
0410
03A3
02C4
0247
0287
030B
0336
02FF
02CC
02E1
032F
0398
03F4
0400
0386
02BB
024E
02FC
0502
07D9
0A6C
0BC8
0BC1
0B00
0A4B
09E6
099E
095B
0950
098E
09BA
0987
094E
09A1
0A4A
0A62
09B8
096E
0A80
0BE4
0B13
06CF
00E1
FC87
FB43
FBCD
FC01
FB3B
FA71
FA9E
FBA0
FC79
FC23
FA3F
F778
F536
F488
F525
F5B4
F554
F488
F46E
F52D
F5CD
F591
F4DF
F486
F4A4
F4C1
F4B7
F4CB
F50D
F52F
F51A
F53E
F5DB
F66B
F634
F55A
F4C7
F4E7
F531
F516
F4DD
F4FF
F534
F4E4
F46F
F522
F7A7
FAEE
FD2F
FDBD
FD5D
FD07
FCF4
FCFC
FD23
FD55
FD30
FC9E
FC4C
FCD5
FDB9
FDD4
FCF1
FC1D
FC05
FBE4
FAE8
FA51
FCAB
027D
08D5
0C26
0C0C
0B22
0B6D
0C3D
0BFD
0ADE
0A6E
0AF4
0AB6
0852
04D8
0296
0260
02F7
0302
02A2
02AB
0334
0391
0370
033C
0347
034B
0305
02DC
034F
040A
042A
0380
02EF
034B
0433
048F
03FC
033C
0321
037D
0393
033F
0328
03A2
040E
03C5
035B
0443
06F9
0A12
0B8D
0B08
0A09
0A18
0AFD
0B64
0ACD
0A13
0A14
0A82
0A93
0A4B
0A59
0ACA
0AC0
09D6
0919
09C0
0B0F
0A84
069B
00CE
FC3A
FA8F
FAD9
FB33
FAE3
FA91
FAF8
FBF3
FCBC
FC97
FB30
F8CC
F657
F4DB
F493
F4BE
F49C
F456
F48D
F543
F5B7
F563
F4B6
F47B
F4DF
F569
F5B6
F5D4
F5D6
F5AF
F58D
F5CA
F644
F63B
F553
F45B
F463
F52F
F569
F483
F39E
F3F9
F4FD
F500
F3E5
F3B7
F615
F9EF
FCB5
FD5C
FD14
FD38
FDA2
FD87
FCFD
FCB6
FCA8
FC21
FB32
FAE9
FBAE
FC6C
FC1E
FB6A
FB91
FC44
FC0A
FB04
FBCF
0074
0727
0BAC
0C03
0A67
0A11
0B54
0C26
0B98
0B0B
0BA9
0C3C
0A9B
06A3
02A9
00EA
0166
0287
0320
0325
0300
02FA
0339
03B2
0401
03C6
0339
0308
0371
03E2
03BE
033E
0322
039C
040D
03F6
039E
037A
036E
0328
02F7
0385
04BF
0595
0521
03E0
0358
0497
0734
09D2
0B51
0B6D
0AAD
09ED
09CC
0A3D
0AAF
0AC1
0AA7
0AB4
0AD1
0AB1
0A67
0A55
0A7C
0A5D
09D2
0993
0A32
0AB1
08F1
0420
FE33
FA48
F9A8
FAD8
FB97
FB39
FACA
FB52
FC74
FCD4
FB78
F8A5
F5A9
F3E0
F3BA
F478
F4FA
F4E5
F4D4
F54F
F5FD
F61D
F59B
F524
F539
F58C
F588
F525
F4E0
F505
F564
F5C4
F621
F66B
F664
F619
F5EC
F5F9
F5BA
F4D8
F3FB
F424
F530
F5C7
F531
F4B2
F630
F9A1
FCC8
FDC7
FD20
FC96
FCDC
FD3B
FD18
FCD4
FCDC
FCE1
FC79
FC04
FC2C
FCBB
FCE6
FC9D
FCA1
FCF1
FC66
FABE
FA2C
FD53
03B7
0990
0BC1
0B14
0A8C
0B54
0BD1
0AC8
0995
0A18
0B92
0B37
07E6
03CF
01E8
02A3
03FC
0434
0371
02B4
0255
0214
0205
0277
033A
03B5
03B2
0396
03AC
03B6
0378
0337
0355
03A6
039F
0334
02FF
035F
03D9
03C7
0354
034C
03EE
0483
0454
03BA
03E5
0597
083F
0A72
0B32
0AB3
09EE
09AB
09F7
0A6F
0AD0
0B28
0B73
0B67
0AD7
0A29
09F2
0A16
09E0
0928
08E5
09EA
0B31
0A42
05D3
FFB7
FB6B
FABC
FC40
FD44
FCA8
FB6A
FAED
FB5B
FBC1
FB23
F949
F6D4
F4CC
F3F3
F436
F4BF
F4C1
F443
F3E7
F402
F442
F448
F432
F44A
F481
F4A3
F4D1
F556
F607
F641
F5AD
F4B8
F415
F3F6
F416
F45D
F4F2
F5AB
F606
F5E9
F5D3
F606
F5F9
F544
F4B7
F5BC
F880
FB68
FCD0
FCDB
FCEC
FD9E
FE29
FDC8
FCE9
FC65
FC59
FC63
FC85
FCF9
FD6B
FD34
FC81
FC58
FD01
FD4B
FC4D
FB7A
FD8B
0304
08F9
0C18
0C19
0B34
0ADE
0A88
098B
08CD
0966
0A88
0A0C
0733
03BE
01D5
01C6
0273
0321
03E0
048D
049B
03FD
0374
038E
03DD
03AB
0321
030D
039F
0413
03D0
0333
02DB
02C7
02AE
02B8
032C
03A9
036E
0289
020D
02C0
040F
04BD
047A
0435
04E2
0673
0842
09CC
0AB8
0ABB
0A00
095C
097B
0A05
0A21
09B9
0997
0A25
0AAD
0A5C
098B
0950
09E4
0A6A
0A70
0A98
0B21
0A9E
0759
01D2
FCD0
FA9E
FADF
FB84
FB5C
FAF5
FB3E
FC16
FC97
FC18
FA87
F83E
F5FE
F4B9
F4BB
F542
F556
F4E4
F4A1
F4E1
F536
F53B
F53A
F591
F5E4
F594
F4E9
F4DB
F596
F60D
F585
F4B2
F49D
F4FE
F4BB
F3C1
F35E
F45A
F5AF
F5D5
F4CB
F3EB
F3EF
F442
F495
F5E0
F8D8
FC4B
FE13
FD8A
FC0F
FB2E
FB17
FB35
FB68
FBEF
FC91
FCCC
FCBB
FCFE
FD85
FD6B
FC7F
FBEB
FC90
FD6F
FD0B
FC0C
FD21
01C7
07FA
0C18
0CA3
0B54
0A8F
0AE7
0B85
0BE2
0C36
0C9C
0CBE
0C42
0AF6
08AD
059C
02D6
01B2
0265
039E
03FD
039D
0394
0423
0459
039E
02B8
029A
02FB
02F3
0284
0289
0342
03DA
03B2
0352
0386
03FF
03C0
02D0
0273
0358
0475
0467
035C
02B0
02FF
0370
031B
0264
0297
0472
076D
0A3D
0BC4
0BAB
0A88
098F
0999
0A4A
0A94
0A1D
09A3
09CA
0A35
0A52
0A65
0AFA
0B9D
0B3C
09E8
093E
0A2F
0B04
08DF
035E
FD95
FACE
FB22
FC13
FBC6
FA9A
F9C7
F9BD
FA2C
FADB
FB9B
FBCF
FAC0
F89B
F681
F55A
F510
F51E
F551
F590
F583
F506
F4A1
F4DB
F558
F535
F464
F3EA
F47E
F572
F582
F48D
F3AF
F3B7
F43B
F47C
F47A
F48B
F48E
F446
F41E
F4C1
F5F2
F690
F605
F504
F488
F487
F46E
F49B
F643
F986
FC99
FD9C
FCB5
FBA1
FB7A
FBD1
FBD5
FB8F
FB94
FC11
FCA8
FD06
FD12
FCB2
FBEC
FB4E
FB7D
FC2B
FC43
FBB8
FC5E
0003
05DD
0AD3
0C92
0BC8
0AF6
0B85
0CA6
0CEA
0C1B
0B32
0AFA
0B3E
0B12
099C
06DE
0407
029F
0309
03FC
03EC
02D0
0206
0277
0374
03BE
0333
02C5
02FC
0359
0357
034C
03AC
041C
03F5
036D
0362
0408
0481
0410
0325
02BB
02FF
033F
032B
0353
0417
04B8
0443
0313
02B2
0436
070D
099D
0AC1
0AA1
0A3E
0A6B
0B1A
0B8E
0B2D
0A31
0977
0987
09FF
0A2C
0A08
0A1A
0A6C
0A6A
0A04
0A29
0B47
0BDD
0997
0432
FE61
FB38
FB13
FBC3
FB84
FAC4
FAB8
FB55
FB9F
FB58
FB44
FBA3
FB64
F982
F68D
F455
F3FC
F4EC
F5C2
F5CD
F562
F512
F50D
F526
F51B
F4CA
F456
F414
F424
F44B
F44C
F44B
F4A4
F555
F5DB
F5C1
F52D
F4B6
F4B2
F4FB
F544
F56F
F572
F544
F504
F4FB
F525
F523
F4E0
F517
F6B1
F98B
FC3F
FD6D
FD05
FC21
FBBA
FBDD
FC1C
FC49
FC7B
FCB9
FCEC
FCFF
FCD7
FC73
FC2E
FCA2
FDC0
FE63
FD6F
FBA4
FBAB
FF7D
05DE
0B17
0C94
0B46
0A1D
0AB0
0C00
0C4B
0B4A
0A48
0A68
0B49
0B5D
0974
05F0
0299
0131
01F8
037D
0414
037B
02E8
0362
047D
04FF
0468
036D
0300
035B
03FE
045D
0441
03BC
0310
02A7
02CF
035E
03D2
03E1
03C1
03AF
038E
0338
02F8
033B
03D9
040C
035A
0258
024E
0406
0704
09DF
0B5A
0B33
0A3C
09A1
09EF
0AA1
0AE3
0A9D
0A6F
0AA2
0AA5
0A00
0946
096B
0A4B
0AAE
0A12
09A6
0A8F
0B90
09C9
043A
FD9E
F9D0
F9D8
FB61
FBE7
FB41
FACE
FB19
FB7C
FB91
FBD3
FC60
FC2E
FA49
F770
F573
F516
F553
F4F1
F41F
F3F0
F4B2
F57A
F567
F4BE
F466
F4A5
F4EB
F4B3
F436
F3FC
F435
F49D
F4F1
F537
F587
F5C1
F597
F4FC
F454
F422
F482
F519
F58A
F5D5
F61F
F646
F5F8
F552
F536
F690
F93B
FBE8
FD47
FD2D
FC74
FC05
FC23
FC84
FCC7
FCB6
FC6C
FC40
FC74
FCD4
FCE4
FC96
FC8E
FD37
FDC3
FCEC
FB02
FA89
FDDB
0442
0A26
0C73
0B74
09EE
09ED
0B04
0BA7
0B4E
0AC3
0ACA
0B2B
0B0F
09DD
07B5
055B
03C8
0377
03FA
0456
0408
0383
038B
0423
0480
0419
034F
02E2
0307
0365
03AC
03D5
03D5
0394
033A
032D
0386
03C4
0361
02A4
0273
0333
0433
0481
0409
0383
0364
0351
02D1
0241
02B6
04DA
07F5
0A54
0AD6
0A01
096D
0A06
0B1D
0B57
0A6B
0982
09A3
0A4C
0A38
0952
08EB
09BC
0AAE
0A67
0972
0996
0AEF
0AE7
0720
00CA
FBCF
FA98
FBBD
FC59
FB94
FAD9
FB41
FC3D
FCDD
FD2A
FD72
FD05
FADA
F759
F46F
F376
F3C7
F3E9
F38E
F387
F430
F4D5
F4D6
F48E
F4B2
F53F
F598
F57A
F540
F534
F523
F4F1
F4FA
F576
F5E0
F58E
F4B0
F430
F476
F4E9
F4D7
F479
F498
F558
F5E5
F57D
F477
F3EC
F49C
F660
F890
FA87
FBD7
FC5B
FC50
FC3A
FC6F
FCCC
FCD6
FC57
FBBA
FBB2
FC6A
FD1E
FCCF
FB7E
FA83
FB42
FD5B
FEAA
FDB9
FC06
FD00
0236
0911
0D1A
0C7E
09AF
0868
09C2
0BB7
0C21
0B2D
0A91
0B1C
0BC6
0B10
08A9
05B0
039A
0317
03C4
04A7
0500
04C0
044C
03ED
0396
0335
0312
0388
0468
04F4
049F
03AE
02DD
02A4
02F2
0381
0417
047A
0487
0461
0462
049A
0492
03D7
02C9
0272
034C
0489
04EB
0458
0421
058D
084B
0AAF
0B67
0ACA
0A41
0A94
0B30
0B29
0A8A
0A30
0A7E
0ACE
0A76
09EC
0A2D
0B1F
0B57
0A08
088F
08F0
0AC3
0ADF
06D7
0044
FB73
FAD2
FC95
FD45
FBCA
FA13
FA1D
FB91
FCB7
FCB6
FC07
FB19
F998
F74B
F4E9
F391
F3A4
F47D
F543
F59C
F5A1
F57B
F548
F528
F52E
F54E
F57F
F5CE
F61B
F610
F582
F4D5
F4A1
F505
F584
F598
F542
F4E1
F4AC
F483
F43E
F3F3
F3DB
F41A
F4AA
F552
F5A3
F56F
F547
F639
F89F
FB64
FCDF
FC7D
FB48
FABA
FB42
FC1E
FC69
FBF7
FB41
FADF
FB2E
FC13
FCED
FD16
FCB2
FC91
FCFF
FD31
FC77
FBDA
FD93
027A
086F
0C22
0C5E
0AFD
0A6E
0B10
0B74
0AA8
0969
0906
09C8
0AB5
0A93
08EF
0662
041B
0317
0377
0462
04C4
0449
038D
0352
03B8
044B
0494
0463
03D0
033E
0325
039E
0426
0419
036D
02C1
02A2
0302
0377
03D3
0424
044C
0406
037C
0353
03D2
0465
044D
0397
031A
0389
04ED
06E4
08F0
0A82
0B1B
0ACF
0A70
0ABE
0B72
0B95
0ACF
09D9
0972
098B
09B6
09F0
0A4C
0A5B
09B0
08EE
094C
0AA2
0AB3
075D
0167
FC1A
F9E1
FA20
FACB
FB0F
FB7C
FC41
FC98
FC2A
FBCD
FC33
FC7C
FB13
F7F4
F51E
F466
F567
F638
F5BA
F494
F40B
F488
F565
F5C7
F571
F4E6
F4D2
F54B
F5B8
F589
F4E9
F491
F4E0
F56C
F5A4
F59E
F5C2
F5EB
F57F
F496
F435
F4F1
F5ED
F5EE
F508
F475
F4D5
F56E
F57D
F59B
F70E
F9DE
FC84
FDA6
FD65
FCBB
FC38
FBF0
FBFE
FC5D
FC97
FC58
FC17
FC85
FD54
FD62
FC73
FBE1
FCBF
FDF0
FD7D
FBE3
FC62
0108
0791
0B9B
0B94
09FE
09D4
0B12
0BAA
0AD8
0A14
0AB1
0BF1
0C24
0AC5
08B2
06C1
0515
03B6
02E7
02C0
02F1
032E
036C
03AA
03B4
0371
0329
0329
033B
02EB
0255
022B
02AC
033B
0344
0325
0384
0432
045E
03E1
0388
03F6
04A2
048E
03B3
031C
0378
0428
041D
0350
02EF
0418
06B8
0993
0B36
0B18
0A07
0964
09CD
0AAA
0B1C
0B14
0B1E
0B57
0B30
0A74
09EC
0A49
0ADF
0A64
090D
08A6
09F0
0ACC
0859
029E
FCF7
FA6F
FAB1
FB2B
FA98
FA1E
FB00
FC7D
FCD6
FBC8
FADF
FB64
FCC1
FD3C
FBCB
F901
F65E
F508
F504
F577
F586
F50B
F486
F46E
F4AE
F4E2
F4FA
F54A
F5F1
F685
F692
F62C
F5BD
F58C
F5A3
F5E4
F60A
F5C1
F511
F493
F4D1
F585
F5CD
F54C
F4B6
F4E1
F596
F5E8
F5A4
F589
F5E9
F607
F56C
F526
F6B3
F9DD
FCA3
FD72
FCD3
FC67
FCD9
FD7D
FDA6
FD6A
FCF9
FC3B
FB83
FBA2
FCB0
FD6E
FCD7
FBC5
FBE3
FD2B
FDB6
FCA4
FC0F
FED6
04C0
0A4C
0C8F
0C0B
0B1B
0ACF
0AA1
0A68
0AD5
0BEA
0C5F
0B5C
09ED
09B5
0A81
0A54
080C
04FB
033D
0341
03C9
03D3
037D
0341
0327
0316
032F
037E
03AB
036A
0307
031F
03B3
041E
03FC
03B4
03C4
03F6
03C7
0347
02FE
031A
0342
0341
035E
03E0
047D
04B4
047E
0459
047A
0463
039A
028E
0270
0407
06DF
09A0
0B20
0B3E
0AC2
0A75
0A61
0A22
09C5
09E0
0AA5
0B4E
0AF7
09DF
093A
09A2
0A45
0A24
09B0
0A33
0B7B
0B31
0760
0122
FBE4
FA08
FAD7
FBE9
FBDD
FB34
FAF3
FB35
FB5C
FB32
FB33
FBD4
FCBC
FCDB
FB4B
F853
F57A
F44C
F4D6
F5AC
F596
F4D1
F46D
F4C5
F536
F53E
F535
F5A1
F62F
F619
F554
F4BF
F4EF
F584
F5EB
F626
F65E
F63E
F577
F48B
F461
F510
F5AE
F590
F522
F51A
F556
F52F
F4BE
F4C8
F55A
F58A
F519
F549
F742
FA2F
FC1B
FC5C
FC30
FCBD
FD8B
FD8D
FCEF
FCC0
FD2E
FD40
FC95
FC05
FC29
FC51
FBE6
FBB8
FCA8
FDB2
FD03
FB2C
FB87
0045
0714
0B56
0B60
09DF
09C5
0AC1
0AD8
09FE
09F9
0B48
0C2D
0B61
0A12
0A15
0AF4
0A68
0795
0464
030F
037F
0405
03CA
035E
033A
0310
02B7
02BE
0387
0474
0490
03DB
0336
031F
0321
02B8
0233
022C
02A5
031C
035D
038E
03AE
0383
0327
0316
0380
03FB
041B
041C
0481
0508
04B2
032C
01CB
0285
05C6
09C3
0C21
0C1E
0AF9
0A6B
0AE4
0B71
0B26
0A47
09C0
09D9
09FD
09C9
09BC
0A6C
0B58
0B59
0A4B
0999
0A5E
0B65
0A04
053E
FF52
FB85
FADB
FB9F
FBE5
FB92
FBAE
FC76
FCEC
FC46
FB24
FAE4
FBF7
FD37
FCFC
FAAA
F754
F4CF
F421
F4AB
F506
F4A3
F438
F494
F57A
F5FD
F5BF
F54C
F53D
F579
F58E
F571
F580
F5CB
F5FD
F5E5
F5B7
F581
F509
F46B
F450
F511
F5FE
F61C
F579
F519
F587
F61B
F5FD
F564
F51F
F545
F546
F54F
F67E
F928
FBD7
FCD7
FC50
FBDD
FC5E
FD1D
FD43
FD1C
FD50
FDA2
FD63
FCDE
FD07
FDC6
FDC1
FC80
FB6B
FBC4
FC9D
FC5A
FBC7
FDD6
03A6
0A2E
0D3C
0C2E
0A33
0A00
0AF4
0B1B
0A59
0A12
0A9C
0ADA
0A67
0A63
0B6B
0BFB
0A11
0618
02E1
0277
03F7
0513
04C8
03D9
0333
02FC
0311
0369
03C9
03C2
034E
030D
0374
040C
0403
0357
02EC
0349
03DD
03D9
034E
02EF
0303
0333
0347
036C
03C3
040C
0413
0412
0455
0492
041C
02EC
0226
031E
05E1
08F9
0AC1
0ACD
0A0F
09B1
09EF
0A1D
09B3
090F
08F3
096C
09C8
09A6
098B
0A0C
0ABF
0AC0
0A1E
0A07
0AF5
0B44
0894
02CA
FCD2
F9D6
FA28
FB80
FBE5
FB83
FB96
FC64
FCE9
FC56
FB38
FAD0
FB7A
FC1E
FB56
F8EE
F62A
F48A
F468
F4D3
F4D3
F484
F4B2
F586
F630
F60A
F57C
F558
F5AD
F5CC
F551
F4AB
F474
F4B2
F505
F553
F5CB
F65C
F6AB
F6A6
F69D
F6A3
F664
F5D7
F592
F5E5
F637
F5DD
F54F
F5AE
F706
F7E8
F753
F667
F734
FA00
FCC2
FDA9
FD24
FCD4
FD46
FDAD
FD6A
FCD5
FC79
FC66
FC8D
FD17
FDDC
FE0E
FD32
FC29
FC35
FD07
FCF4
FBB0
FB99
FF17
0539
0A4A
0BE2
0B28
0AB7
0B4A
0B9A
0AE1
0A09
0A08
0A6A
0A5B
0A39
0AE6
0BD5
0B2A
0825
0478
0288
02CA
039A
037F
02BE
0273
02EE
0381
039D
0360
031F
02F6
02FC
0358
03E9
0426
03A4
02B6
022D
027A
0336
03AA
038A
0314
02A8
027F
02A9
0310
0386
03FA
0489
0523
053A
0430
0251
0113
01EA
04BF
07E7
09BD
0A2C
0A58
0B18
0C0B
0C42
0B64
0A10
092E
0917
0972
09C1
09EC
0A28
0A7D
0AA3
0A75
0A5D
0AD1
0B4E
0A35
0649
0084
FBC1
FA38
FB65
FCDA
FCE4
FC00
FB95
FBEF
FC16
FB68
FAB4
FB2F
FCB9
FD9D
FC4E
F907
F5A2
F3DC
F3F1
F4C3
F52F
F502
F4B1
F483
F456
F41F
F430
F4C4
F587
F5E0
F5A0
F526
F4DE
F4D4
F4E3
F510
F56B
F5B8
F5A4
F54B
F52A
F567
F597
F56E
F53B
F563
F5CE
F621
F658
F693
F68F
F5DD
F4EA
F51B
F749
FA6B
FC87
FCF0
FCB5
FCD3
FCFE
FCC0
FCA6
FD64
FE61
FE4A
FD09
FC0D
FC50
FD04
FCF5
FC70
FC8F
FD1C
FCD0
FC02
FD3E
0205
081C
0BB8
0BD9
0AEE
0B38
0C2C
0C17
0B08
0A8D
0B16
0B5D
0AB3
0A49
0B21
0BF5
0AA0
0725
03F0
02FB
03CC
049C
047D
03D9
035E
033B
0361
03C3
0417
03F7
037F
0353
03AB
03E0
0372
02EA
030B
0396
039C
02FE
02B9
0372
046C
0475
0386
02C6
02ED
0365
0359
02F5
02F8
0366
0379
02DC
0260
0328
056D
083E
0A5C
0B2F
0B06
0A8E
0A37
0A0D
09FB
0A00
0A1D
0A2B
09FD
09BC
09E4
0A9E
0B3E
0AEE
09EE
0990
0A74
0B2A
095B
0469
FE88
FACB
FA52
FBA1
FC94
FC72
FBF7
FBCF
FBBE
FB48
FAB0
FAD4
FC00
FD34
FCD9
FA59
F6E0
F463
F3DC
F4A4
F574
F5BF
F5DC
F622
F64A
F5E2
F509
F46D
F48A
F528
F5B7
F5E1
F5BB
F584
F569
F57D
F5B4
F5E6
F5F3
F5ED
F5F7
F600
F5C6
F53D
F4CA
F4E0
F56F
F5F8
F630
F648
F672
F676
F626
F609
F718
F97C
FC06
FD46
FD19
FCA1
FCC2
FD2F
FD34
FCDB
FCCC
FD3B
FD93
FD48
FC92
FC12
FC14
FC7D
FD1A
FD90
FD38
FBF8
FB4C
FD74
02E6
0917
0CAC
0CBF
0B58
0ABF
0B3B
0BB4
0BB1
0BAB
0BC5
0B80
0AE0
0AC4
0B63
0B57
0937
05C2
034D
0315
03F5
0423
036A
02F9
0380
0456
049C
0451
03EB
0384
0319
0305
0394
0450
046D
03D6
033D
0318
0314
02C9
0272
0291
0307
0321
0299
0211
0237
02E5
037A
03BF
03E7
03EB
037B
02BC
029B
0401
06BF
0976
0AC3
0A7C
09C3
09C4
0A7F
0AFF
0A91
099A
0909
0939
09AD
09DF
09F2
0A2A
0A2E
098B
08D4
0940
0AA9
0AC6
075D
012C
FBAA
F9AD
FABF
FC32
FC4D
FBA6
FB86
FBF1
FBDF
FAEC
FA01
FA38
FB83
FCA1
FC41
FA2E
F77D
F590
F4D7
F4AF
F462
F411
F452
F52D
F5E4
F5DD
F565
F534
F55D
F547
F4C0
F46E
F4EB
F5D9
F65C
F63E
F60C
F625
F639
F5EC
F584
F595
F62A
F6A9
F6A7
F66A
F666
F68C
F672
F608
F5C0
F5F0
F652
F664
F625
F63A
F749
F93C
FB38
FC54
FC68
FC1E
FC4C
FD2A
FE2D
FE93
FE15
FD17
FC44
FC0B
FC77
FD42
FDF3
FE0A
FD67
FC9D
FC92
FD6C
FE1B
FD74
FBF5
FBE2
FF1B
04D5
0A01
0C3D
0BF5
0B50
0B7E
0BCF
0B58
0A75
0A1B
0A64
0AAB
0AC6
0B39
0BEC
0B99
093B
05BB
0350
030F
03D8
03F0
031F
028E
0305
03FD
047B
0429
0375
02F5
02F1
035B
03E2
0422
03F2
0394
036D
0391
03AB
037E
0333
0309
02FF
02F9
0318
0385
0411
0447
03EC
0349
02E6
0311
0388
03A4
0301
021A
0209
0382
060D
0869
09B4
0A1A
0A3C
0A52
0A30
09F5
0A06
0A59
0A71
0A3C
0A5C
0B0D
0B7C
0AD5
09A3
0942
09F4
0A6E
09BD
08E4
0983
0B24
0B06
0736
0110
FBFF
FA21
FAD4
FC14
FC7A
FBF2
FB3A
FAFC
FB3E
FB7A
FB61
FB5C
FBF8
FCC1
FC3F
F9A8
F64E
F482
F4FB
F615
F60A
F510
F48D
F4F2
F55B
F52A
F4E1
F523
F59C
F583
F4E1
F498
F520
F5D8
F5EB
F569
F4FF
F4F3
F4FE
F4ED
F4FB
F561
F5FD
F67B
F6A9
F696
F674
F662
F64F
F619
F5C7
F592
F5A0
F5CF
F5F0
F637
F73F
F94E
FBBE
FD5D
FD9C
FD1A
FCD9
FD1B
FD5E
FD39
FCE1
FCC1
FCE2
FCF7
FCD9
FCCC
FD12
FD70
FD5C
FCDC
FCC0
FD8F
FE7A
FE26
FCC2
FC9C
FFD6
05A7
0AA8
0C4D
0B64
0AA3
0B40
0C18
0C0A
0B98
0BA3
0BC2
0B1A
0A19
0A0A
0AE8
0AE8
08C0
0586
0374
0341
03A2
0369
02EF
0307
038D
03D9
03DE
03FD
041E
03DA
0356
0322
0353
0361
0316
02F8
0375
0415
0417
0396
0366
03C9
040C
03BD
0361
037C
03A5
0345
02B2
02AE
0326
0356
02FF
02B1
02CB
02E7
02C0
0316
04EF
0803
0AA6
0B9F
0B5F
0B17
0B30
0B43
0B03
0A90
0A26
0A09
0A78
0B2B
0B47
0A57
0920
08E1
09AA
0A2E
098D
08BD
0938
0A7B
09FE
0634
00AA
FC79
FB19
FB84
FBF7
FBB9
FB2B
FAEF
FB43
FBDE
FC2E
FBF0
FB87
FB91
FBFD
FBCB
FA1F
F771
F53C
F463
F468
F474
F472
F4BC
F53E
F58F
F5A9
F5D9
F61F
F618
F5A8
F541
F54B
F59B
F5B3
F57A
F54F
F56F
F59C
F585
F54F
F55F
F5D0
F661
F6BA
F6A1
F61C
F57F
F534
F542
F550
F537
F54A
F5BF
F62A
F606
F5B3
F657
F88E
FB73
FD69
FDBB
FD24
FCB5
FCB8
FCDC
FCEE
FCF9
FCE1
FC72
FBD0
FB77
FBB7
FC5F
FCE4
FCE2
FC93
FCA0
FD39
FD9B
FCFF
FC28
FD53
01DD
0825
0C90
0D13
0B3D
0A20
0AC7
0BBF
0BD3
0BA0
0BF7
0C37
0B71
0A57
0A6C
0B83
0B7B
08EF
053E
0305
0324
0426
047B
041A
03B8
0370
0308
02BD
02E2
032A
0322
02F8
031C
0368
035E
0312
0325
03C5
0451
0435
03BC
038C
03A5
038E
0353
037E
03F1
03D1
0303
02A0
034B
0403
0399
0293
026E
035A
03F3
0379
0330
04D1
0822
0B08
0BED
0B32
0A24
097D
0967
09F1
0ACA
0B31
0AF3
0AD8
0B64
0BD7
0B53
0A5D
0A3B
0AE9
0AF4
09C1
08D7
09CC
0B65
0A61
0577
FF33
FB20
FA24
FA94
FAE3
FAE8
FAED
FAF0
FAF5
FB3A
FBB8
FBFD
FBD9
FBAC
FBA8
FB19
F936
F68E
F4CF
F4D4
F5A2
F5DC
F566
F501
F4F6
F500
F512
F558
F59C
F56D
F4ED
F4CE
F549
F5A0
F520
F44C
F44E
F558
F63A
F5F4
F4F3
F453
F473
F4E9
F55A
F5C0
F603
F5FF
F5E0
F601
F668
F6BF
F6E3
F708
F72F
F6EE
F635
F5FD
F76D
FA35
FC78
FCD9
FC0C
FBC7
FC91
FD6A
FD6E
FCEF
FCB2
FCBE
FC9A
FC4A
FC65
FD0D
FD75
FD02
FC65
FCD9
FE41
FEE9
FDCB
FC71
FDB2
025A
07EC
0B31
0B8A
0B10
0B96
0C96
0C89
0B6B
0ABC
0B37
0BCE
0B6E
0AB2
0AE5
0BD6
0BCC
09BB
06A2
0469
03D0
0408
03FB
0372
02E1
02AE
02F9
039F
042D
0426
039C
032C
0320
0316
02CC
02AE
0327
03D4
03FD
03AC
038E
03DB
03ED
0363
02F3
037C
048C
04CE
0405
0362
03A2
03E9
0352
0289
02C2
03B1
03E2
0305
02B8
047F
07B0
0A34
0AEE
0A97
0A50
0A63
0A9F
0B01
0B55
0B12
0A45
09E3
0A79
0B34
0B10
0A78
0A9A
0B6B
0B85
0A5E
096D
0A0F
0AE9
0901
03A3
FDB2
FA6B
F9F8
FA49
FA36
FA55
FB19
FBC7
FBA2
FB13
FAF7
FB5F
FBBC
FBF1
FC54
FC8C
FB74
F8A9
F58C
F3F6
F439
F51E
F588
F565
F524
F4F9
F4DA
F4C8
F4C5
F4C0
F4B2
F4BF
F502
F549
F53F
F4ED
F4C7
F510
F577
F595
F575
F572
F59B
F5A8
F56E
F51F
F51C
F594
F651
F6D3
F6BF
F64F
F62D
F6A6
F726
F6D2
F5C9
F575
F725
FA61
FD28
FDF7
FD38
FC75
FC80
FCED
FD16
FCFA
FCE5
FCD4
FC9B
FC74
FCC7
FD71
FDB2
FD30
FCAF
FD28
FE44
FE86
FD66
FCB3
FEF8
0469
0A20
0CF1
0C94
0B7A
0BA8
0CA4
0CCB
0BCF
0AF8
0B09
0B25
0A4B
0915
0904
0A4A
0B26
09D6
0696
035C
01DA
0225
0328
03DC
03E9
0381
0317
0312
0379
03F0
041B
03F7
03AB
0340
02BF
0269
027F
02E2
0323
0313
02FA
032D
0390
03BD
0392
0357
0346
0342
032B
032A
036C
03C2
03DC
03BD
03A4
0396
0355
02EB
0300
0460
0711
09FB
0BB4
0BB1
0AB5
0A05
0A39
0AD7
0B07
0A94
0A09
09DF
09E5
09B7
0997
0A1B
0B09
0B3E
0A38
0924
098E
0B19
0B45
0811
026C
FD6A
FB34
FB44
FBB0
FB73
FAF4
FAD3
FB12
FB5D
FB8E
FBA2
FB94
FB80
FBB0
FC35
FC76
FB88
F92B
F654
F476
F43D
F518
F5EB
F60B
F59A
F526
F504
F513
F50B
F4EE
F4FB
F547
F578
F52D
F48A
F42F
F491
F570
F611
F5F6
F54B
F4AA
F487
F4E2
F567
F5B5
F5A9
F577
F56A
F59A
F5DD
F610
F653
F6BA
F6F5
F68E
F5B5
F577
F6CD
F96A
FBCA
FCA8
FC46
FBF4
FC87
FD8B
FE16
FDE8
FD7F
FD46
FD30
FD28
FD54
FDB0
FDCD
FD5A
FCCF
FCE9
FD83
FD91
FCBC
FC9A
FF4A
04CB
0A54
0CF3
0C6F
0B0C
0ABD
0B54
0B8D
0B1B
0ADF
0B5A
0BD7
0B75
0A81
0A18
0A9C
0B0D
0A24
07CA
0532
03A9
036E
03BD
03C1
0360
0318
034C
03C8
0408
03CA
0353
0324
0372
03FB
0450
0439
03E2
03AC
03D2
0428
0435
03B6
0310
02F7
039E
0460
0480
0412
03E4
0479
0554
058D
04DA
03D3
0327
02F4
02F1
02E6
02D1
02C4
02FB
03E5
05C9
082F
0A0B
0A99
0A1E
097F
0957
098D
09CB
09ED
09F5
09DF
09C7
09F8
0A7F
0ADC
0A98
0A15
0A37
0AD5
0A1F
065C
005B
FB49
F9AD
FAE4
FC3E
FC21
FB5E
FB5F
FC09
FC23
FB4F
FA9C
FAEF
FBCF
FC30
FBE8
FB98
FB83
FB4C
FAE7
FAF6
FBB9
FC27
FADB
F7E7
F521
F43D
F516
F622
F641
F59D
F4FD
F4C9
F4D9
F4DB
F4AC
F46F
F468
F4BC
F531
F556
F509
F4BA
F4EA
F572
F5A5
F545
F4F8
F574
F67A
F70B
F697
F596
F4EF
F501
F581
F5F4
F629
F628
F603
F5DD
F5E4
F625
F65D
F63A
F5CB
F59F
F670
F888
FB5D
FDC1
FEB6
FE49
FD81
FD53
FDBB
FDFF
FDBD
FD59
FD54
FD8C
FD85
FD4C
FD6F
FE04
FE3A
FD82
FCE0
FE54
0298
07E4
0B67
0BF8
0AEF
0A59
0AC7
0B40
0AF4
0A56
0A58
0B1C
0BD2
0BDB
0B85
0B7A
0BD1
0BFC
0B96
0AF0
0AB5
0B17
0B6F
0ABF
08A6
05E5
03E6
038A
0462
051C
04DB
0402
038C
03CE
0434
0433
03EF
03CC
03BC
036A
02E7
02A0
02CA
0323
036F
03D8
0486
0519
04FE
0440
038A
0343
0332
031C
0342
03D3
045B
044C
03C8
0370
0379
0380
0351
033F
0373
0362
02AD
0239
0375
065C
0919
0A1F
09DB
09BB
0A2E
0A84
0A61
0A48
0A94
0AC6
0A67
09E1
09D0
09E1
0965
08D9
0982
0B08
0AC4
06B0
005F
FBB0
FAA2
FB9B
FBFB
FB4D
FB04
FBDE
FCCC
FCAA
FBD4
FB5E
FB63
FB23
FA71
FA11
FA87
FB52
FBAD
FBA5
FBDA
FC59
FC23
FA37
F6F8
F42D
F36C
F495
F605
F63A
F532
F41D
F3EE
F46A
F4BB
F499
F482
F4D8
F551
F57A
F56C
F596
F609
F65B
F63B
F5D5
F586
F570
F576
F581
F59B
F5C4
F5F0
F61C
F656
F68A
F688
F657
F641
F679
F6CC
F6EC
F6D9
F6BD
F689
F607
F56A
F57B
F6EE
F979
FBD9
FCE5
FCA3
FC21
FC40
FCD8
FD29
FCF4
FCC8
FD32
FDE9
FE19
FD88
FCE4
FCBE
FCA5
FC00
FBA8
FDA0
02A9
08B6
0C92
0CF6
0B78
0A76
0ABA
0B6E
0BBA
0BB0
0BA9
0B9E
0B6F
0B56
0B8D
0BDD
0BDB
0B6C
0AC7
0A41
0A48
0B1E
0C2F
0C00
0997
05F2
0377
0375
04B5
050D
0416
034E
03AF
044E
03F7
0313
02E8
0390
03DD
0340
02A1
02F7
03D1
040C
0396
0383
0455
0529
04FF
0415
0356
0306
02BF
026E
0282
030D
037C
0368
0322
0329
0356
032B
02BB
02AD
032E
0384
0324
02BD
039D
0613
08F5
0AC7
0B0D
0A65
09B6
0987
09DF
0A79
0B07
0B60
0B8D
0B93
0B43
0A84
09D2
0A13
0B7C
0C9B
0B3B
068E
006B
FBE6
FA97
FB67
FC1D
FBBF
FB1A
FB34
FBD7
FC14
FBAE
FB4A
FB58
FB73
FB2D
FADC
FB0D
FB87
FB92
FB2D
FB4B
FC64
FD4C
FC4B
F944
F61F
F4CB
F557
F657
F6A4
F627
F559
F4A8
F45F
F48F
F4E3
F4DB
F473
F447
F4C3
F568
F55B
F49E
F42A
F496
F544
F54C
F4BE
F475
F4D8
F573
F5BB
F5B0
F5A9
F5BE
F5C7
F5BD
F5D0
F612
F64A
F63D
F5F0
F594
F55B
F572
F5D9
F644
F690
F749
F91E
FB9C
FD18
FC99
FB46
FB3A
FCE5
FE83
FE7F
FD85
FD5C
FE42
FEBD
FE12
FD60
FDA0
FDE4
FCFB
FC15
FE07
0397
09CD
0CEB
0C57
0AB0
0A5B
0B3D
0BFD
0C29
0C34
0C34
0BC8
0B07
0A91
0AA3
0ADE
0B00
0B39
0B8F
0B8C
0B06
0AA9
0B04
0B3E
09C1
067B
0379
0294
0346
039F
02F2
026D
030C
0418
043B
036B
02DB
0332
03C1
03C0
0375
0398
041C
0451
03FC
039B
0394
03BB
03D4
03FD
0450
0475
0410
037A
0369
03D9
03EF
0331
0261
0287
0381
0431
040B
03B7
03DA
03F9
0345
0243
02AA
054D
08C5
0ADA
0ADA
0A08
09C4
0A1A
0A4B
0A20
0A19
0A72
0ABD
0A82
09DD
093D
0908
098A
0AC0
0BB6
0A9E
0673
009F
FC33
FB02
FBEB
FC79
FBCA
FB10
FB53
FBED
FBC7
FB21
FB22
FBFF
FCA2
FC4A
FB9C
FB98
FC19
FC2A
FB8C
FB22
FB88
FC06
FB62
F95A
F6D0
F4DE
F423
F4A2
F5C1
F67B
F633
F55B
F4EE
F53B
F59C
F57E
F548
F5B6
F685
F6AA
F5D7
F502
F500
F562
F54D
F4D9
F4C9
F541
F594
F55D
F514
F537
F57B
F566
F540
F5B8
F6A6
F70B
F67B
F5BB
F589
F598
F55A
F50F
F53C
F5A5
F5C9
F62E
F801
FB20
FD8B
FDA4
FC6A
FC3D
FD9E
FEA5
FDF3
FCAD
FC93
FD5F
FD84
FCE6
FCFF
FE34
FEC0
FD63
FC04
FDF7
03B5
09CF
0CB6
0C5D
0B43
0AF3
0AF3
0A9D
0A6D
0AF7
0BC7
0BFC
0B8C
0B2A
0B1D
0B00
0AAA
0A99
0B12
0B89
0B80
0B68
0BD7
0C33
0B0D
080F
04C0
02F6
02EE
036A
0373
0344
036B
03BA
03A4
0338
0311
0366
03AD
036D
02E9
02B0
02D6
02F6
02DF
02D6
0313
0365
0389
039B
03DC
0433
0441
03F2
039B
0375
0344
02D7
0291
02F8
03D6
0444
03CE
030B
02C9
02FA
02F3
02B3
032F
052C
081D
0A84
0B69
0B10
0A58
09DB
09C4
09F7
0A2F
0A27
09F8
0A01
0A43
0A3C
09CE
09CA
0AE4
0C0A
0ABB
05C2
FF34
FACE
FA2F
FB89
FC30
FB97
FB17
FB91
FC5E
FC88
FC0C
FB92
FB72
FB8B
FBC2
FC18
FC54
FC1C
FB9B
FB88
FC37
FD08
FD12
FBFE
FA05
F797
F578
F4A6
F56F
F6B9
F6EE
F5C1
F48F
F497
F565
F593
F4DE
F475
F524
F621
F637
F570
F4C4
F4A1
F49E
F484
F4B4
F559
F5E6
F5C8
F549
F52A
F595
F5FD
F622
F663
F6E4
F71B
F6AD
F626
F635
F698
F694
F621
F5E8
F619
F619
F5AF
F5D0
F77D
FA21
FBFE
FC52
FC34
FCDC
FDF2
FE4F
FDD2
FD71
FDA6
FDD6
FD86
FD3C
FD9A
FE20
FDBB
FCB5
FD0C
0052
059B
0A2B
0C19
0BC5
0ADA
0A89
0AE7
0B79
0BD7
0BE1
0BAC
0B78
0B7D
0BA5
0B90
0B08
0A6F
0A65
0B05
0BAC
0BBE
0B65
0B3B
0B46
0AA4
0887
0572
0303
025F
030A
03A6
039A
0379
03DA
0463
045C
03C3
0341
032B
031E
02C5
027E
02D8
039F
0400
039C
02FF
02D2
0307
0327
031B
033A
03A2
0409
043B
0462
049E
04A4
0419
0330
0295
02AA
030F
0332
0306
02EF
0323
037B
03F1
04EC
06CF
094D
0B54
0BE0
0AF8
09BF
095A
09D6
0A4B
0A10
097F
0957
09AD
09DF
09B6
09E4
0AE6
0B9E
09FA
0552
FFA8
FBEF
FB3C
FC18
FC72
FBB0
FABF
FA94
FB2F
FBEA
FC41
FC15
FB86
FAE7
FAB2
FB1F
FBCC
FBFD
FB62
FA82
FA4F
FB35
FC7F
FCBF
FB07
F7F3
F53C
F42B
F47E
F4EE
F4B6
F44F
F48B
F55B
F5D3
F55C
F46A
F3E0
F419
F4C6
F578
F5E8
F5F8
F5BE
F590
F5B6
F5F9
F5C9
F4FC
F439
F45A
F577
F6C4
F769
F734
F67F
F5B7
F53C
F551
F5D9
F648
F62C
F5BC
F58A
F5CC
F624
F634
F618
F626
F664
F699
F6DF
F7BC
F983
FBC6
FDAA
FE94
FE76
FDB9
FD04
FCD6
FD20
FD66
FD6B
FD84
FDF5
FE52
FDF5
FD0B
FC87
FCD4
FD1E
FCAF
FC9E
FF12
0461
09FA
0CD6
0C90
0B49
0AE5
0B47
0B5C
0AD1
0A4B
0A4C
0AB6
0B4A
0BEF
0C5E
0C39
0BB0
0B81
0BE9
0C25
0B9B
0AF3
0B2E
0BF7
0BBA
0999
06A6
04A6
041C
0423
03F5
03BB
03B8
03A2
033E
0313
03A7
0487
04C1
0436
03B6
03BE
03D0
0353
029D
028B
033B
03DA
03C7
035B
0342
037C
038B
0349
030E
0319
0359
03B0
0413
0448
03FE
034C
02D4
0313
03AB
03BC
0308
024F
024E
02C0
02D6
028B
02E6
04B9
0771
0990
0A41
0A1A
0A36
0AC4
0AF1
0A37
094C
094F
0A46
0B0E
0AD0
0A07
09A8
09C5
09A9
0938
0958
0A64
0ACA
0848
02C5
FD0C
FA2A
FA77
FBBA
FBF1
FB24
FA95
FADE
FB75
FBA5
FB5F
FAFE
FAB6
FA8E
FAAF
FB43
FC07
FC62
FC00
FB49
FB0D
FBAC
FC7C
FC2D
FA19
F726
F50D
F48F
F4C8
F471
F37E
F311
F3DB
F528
F5BF
F55F
F4D0
F4B7
F4EB
F50B
F525
F558
F572
F55C
F582
F648
F735
F755
F67B
F5AB
F5EF
F71C
F80F
F808
F74A
F676
F5D7
F585
F5AC
F63F
F6C1
F6C9
F681
F650
F641
F629
F625
F675
F6E3
F6E1
F677
F6AB
F86B
FB3E
FD93
FE6B
FE2D
FDBC
FD71
FD52
FD97
FE4A
FEDF
FED0
FE6A
FE58
FE8A
FE43
FD52
FC86
FC77
FC87
FC19
FC5B
FF69
053E
0AC2
0CEF
0C16
0AF8
0B39
0BF3
0BC6
0AF6
0ABF
0B6C
0C1B
0C3A
0C31
0C59
0C4D
0BBD
0B1A
0AD0
0A7E
09CE
097B
0A6B
0BEA
0BE3
0951
05BB
0399
039E
0455
044C
03B4
038A
03FA
0459
044D
0424
042F
0459
0470
045D
0406
0367
02D2
02C4
0353
03E4
03CD
0329
02B7
02E6
0352
0360
0307
02B9
02C7
032B
03B1
040D
03F3
036C
02FE
0318
037F
0384
02F2
0267
0289
031E
0345
02B6
0260
0377
05FF
08A6
0A18
0A3C
0A02
0A2B
0A77
0A25
0935
08A4
093A
0A51
0A93
09CB
0936
09B0
0A66
0A1C
0941
0986
0B09
0B22
0731
004F
FAC0
F964
FAE2
FBF8
FB74
FAB9
FAED
FB62
FAFE
FA1A
F9F5
FAD9
FBC1
FBEA
FBD0
FC34
FCCD
FCAF
FBB2
FAC8
FAE5
FBE7
FC95
FB9F
F8CC
F574
F387
F3C1
F4FB
F588
F511
F4A9
F525
F5E9
F5CE
F4D7
F43C
F4C6
F5D9
F670
F65C
F60A
F595
F4E6
F45B
F49B
F595
F65F
F637
F570
F4FF
F550
F5EB
F62C
F604
F5D6
F5D4
F5DE
F5BE
F561
F4F3
F4D8
F544
F5DC
F60F
F5F3
F636
F6F8
F755
F6A3
F5D6
F6BD
F9CB
FD34
FEBE
FE1A
FCDA
FC56
FC8C
FCF4
FD74
FDFD
FE1B
FDA6
FD45
FD8D
FE10
FE0A
FDA8
FDAC
FDF1
FD6B
FC43
FCD0
0125
07E2
0D01
0E2A
0CF6
0C30
0C47
0BC7
0A55
097A
0A4D
0BE7
0CB7
0C87
0C3C
0C34
0BEF
0B48
0AD4
0AC5
0A81
09ED
0A10
0B5E
0C4E
0AE1
0764
045B
0383
03FC
03EA
030D
02B6
037F
0454
041B
035C
035B
0439
04D4
0461
0348
0275
0262
02EB
03A1
041B
0430
0407
03E7
03DF
03BD
0377
0358
0395
03D0
0381
02D4
0292
02F8
033C
02B4
01EF
0206
030F
03FF
040C
039D
037C
039F
0349
025D
01FE
0363
0651
0924
0A69
0A1F
096F
095A
09DC
0A50
0A6D
0A9C
0B2C
0B8E
0AFC
09C1
0917
097A
09E4
094E
086D
08CE
0A2B
09CC
0599
FF3D
FAF1
FAE8
FD1A
FE18
FD04
FBB6
FBA4
FC28
FC10
FB8C
FBB4
FC9D
FD16
FC64
FB71
FBA3
FCEF
FDD4
FD4A
FC06
FB7F
FC03
FC3A
FAAB
F79A
F502
F479
F564
F5B8
F47D
F2E9
F2BB
F40C
F54F
F54E
F46D
F3E2
F431
F4EC
F59B
F63C
F6C7
F6D9
F646
F584
F521
F523
F533
F52B
F51D
F50C
F504
F549
F5F7
F6A5
F6B4
F627
F5B8
F5EB
F650
F627
F575
F4F2
F4EE
F50E
F540
F5FF
F740
F7FF
F7A8
F75A
F8B9
FBB0
FE4D
FEFB
FE31
FD73
FD52
FD47
FD1C
FD5B
FE18
FE7A
FE07
FD84
FDC0
FE59
FE70
FE05
FDA7
FD35
FC3B
FB9C
FD84
02BC
08D5
0C40
0C23
0ADA
0A8D
0AC3
0A26
091B
0921
0A54
0B36
0AF5
0A7D
0AD7
0B87
0B71
0AA8
0A4C
0AAF
0AEC
0A9C
0AAF
0BB3
0C55
0AC4
0746
041D
02F4
034F
03D1
0408
0467
04EF
04E8
03FC
02DC
0262
0286
02AA
028B
025A
022F
01EF
01AF
01BD
0239
02F8
03C2
046F
04D4
04CE
0489
046F
049C
049C
0400
031B
02B7
02F7
0316
0290
01FD
0243
0332
03A9
0320
025F
0262
02F1
02FA
0232
01CF
0330
061A
08CC
09DF
0992
092D
096B
09F4
0A3D
0A55
0A9D
0AF5
0ACD
0A13
0995
09F0
0A84
0A2B
08FC
088B
09CA
0B3C
0A13
0559
FF52
FB60
FACF
FC1C
FD10
FCE5
FC36
FBB6
FB87
FB89
FB9A
FB91
FB5F
FB43
FB91
FC33
FC96
FC5A
FBD2
FBAF
FC22
FC89
FC0E
FA6C
F825
F61A
F506
F510
F59C
F5C7
F540
F494
F47C
F509
F5B5
F61A
F63E
F63F
F610
F5BA
F594
F5DF
F634
F5D3
F4A6
F3A3
F3D0
F506
F610
F5FE
F517
F471
F4C7
F5D6
F6CA
F724
F722
F731
F744
F6FB
F657
F5E7
F60C
F65C
F626
F589
F58A
F6BE
F84A
F8D4
F853
F839
F99F
FBF0
FDD0
FEB4
FEFA
FED3
FDFB
FCA2
FBD3
FC5C
FDAF
FE79
FE2F
FD7B
FD1D
FD1F
FD56
FDD6
FE6C
FE62
FD9D
FD94
0017
04F6
09AE
0BE2
0BAE
0B06
0B2D
0BA6
0B92
0B1C
0AF8
0B33
0B4D
0B21
0B02
0B12
0B24
0B34
0B71
0BA4
0B32
0A11
0950
09E7
0B21
0B00
088F
052B
0309
02D1
035F
0378
030C
02AA
0291
0293
02A0
02D8
0332
0369
036C
0376
039F
03A4
0356
0300
0304
0348
0365
034A
034B
0389
03B6
0392
0362
039A
0422
045F
03EC
0308
0221
015B
00C8
00C3
018B
02A6
0328
02C0
0220
0206
0244
0234
0203
02D9
0558
0877
0A75
0ABF
0A59
0A5B
0AB8
0ADC
0AE9
0B83
0C71
0C77
0B00
0956
093A
0A7D
0AFE
096B
0747
072C
0936
0A41
0745
00FD
FB54
F956
FA5D
FB79
FAF7
F9DA
F9F0
FB5A
FC7E
FC1F
FAD2
FA25
FAB7
FBA8
FBDA
FB50
FB05
FB8D
FC59
FC8B
FC1D
FBC2
FBA2
FAE1
F8C4
F5FF
F448
F47B
F59A
F5F4
F513
F40A
F3FA
F4CA
F59D
F5FC
F623
F64C
F654
F624
F611
F663
F6C5
F685
F587
F483
F44A
F4EE
F5E3
F6A8
F70F
F70F
F6B4
F64B
F646
F6C2
F759
F7A3
F7BC
F808
F880
F8AA
F847
F7B0
F741
F6E4
F680
F6AA
F837
FAED
FD43
FDE2
FD2B
FCAA
FD16
FD99
FD2A
FC08
FB31
FAF6
FACD
FA88
FACB
FBE9
FCFE
FD11
FCE9
FEA6
0318
0847
0B4C
0B62
0A65
0A65
0B87
0C90
0CC2
0C8D
0C92
0CBD
0C99
0BFF
0B24
0A49
09BD
09CE
0A5C
0AB9
0A66
09E1
0A1F
0B12
0B40
095B
060A
0371
02F0
03D9
048D
0459
03C3
0378
03A2
0428
04EB
0593
058F
04BA
03B2
0338
0354
0379
0373
03A1
0412
041E
035A
0270
0271
0353
03EB
037C
02B0
0295
0314
031B
023D
015B
0170
024D
0310
0375
03F0
049D
04DE
044F
03A5
040D
05CE
07FB
0983
0A1F
0A22
09CE
0939
0895
082E
0829
0880
0918
09AE
09C8
0937
08AD
0936
0AAC
0B0E
0846
02AF
FD44
FAC2
FB20
FC22
FC1A
FB4B
FACA
FAE8
FB29
FB42
FB55
FB55
FAF7
FA69
FA5E
FB08
FB8B
FB11
FA13
F9E3
FAF7
FC52
FCB5
FBE4
FA63
F879
F63F
F45D
F3CF
F492
F55E
F529
F477
F480
F560
F606
F5C6
F537
F52A
F56F
F552
F4F4
F53E
F66F
F784
F787
F6DA
F687
F6C0
F6BE
F600
F4FF
F487
F4D7
F59C
F676
F721
F762
F729
F6CF
F6C6
F6FA
F6FA
F6B3
F68D
F693
F645
F5B0
F5FD
F827
FB4D
FD48
FD1B
FC14
FC14
FD3A
FE12
FDC3
FD03
FCB7
FCBE
FCA2
FCA4
FD1B
FD6A
FCCC
FC1B
FD97
0234
07E2
0B6E
0BE0
0B0E
0AF5
0B96
0BE9
0BD0
0BFE
0C81
0C93
0BF5
0B70
0B92
0BAF
0AE9
09B8
0977
0A6A
0B35
0AC7
09ED
0A18
0AFD
0A94
07B9
03E7
01BB
020E
034C
0397
02D6
0264
031B
0468
0526
04ED
0440
03DF
041B
04BF
054D
0559
04D2
040F
038A
037C
03BD
03F7
03EE
0394
02FF
0273
0243
0282
02C5
0281
01A7
00D8
00BC
0159
0224
02C0
034A
03DA
040A
037B
02AD
02F1
0525
0896
0B70
0C6B
0BD8
0B0E
0AE6
0B0F
0AD5
0A2F
09C8
0A0F
0A80
0A3F
095D
090B
0A1C
0B76
0A9B
063A
FFF6
FB26
F9B8
FAA4
FB84
FB3D
FA9B
FAA2
FB27
FB66
FB40
FB3D
FB8C
FBB3
FB6A
FB2F
FBA1
FC87
FCED
FC50
FB4C
FAEF
FB93
FC86
FCA0
FB32
F8A2
F645
F54D
F5A5
F605
F572
F45E
F401
F4AB
F560
F540
F4C4
F4F4
F5C8
F61F
F578
F4C8
F51D
F611
F656
F587
F499
F47E
F501
F55F
F56F
F5AE
F650
F6EF
F733
F739
F729
F6E3
F673
F642
F678
F68E
F612
F57D
F596
F62B
F635
F573
F532
F6C6
F996
FBA5
FBFD
FBB5
FC25
FD1C
FD85
FD28
FCCA
FCD2
FCD6
FCA5
FCC3
FD58
FD73
FC5D
FB68
FD1A
0220
07EC
0B3F
0B80
0ACB
0B02
0BEA
0C47
0BCF
0B45
0B30
0B40
0B18
0AEF
0B10
0B41
0B2A
0B0A
0B5F
0C02
0C32
0BB3
0B4E
0BBF
0C77
0BF1
096E
05FF
0385
02DA
0340
038B
035D
031D
0323
035D
03AA
0418
0498
04D0
047E
03FB
03E5
0453
04A1
0449
03A2
036C
03C4
03F9
037F
02B6
0263
02B1
0320
034B
0351
036E
0385
0366
0341
0375
03F0
0424
03CB
035B
0361
03AE
039D
033B
0393
0579
084A
0A4C
0A81
09BF
09B2
0ADA
0C01
0BD5
0A91
0994
097F
098F
090C
08B8
09D1
0BBC
0BB0
0791
00D4
FB8E
FA6E
FC47
FDF2
FDD5
FCE5
FC92
FCE0
FCD6
FC14
FB3D
FAE9
FADE
FA8E
F9F1
F986
F9AD
FA51
FB0E
FB8E
FBD1
FC24
FC9E
FC8F
FAF2
F7D2
F4ED
F443
F5E1
F7A2
F77B
F5AD
F438
F454
F546
F5C5
F5B8
F5E0
F65F
F679
F5C9
F4FB
F4EC
F585
F5E1
F577
F4B2
F451
F47F
F4BF
F4A6
F450
F435
F4A2
F565
F5ED
F5E1
F595
F5BA
F66D
F6F4
F6A6
F5DF
F5A2
F636
F6A4
F5F3
F49F
F453
F619
F926
FBC4
FD00
FD2E
FD13
FD0E
FD26
FD5C
FD93
FD7A
FCF5
FC74
FC73
FCA2
FC1C
FADD
FAA9
FD99
038A
098B
0C7A
0C0E
0ABA
0AB4
0BC3
0C47
0B9D
0AC1
0AB3
0B2F
0B69
0B53
0B6C
0BA5
0B65
0AB4
0A7F
0B32
0BE6
0BA6
0AF8
0B2A
0C18
0BD1
090B
052E
02FA
034C
0458
0439
0334
02BF
033D
03AF
036F
0311
0354
03FA
044B
042B
041B
0449
0452
0408
03CF
03E8
03EE
0386
0314
0331
03A8
03AF
0315
0295
02BF
0325
0304
0272
0252
0307
03DC
03FC
038D
0359
0392
039F
0333
0309
0431
06C3
097C
0ADE
0A96
09B9
0986
0A1A
0A9A
0A77
0A29
0A5B
0AC2
0A59
0907
084A
096C
0B38
0A93
05E6
FF49
FA94
F98C
FAAE
FB97
FBA4
FBC9
FC88
FD2D
FD0A
FC77
FC34
FC50
FC4D
FC00
FBB5
FB89
FB42
FAD5
FA98
FAC7
FB25
FB6C
FBB7
FC16
FBDD
FA34
F76C
F52A
F4B0
F571
F5E2
F572
F4FA
F538
F5A2
F546
F446
F3AF
F3FA
F472
F465
F432
F493
F566
F5D3
F597
F55B
F5A1
F5EF
F59A
F4E2
F4AE
F53B
F5C1
F59D
F52A
F513
F555
F577
F57E
F5DB
F68A
F6DD
F66E
F5C4
F591
F5AF
F586
F55B
F650
F8D7
FBAC
FD18
FCBF
FBC9
FB72
FBFA
FCDA
FD6E
FD57
FCB9
FC46
FCA9
FD88
FDA0
FC82
FBFA
FE7C
0402
096A
0BB5
0B29
0A58
0ABC
0B6B
0B26
0A50
0A25
0AD5
0B72
0B91
0BCA
0C57
0C70
0BA6
0AF6
0B7A
0CA1
0CCF
0BA4
0A8D
0AC1
0B92
0B4D
0963
06DA
04D6
0386
02B2
0284
031A
03EC
0455
0463
047F
0494
0437
038D
035C
03F4
049B
0476
03B8
036F
0419
050F
056D
0525
04B9
0469
0410
039B
032D
02E3
02CC
02FC
0362
039C
0353
02B6
0256
0271
02AC
02A9
0293
02B8
02DF
02BD
02F3
04AE
07DE
0A9F
0B33
0A27
0991
0A53
0B1F
0AA3
0997
09B2
0AFD
0B97
0A77
0930
09C5
0B62
0AB1
05CF
FEF3
FA54
F9DF
FBB7
FCD1
FC2C
FB0C
FAC4
FB36
FB77
FB2D
FACD
FAD2
FB30
FB91
FBBE
FBB0
FB73
FB31
FB24
FB70
FBF9
FC86
FCE2
FCCE
FBF8
FA48
F834
F681
F58D
F50A
F48E
F441
F491
F560
F5EF
F5C5
F53D
F4E7
F4BE
F46E
F420
F45F
F532
F5D8
F5AD
F50B
F4C9
F504
F510
F4A6
F464
F4D6
F591
F5C3
F560
F51C
F561
F5E4
F63C
F669
F68C
F67F
F61D
F5B2
F5AB
F5CC
F56D
F499
F466
F5C5
F85C
FAF4
FC9E
FD21
FCBC
FC06
FBD9
FC99
FD7F
FD44
FBDA
FAE0
FBAF
FD51
FD8C
FC19
FB9B
FEAA
0496
0A0F
0CAF
0CD8
0C4B
0C00
0BDD
0BCB
0C03
0C6E
0C7F
0BFF
0B71
0B4D
0B48
0AE3
0A3F
09EB
0A10
0A64
0AC5
0B4A
0BAC
0B21
093F
06B6
04CF
0426
0436
0437
03F1
03A2
0369
033E
0347
03B5
0452
048E
0428
0383
033A
036E
03A8
036F
02E5
02B0
0337
0415
0476
03FD
032E
02DC
0333
038E
0359
02D0
0299
02BD
02AE
0246
023B
0309
03F6
03DB
02EC
02EC
0521
0892
0AE3
0AF2
09E2
0967
09BC
09EF
09A9
09B6
0A82
0B20
0A7F
0934
0908
0A5D
0AFC
0841
0267
FCC7
FA72
FB27
FC2D
FBB5
FA7C
FA1D
FACF
FB82
FBA0
FBA0
FBED
FC17
FBAC
FB33
FB85
FC5A
FC7E
FB99
FAED
FBA8
FCF9
FCC0
FA14
F667
F3F7
F3A0
F480
F556
F5AA
F5A4
F570
F51A
F4D0
F4C5
F4F5
F526
F52F
F503
F4B5
F488
F4C9
F566
F5DC
F5C7
F566
F548
F590
F5C9
F598
F542
F541
F58D
F5B1
F590
F591
F5EE
F643
F630
F5E6
F5BD
F593
F51E
F4C1
F56C
F785
FA37
FC26
FCB5
FC6D
FC37
FC7E
FD05
FD4E
FD08
FC79
FC6B
FD4F
FE5C
FE3D
FD0E
FCFA
001C
05DA
0B1D
0D50
0CB3
0B79
0B29
0B87
0BC4
0BB5
0B98
0B58
0ACA
0A3C
0A24
0A75
0ABA
0AC3
0AC4
0AD7
0AD6
0ACB
0B09
0B7E
0B42
0970
0670
03DC
02DF
031C
036C
034F
0322
0339
0379
03B8
0402
044F
0457
03EE
035C
0314
0315
02DF
022C
017B
019B
02AE
03EB
045D
03CC
02EF
02B2
0348
0402
0423
03C3
038B
03AF
03AE
0341
02FC
0382
0455
0449
034C
0308
0505
0887
0B12
0B3A
0A11
0977
09D3
0A35
0A31
0A5B
0AEE
0B11
0A23
091F
097F
0ACA
0A5C
065D
0053
FBDD
FAEB
FC09
FC87
FB92
FA8F
FAD8
FC11
FCE9
FCD8
FC6A
FC1E
FBB4
FADD
FA14
FA29
FB14
FBDA
FBC7
FB56
FB74
FC0F
FBE2
F9F4
F6F4
F4B4
F44E
F52D
F5ED
F5EB
F5AB
F5D3
F645
F664
F5FE
F594
F5AC
F61E
F657
F621
F5E4
F606
F64B
F62D
F5A9
F553
F588
F5EE
F5FE
F5C5
F5C3
F61B
F656
F617
F5A9
F590
F5C4
F5CC
F59C
F5BD
F661
F6DF
F68B
F5D5
F601
F7B8
FA48
FC52
FD15
FCDF
FC87
FC9F
FD13
FD62
FD32
FCCD
FCE5
FD8F
FDCC
FCC1
FB74
FC66
00D8
06FE
0B96
0D10
0C8C
0BF0
0BDE
0BDE
0BB2
0B99
0B86
0B12
0A78
0A9B
0BAA
0C77
0BEC
0A93
09DB
0A37
0AD4
0B0D
0B37
0B96
0B57
0976
066A
03FD
034B
03AC
03F5
03F5
0418
0440
03EA
0340
0307
037E
03E5
0390
02D5
028B
02CD
02EE
0295
0254
02CA
03AF
042E
03EC
034C
02D2
02B5
02DD
030A
0301
02D4
02DC
0339
0391
0384
0342
0352
03B4
03BF
0347
036C
056B
08B5
0B23
0B69
0A7E
09FF
0A19
09EE
097F
09DA
0B27
0BE2
0AE6
0969
0989
0AEA
0A6E
0609
FFBE
FB96
FB1A
FC29
FC33
FB2D
FAC2
FB86
FC45
FBF0
FB0C
FABD
FB1F
FB5F
FB20
FAEB
FB3E
FBC2
FBD5
FB72
FB36
FB96
FC36
FC32
FAF4
F8CC
F6AE
F56C
F516
F524
F521
F522
F567
F5C7
F5C7
F55A
F516
F56B
F5FA
F618
F5BC
F591
F601
F6A6
F6D5
F67B
F610
F5E1
F5CC
F5C0
F5F5
F66B
F6AF
F676
F62D
F678
F72F
F768
F6AA
F59F
F54F
F5CF
F63E
F603
F5A8
F62E
F7E8
FA24
FBE7
FCB5
FCCF
FCE8
FD77
FE2C
FE3A
FD6A
FCAC
FD1F
FE6D
FED4
FD64
FBD5
FD28
0233
084A
0BEC
0C4A
0B77
0B84
0C58
0C98
0BC7
0ABF
0A64
0AB2
0B38
0BC2
0C38
0C4E
0BE5
0B69
0B4D
0B5A
0B0E
0A8F
0AA0
0B65
0BBF
0A64
0780
04B3
0350
0330
0359
034A
0332
033E
0352
0364
0397
03E3
03EF
038E
030D
02E4
031D
0352
0341
031C
032A
035D
0373
0351
0308
02BE
02A5
02DD
033A
0363
034C
0354
03B0
03FF
03D0
0364
036E
03F4
0411
035F
0313
04C7
082A
0AE1
0B3C
0A1C
097E
09EE
0A5A
0A16
09CB
0A10
0A46
09BF
0938
09DC
0AD8
0974
0470
FE37
FA85
FA65
FB9B
FBCF
FB14
FAE4
FBB1
FC74
FC58
FBC4
FB7C
FB7C
FB40
FAC8
FA9D
FAF7
FB74
FB9C
FB6A
FB35
FB56
FBB9
FBB9
FA8B
F828
F5AF
F481
F4D8
F590
F588
F4EE
F4CA
F571
F61F
F632
F609
F633
F668
F5FA
F518
F4C3
F566
F629
F60B
F53E
F4D6
F548
F5DF
F5E4
F59E
F5C2
F653
F6AF
F687
F63E
F634
F63D
F60C
F5D6
F612
F6AB
F6DF
F629
F515
F4E1
F656
F8FF
FB81
FCAF
FC7B
FBF4
FC30
FD1A
FD94
FCF0
FC03
FC2A
FD58
FDE3
FCD9
FBF0
FE04
0386
096F
0C6B
0C48
0B85
0BE8
0CB7
0C89
0B98
0B3A
0BBA
0BF6
0B4B
0A9C
0AD7
0B71
0B5A
0AB0
0A83
0B15
0B7A
0B2B
0AF0
0B7C
0BDF
0A6B
0728
042B
0326
0383
039F
030B
02AC
0312
03BD
040D
040A
0400
03E2
0383
0310
02E5
02FF
0302
02DF
02EB
033D
0376
0362
0344
0339
02EE
0258
0218
0290
0324
0306
027A
0276
0324
0390
031D
0286
02B9
033D
02F9
0265
0374
06C9
0A4F
0BA0
0ADF
0A0D
0A33
0A93
0A67
0A14
0A18
0A02
0961
0902
09C9
0A7F
086C
02E5
FCEE
FA26
FADA
FC53
FC71
FBA1
FB43
FB9A
FBDF
FBAC
FB66
FB65
FB7C
FB79
FB8E
FBDD
FC1B
FBF9
FBAA
FB8E
FBC0
FC32
FCD1
FD0E
FBEA
F91C
F5F1
F44F
F4BC
F5EC
F659
F5E3
F575
F591
F5D2
F5E0
F600
F66B
F6AF
F65A
F5C9
F5B9
F62D
F66D
F612
F58B
F577
F5DB
F634
F621
F5C6
F588
F5A4
F607
F673
F69E
F662
F5E1
F573
F551
F570
F5AE
F5E0
F5C6
F54B
F505
F5F8
F868
FB23
FC88
FC42
FB9B
FBDF
FCD9
FD53
FCDB
FC4E
FC7A
FCD3
FC49
FB36
FBAD
FF56
0548
0A8B
0CC9
0C4C
0B2F
0AF6
0B5A
0B65
0B01
0AE9
0B56
0B9E
0B45
0AC7
0ADC
0B63
0B9B
0B4C
0AFF
0B16
0B33
0B02
0B02
0BC1
0C79
0B81
0878
052C
03B1
040D
0491
0421
0349
0308
035C
0383
032D
02D3
02DA
0313
032A
0330
034F
0357
030D
029F
0275
02A2
02EA
0324
0352
0370
0370
0362
035B
0350
0328
02FB
0300
033B
0367
0360
036E
03B9
03CA
0328
0281
034D
05EF
08E1
0A5A
0A4B
0A0F
0A85
0B3C
0B76
0B2A
0AB1
0A25
09A9
09CA
0A97
0A84
0788
01EE
FCEF
FB7A
FD06
FE83
FE14
FCC5
FC7F
FD7C
FE6C
FE67
FDD6
FD6D
FD3C
FD07
FCE8
FD09
FD2A
FD06
FCD5
FCE5
FD0F
FD0F
FD22
FDB5
FE90
FEE6
FE66
FDB5
FD96
FDE1
FDD0
FD30
FCAB
FCCE
FD54
FDC4
FE19
FE66
FE62
FDDB
FD50
FD68
FDFD
FE38
FDBA
FD1B
FD0E
FD66
FD6C
FCF3
FC92
FCBB
FD2C
FD80
FDBB
FDF1
FDE8
FD7A
FD0E
FD14
FD60
FD7C
FD68
FD8B
FDDA
FDBD
FCF8
FC40
FC61
FD15
FD67
FD2B
FD2F
FDD1
FE48
FDED
FD63
FD89
FDE1
FD35
FBDB
FC2B
FFDC
0593
09F4
0B1F
0A54
09E3
0A77
0B0B
0ADF
0A65
0A54
0AA1
0AC0
0A7D
0A2C
0A31
0A85
0AC5
0AA6
0A50
0A20
0A3B
0A5E
0A34
09D3
09B1
0A0E
0A8F
0AB7
0A9E
0ABE
0B10
0AF8
0A4C
09BB
09C3
09DA
0952
08B0
0928
0A8C
0AA4
0777
01ED
FD42
FBB4
FC73
FD38
FD04
FC91
FC9B
FCD6
FCB0
FC4B
FC35
FC89
FCD6
FCC4
FC8C
FC93
FCDE
FD15
FD01
FCC5
FCA0
FC9F
FCA2
FC8A
FC6B
FC81
FCDC
FD37
FD4B
FD4A
FD8E
FDE4
FDAB
FCDB
FC64
FCF4
FDC1
FD67
FC14
FC12
FF5A
04EF
0987
0AEF
0A13
094A
0986
09EF
09C5
097B
09CA
0A7C
0AB5
0A29
0979
0952
099A
09C1
0992
096B
09A0
0A05
0A27
09E0
097E
095E
0977
095E
08E1
086D
0886
0904
093B
08FD
08E1
0945
0990
090F
0842
086E
099E
09C7
06D2
0158
FC72
FA95
FB34
FC03
FBCB
FB44
FB68
FC01
FC36
FBE1
FBB0
FC19
FCB4
FCC9
FC47
FBC3
FBA9
FBC7
FBAE
FB56
FB21
FB5E
FBEC
FC64
FC86
FC6A
FC38
FBF2
FBAA
FBB7
FC54
FD08
FD08
FC54
FBF3
FC97
FD6E
FD04
FB7B
FB1A
FDFE
036F
0844
0A0C
0954
0873
08C1
0997
09CB
0945
08D3
08EA
0926
08FD
0888
085A
08B1
091B
091C
08E0
08F7
0978
09BD
0937
0845
07D5
083D
08C6
08AA
0827
0814
088F
08D2
0871
080C
0845
08B0
0880
07FD
084A
0970
098B
06A3
013D
FC46
FA30
FAAC
FB91
FB76
FACD
FAA6
FB34
FBB9
FB91
FAF1
FA9A
FAF0
FB7F
FB93
FB26
FAEC
FB60
FC1A
FC51
FBE2
FB70
FB7B
FBB6
FB95
FB2F
FB0E
FB3F
FB43
FB01
FB0F
FBA7
FC0D
FBAE
FB27
FB6B
FC20
FBE8
FAA1
FA63
FD59
02E3
07D8
09CE
094E
0878
085E
0889
0877
086B
08B4
090E
0910
08CB
08A4
08BA
08CA
089E
0855
0825
0818
081F
0837
0857
0855
081B
07D5
07B6
07D1
081F
0874
086C
07CB
0717
073B
083E
08E2
0828
06F4
0727
08E8
099F
06AE
00D2
FBBA
FA0C
FADD
FB91
FB2E
FAC4
FB26
FBA4
FB50
FA79
FA33
FACF
FB7F
FB7E
FAFE
FAAC
FABF
FAE5
FADC
FABB
FAB1
FAD6
FB22
FB69
FB76
FB50
FB30
FB25
FAFF
FAC1
FAC3
FB2A
FB87
FB61
FB0A
FB3E
FBEA
FBF7
FAED
FA64
FCB2
01EC
0731
098F
08FF
07D7
07C0
0848
0844
07A4
0751
07C5
0878
08B5
087F
0853
086D
089C
08A3
087E
084F
0841
0863
0883
085A
07FE
07D4
07F6
0801
07B4
0757
0748
0763
074A
0710
071A
0757
0735
06AE
06C3
07FF
08D7
06C8
0181
FBF0
F945
F99E
FA89
FA4C
F988
F996
FA74
FB01
FAB6
FA2E
FA05
FA08
F9D2
F99E
F9DF
FA6B
FAA7
FA61
FA00
F9E9
FA22
FA65
FA66
FA16
F9D0
FA07
FAAE
FB28
FB0B
FAAC
FAA0
FADB
FACC
FA6B
FA78
FB2E
FB6F
FA48
F926
FAEA
0041
0615
08C6
081A
06E2
0720
080C
07FF
0709
068D
0704
076C
070A
0683
06B9
0764
07A2
0759
072B
075C
0794
079D
07A5
07CF
07F9
07FE
07E4
07B8
077F
0746
0723
070A
06CB
0675
066C
06DC
0746
0733
0725
07CF
084C
066E
0191
FC31
F985
FA07
FB6B
FBA8
FAF4
FA8B
FAA9
FA9D
FA4B
FA60
FAFA
FB3E
FAAF
FA0D
FA1D
FA6D
FA23
F96F
F93D
F9C4
FA51
FA63
FA41
FA5E
FAA9
FAC9
FAA3
FA6F
FA5F
FA76
FAB6
FB07
FB10
FAA2
FA2F
FA3E
FA66
F9E7
F983
FB68
0052
05CC
087C
07CC
0634
05FA
06EA
077A
0733
06E7
0708
0711
06B9
0696
06FE
0742
06D3
065A
06BF
07A8
07F8
076C
06D6
06D0
0713
0716
06D9
06B3
06BF
06D5
06DA
06D4
06AE
0659
0618
062E
064C
060D
05FD
06E7
07DD
0658
015F
FB85
F878
F8F7
FA76
FA94
F99A
F930
F9B6
FA1B
F9D7
F9A3
F9FE
FA3E
F9C7
F934
F959
F9E8
FA0C
F9C6
F9B9
F9FB
FA0D
F9D9
F9DE
FA4D
FAA5
FA6E
F9EC
F9C0
FA0F
FA68
FA7A
FA5A
FA24
F9E7
F9F9
FA86
FAC7
F9D7
F8B3
FA04
FEE3
04C3
07EB
0790
0639
0641
074D
07AB
0704
068C
06E7
074E
070F
06BA
070C
079B
0790
06FC
0698
0699
06A8
06B2
06EA
0724
06FA
067B
0636
0676
06D8
06D8
066F
05FC
05AE
0588
05B4
063E
069F
0651
05E8
0667
072E
05E0
015D
FBD9
F8B7
F8C8
F9E1
F9E7
F910
F8C3
F951
F9CB
F9A5
F96E
F9A8
F9EA
F9B0
F949
F93D
F969
F95B
F92B
F933
F962
F96C
F961
F97E
F9B4
F9CB
F9CC
F9D7
F9CD
F98D
F963
F9C3
FA70
FA88
F9D1
F95C
FA11
FAF6
FA6E
F933
FA46
FF0F
04E9
07FD
07A2
066A
0672
073A
0754
06B3
0655
0685
0697
0646
0632
06A5
06F0
0694
062B
0667
06E6
06E9
0693
0686
06CE
06FD
0700
0712
071E
06D8
066C
0658
069A
068C
05ED
0577
05CF
0653
060B
058A
063F
0793
06A0
01D9
FBBE
F83F
F845
F959
F94F
F89C
F8B1
F98B
F9F7
F999
F94E
F997
F9D1
F97A
F92A
F97D
F9F6
F9DB
F97B
F994
FA0A
FA1D
F9AD
F952
F95B
F973
F949
F90A
F902
F92C
F95D
F98D
F9B0
F985
F906
F8CD
F947
F9A9
F8DF
F7C5
F900
FDB5
037B
06C8
06D6
05E1
05EB
06AB
06DB
0652
05F9
062C
0647
05EA
05A6
0604
0694
06A2
064B
0626
0653
0683
0697
06A3
0692
0659
062B
062D
0623
05E1
05AC
05D1
0605
05C3
053B
054F
063F
06F5
067E
05B6
0623
072A
0601
0151
FB8E
F86F
F8C4
FA1F
FA3F
F954
F8C0
F8EA
F917
F8D8
F88A
F87E
F86E
F82E
F823
F88F
F902
F903
F8CE
F8CF
F8E5
F8C1
F88A
F88D
F8AA
F89E
F888
F8AD
F8EB
F8F1
F8EA
F94C
F9F2
FA04
F933
F87A
F8D3
F98B
F933
F847
F95B
FDC5
0363
06DF
075E
06B4
0686
06A9
066A
060D
0645
06E1
0700
067D
0622
065D
0691
0630
05A9
059F
05EB
0607
05FB
0610
0628
0611
0613
067F
06F1
06C3
0617
05C0
060B
0649
05E9
056E
059A
0605
05B5
04FB
0532
062E
0580
0178
FBE2
F848
F7F2
F8FF
F93E
F894
F832
F88E
F904
F91F
F915
F909
F8B8
F843
F852
F8F9
F955
F8E4
F868
F8A9
F92F
F91D
F8AE
F8C3
F953
F970
F8E6
F8B0
F95F
F9F4
F977
F919
FB46
003B
0512
06FB
0655
057D
05A7
0624
063C
062F
064C
063C
05BC
0547
0579
0614
0655
0617
05EF
0614
060F
05C4
05C7
0643
0673
05E6
0574
05F1
06B9
0697
05CE
05D3
06C2
0662
02B2
FCDC
F86A
F76D
F894
F960
F913
F894
F87D
F88A
F88E
F8CB
F942
F97F
F94D
F90A
F90F
F928
F8FC
F8A7
F88E
F8AE
F8B2
F89D
F8C5
F909
F8D9
F84C
F846
F8FF
F953
F884
F80F
FA62
FFB2
051C
0793
06FA
05B0
0576
05DA
05BD
052D
04F4
053E
0586
0590
0598
05B3
05B7
05A4
05A5
05B8
05AE
0598
05B5
05E8
05AF
04FC
049D
0534
0607
05E4
0511
0519
061F
05C9
020B
FC3E
F810
F779
F8DF
F990
F8E6
F83A
F871
F8EE
F8EF
F8C6
F903
F961
F94B
F8DC
F899
F897
F897
F899
F8BC
F8C9
F886
F847
F88A
F911
F90B
F86A
F83A
F909
F9A7
F8CC
F7B5
F972
FEDB
04CC
0788
06E0
05A8
05C7
0682
0684
0602
0601
0680
0692
0602
05A6
05E5
0615
05BF
0579
05C4
060A
059E
04FA
04FB
0576
059A
055B
0564
05C5
05C1
0537
0524
05DC
058F
021A
FC51
F7D3
F6F4
F837
F8CA
F833
F803
F8DC
F987
F909
F811
F7D8
F86E
F8EE
F8E7
F8BB
F8B8
F8A6
F873
F872
F8A2
F883
F812
F80A
F8A5
F908
F8A2
F842
F8BE
F963
F902
F85D
F9EC
FEB1
0442
072A
06C9
059F
05C4
069C
0695
05C1
0564
05D9
064A
062F
05E4
05D2
05DE
05DC
05E1
05F3
05E2
05A4
0594
05E3
0612
05A0
04F8
04F4
0576
0582
050D
0548
0661
063C
02CF
FD28
F8B4
F779
F83C
F899
F7F4
F77C
F7E5
F87A
F874
F825
F82F
F878
F891
F888
F899
F899
F85F
F84C
F8AF
F912
F8DD
F863
F879
F922
F96E
F8F1
F884
F8E7
F952
F8A5
F7DC
F99C
FEAF
0449
0702
0694
0584
059C
064E
065B
05CB
0587
05DF
0653
0685
069F
06AC
0669
05EE
05C3
05F4
05D7
0537
04E2
056A
0614
05EF
0549
051C
0570
055F
04D7
04FB
0618
0629
02D9
FCE5
F800
F6D0
F828
F919
F894
F7D8
F7F6
F87E
F89B
F857
F83D
F862
F878
F86C
F882
F8C5
F8EC
F8DE
F8CF
F8C3
F882
F836
F85E
F8E9
F90F
F89C
F875
F920
F996
F8B6
F791
F8E5
FDC4
03B6
0713
06EC
0595
0562
0631
0696
063A
05ED
0610
0628
05E7
05A0
05A9
05D9
05E6
05CC
05AC
0590
057B
058C
05B9
05A6
051F
04A7
04D3
0542
050E
046B
04AE
0603
063A
0311
FD59
F87E
F6F4
F7E4
F8CE
F88F
F7F8
F7F5
F84B
F872
F885
F8C4
F8DD
F880
F810
F81B
F872
F884
F84B
F834
F854
F85B
F843
F86A
F8D9
F907
F8B5
F888
F909
F97D
F8DA
F800
F977
FE36
03C8
06C5
068A
0553
051C
05BA
060F
05EB
05E6
0619
0601
0598
058D
0619
0682
0634
05A4
0571
0572
053F
0512
0548
0590
0563
050A
053D
05DD
05EA
0528
04C3
057E
05CF
0347
FDFB
F920
F77B
F862
F934
F8CE
F82A
F836
F889
F876
F839
F863
F8C2
F8AA
F81B
F7D4
F82F
F8A9
F8BD
F894
F86B
F81B
F7B0
F7BC
F875
F91A
F8FB
F88D
F899
F8D5
F865
F7C6
F909
FD59
02E1
0653
067F
054A
04F0
0583
05CF
058A
0570
05BC
05DE
058B
0541
056E
05D6
0604
05F3
05DD
05BE
0571
0526
0531
0570
0570
053C
0557
05AD
0589
04F0
0504
061A
0662
03AC
FE5B
F96F
F767
F7DD
F8AD
F8B3
F87A
F89E
F8BE
F869
F806
F81E
F86C
F875
F860
F896
F8E9
F8E8
F8AE
F8A7
F8C3
F891
F81D
F802
F86C
F8AC
F84C
F7FA
F882
F942
F8E8
F7F5
F8F5
FD43
02CA
0623
065F
0569
0526
0584
0591
053C
0530
0587
05AB
0569
0541
056B
0573
0526
0516
058E
05EC
059F
0526
053A
0594
0581
0523
0537
05B0
05A0
04DF
04AB
05C3
0674
041B
FEB3
F978
F757
F7DF
F89C
F86B
F814
F853
F8BB
F8BE
F891
F897
F8A2
F857
F7F6
F80D
F884
F8AE
F85F
F82B
F85E
F882
F850
F84C
F8BE
F903
F89B
F838
F8B6
F97B
F930
F823
F8B4
FC90
0221
05F1
066E
054F
04F2
05A3
0628
05F6
059D
058B
058C
056F
0564
0583
0594
0578
0560
056B
0567
0533
0517
0557
059B
0561
04F0
050F
05A6
05B5
050D
04F3
060E
069F
0426
FEB2
F959
F706
F791
F896
F87B
F7C1
F778
F7AF
F7DE
F7F5
F831
F86C
F861
F838
F846
F876
F882
F87F
F8A6
F8C8
F88B
F823
F82B
F8AC
F8DD
F856
F7F1
F89B
F994
F93B
F7D4
F819
FBFA
01CF
05F3
06C2
05D1
0559
05C5
0621
05FD
05DC
060B
0621
05D5
058D
05A4
05D3
05C6
05AB
05B5
059B
053F
0525
05A2
0619
05C6
0507
04E8
057F
05A9
04E4
0464
0546
062D
0446
FF15
F9B3
F769
F813
F910
F8DE
F849
F866
F8E3
F8DA
F84E
F7FF
F82B
F84F
F825
F805
F833
F868
F87D
F8BB
F92A
F93C
F8C0
F865
F8AB
F907
F8CF
F874
F8C6
F953
F8CD
F769
F79E
FB73
0175
05C7
066A
0527
04C3
05AE
066C
0641
05DF
05E0
05F1
05B2
0574
0598
05E2
05D0
056C
052F
053C
0544
0532
054E
058B
057D
0538
055C
05E6
05EB
052F
04F1
060E
06EC
04CE
FF59
F99A
F6EE
F781
F8C9
F8EA
F866
F85F
F8AE
F88C
F810
F7EB
F82C
F84E
F832
F836
F874
F8A6
F8B8
F8E2
F91A
F901
F888
F837
F866
F89C
F859
F829
F8DD
F9D1
F961
F7B7
F79B
FB43
012D
0582
0654
0537
04AF
054A
05EA
05E5
05BD
05E6
0608
05D7
05B0
05DC
05F3
059F
054E
0571
05A8
0567
04F5
04EC
0536
0548
052B
0570
05FC
05E3
04EE
047A
05A1
06E4
0541
0011
FA67
F7B2
F809
F8E3
F8A1
F7EA
F7D7
F846
F879
F850
F83D
F854
F842
F80D
F828
F8AA
F909
F8FE
F8EB
F912
F913
F8B4
F870
F899
F8AE
F838
F7D0
F83F
F8FA
F8AA
F77C
F7C7
FB81
0169
05F3
0713
0616
0571
05D6
0654
0652
062E
062F
060F
05AC
0564
0582
05C4
05CA
059A
0581
058B
0580
055E
055C
0573
0561
0539
055B
05A3
0571
04D2
04DC
0604
06B1
049C
FFA6
FA6A
F7A7
F79E
F86C
F88E
F839
F83E
F89F
F8C6
F88E
F858
F85C
F879
F88F
F897
F87C
F83C
F815
F848
F8B1
F8F0
F8EC
F8DA
F8D0
F898
F83C
F84D
F918
F9C6
F92D
F7BE
F7C9
FB1B
00AF
0579
0764
06E9
05DF
056A
0566
055B
0540
0552
058D
05B7
05BB
05AE
05A1
0591
0584
0582
058C
05A3
05B4
0589
051A
04EC
059E
06AF
0644
02D4
FD3F
F88B
F71B
F85C
F9AD
F95F
F82F
F7B2
F82D
F8A2
F881
F84F
F8A1
F921
F91A
F888
F827
F869
F8D9
F8CE
F865
F85D
F8F8
F974
F8F9
F7FE
F854
FB76
00B8
0572
074B
0663
04F6
04E2
05EE
06A8
0664
05D0
05B8
05E8
05B9
0539
051B
0592
05E4
0583
04F6
0522
05E5
0625
056F
04CD
0574
06C9
0681
0307
FD83
F8FA
F772
F840
F935
F905
F83A
F7F1
F858
F8A9
F86A
F810
F841
F8CF
F8F4
F876
F803
F83B
F8C8
F8E0
F87C
F870
F91E
F99E
F8DE
F77E
F7CA
FB54
00E2
055B
06BD
05D9
04FE
0564
0652
068E
05F1
0555
054B
0589
0596
058B
05CD
0649
066F
0602
0584
058C
05E7
05D6
053E
050D
0604
0732
0661
026C
FCD4
F8A3
F796
F8B7
F9C0
F98A
F8C1
F878
F8BD
F8D4
F868
F7FD
F81C
F890
F8C2
F88B
F865
F8AB
F915
F925
F8E1
F8C7
F8FB
F8EB
F82E
F795
F8D5
FCBD
01E9
05BB
06BA
05CD
0506
0563
0623
062C
0580
050A
0547
05C0
05DA
05B1
05CF
0641
0670
05FF
055F
053C
058B
05A5
0559
0557
0627
06E4
05A4
017D
FBEE
F7D2
F6C5
F7D6
F8DC
F8CB
F854
F87B
F91C
F948
F8AE
F811
F83B
F8F3
F951
F8FB
F884
F892
F900
F932
F907
F8F3
F920
F8FB
F815
F74F
F87F
FC89
01FD
0610
0729
0638
056A
05CF
06A5
06CA
063F
05E5
0625
0671
0632
05AC
0587
05C4
05BF
0530
04AF
04D6
0558
0567
04FE
0515
0634
072E
05EA
01A1
FC13
F81F
F72B
F827
F903
F8C7
F81E
F801
F876
F8BE
F875
F80C
F819
F886
F8C8
F8BB
F8C6
F925
F972
F940
F8DE
F900
F99B
F9B2
F8B0
F7B3
F8E0
FD13
0294
0680
0770
0674
0593
05B6
0638
0633
05A7
053B
054C
058C
059D
0598
05C7
060F
0607
0599
053D
0555
058F
054F
04B2
04AD
05BF
06BD
058A
0155
FBD0
F7D8
F6D9
F7D0
F8BF
F8BB
F85C
F876
F8F5
F92B
F8D2
F861
F85A
F8AF
F8FA
F919
F939
F95D
F93E
F8C3
F86B
F8C9
F994
F9B3
F8A1
F79C
F8D8
FD27
02B7
0692
0759
064D
058E
05DC
0651
0602
0541
04FB
0564
05D2
05C4
058D
05B4
0615
060B
056C
04E2
0504
057C
0578
04EF
04E1
05EB
06EA
05B0
015E
FBC5
F7ED
F745
F882
F95E
F902
F862
F882
F916
F924
F884
F81B
F897
F97F
F9D6
F964
F8DD
F8D8
F91B
F925
F90A
F93C
F990
F930
F7E9
F729
F901
FDD2
0360
06AB
06B8
053C
0482
0512
05B8
057B
04DF
04FA
05D9
0670
0610
0553
053C
05D1
0621
05A7
04FD
04F1
055E
057A
053C
058C
06C6
0776
0572
006E
FADB
F7BF
F7D0
F921
F986
F8C7
F839
F8A5
F957
F93C
F86B
F7F3
F876
F95E
F9BB
F96B
F917
F92F
F95F
F933
F8DC
F8E4
F92F
F8E9
F7D5
F750
F950
FE19
0365
0653
0630
04EC
04C1
05DC
06B9
065B
0578
0543
05C5
0600
0580
04FA
053C
05FD
0644
05BB
0519
050C
054A
0526
04C6
0515
0650
0704
052E
0079
FB07
F7B2
F773
F8B9
F954
F8B1
F7F7
F832
F8FE
F939
F89A
F801
F82E
F8C1
F8DA
F871
F85E
F909
F9BB
F99A
F8F0
F8BE
F92D
F92E
F822
F764
F943
FE44
0408
0765
0778
0627
05B0
0659
06CE
0638
0545
0509
0587
05DA
058C
0531
0572
0610
0638
05BB
0557
05A7
063A
062F
058E
0564
062F
06A0
0497
FFA3
FA09
F6D8
F708
F8C0
F991
F8E5
F809
F821
F8D4
F91E
F8CD
F89C
F8F6
F950
F909
F872
F86B
F913
F98A
F928
F879
F873
F8FE
F8FD
F80D
F7AA
F9E4
FEE4
0441
0727
06F9
0594
050A
05A1
0627
05D4
0534
0536
05D9
0640
05ED
0561
0555
05AC
05AD
052D
04DF
0551
05FF
05FD
055F
0544
0627
06A2
049A
FFC5
FA7A
F792
F7B5
F913
F9A2
F917
F893
F8DB
F97C
F9A2
F939
F8DE
F8E7
F901
F8C9
F876
F887
F8F9
F934
F8EB
F89E
F8EF
F997
F98C
F88C
F813
FA21
FEEC
0424
0704
06E4
057B
04C9
052B
05AD
05A6
056F
0588
05BD
058C
0518
0511
05B2
0648
060B
0539
04D8
0565
062A
063B
05C4
05CF
0694
0692
03ED
FEC9
F9B2
F757
F801
F997
FA06
F92F
F863
F86F
F8D3
F8D4
F892
F8AF
F932
F965
F8E4
F841
F84B
F8F6
F969
F92F
F8D4
F90B
F987
F94E
F84B
F812
FA7E
FF78
048F
0714
069A
051C
04BE
05BF
06BB
069C
05CA
055D
05B6
0645
0677
065E
063B
05FA
056E
04F4
0530
0614
06A2
0619
0516
04FB
0600
0666
0422
FF3A
FA1C
F75D
F76C
F8A3
F948
F913
F8BD
F8AF
F8A4
F863
F842
F8AA
F95A
F99C
F933
F8AE
F8A7
F8EF
F8E2
F86D
F847
F8E5
F998
F954
F85E
F8A8
FBDE
013D
05E1
0782
0691
055D
056E
063B
066D
05CA
054F
05A8
0653
0674
0607
05C9
0613
066B
0650
0602
0611
065F
0621
0510
042D
04B4
0649
06B7
0402
FEB4
F9B0
F78B
F83E
F9A0
F9DB
F90B
F866
F86E
F891
F84E
F80E
F86E
F92E
F974
F903
F89B
F8ED
F997
F9AA
F8FD
F871
F8AD
F924
F8DC
F81C
F89A
FBB2
00A0
04ED
06B9
0659
05A4
05CE
0661
064F
058C
051A
059A
0671
069E
0614
05AF
05E9
0630
05D5
0535
0544
060A
066A
05B6
04E4
0558
06B5
06B2
0389
FE32
F9A2
F7EC
F87F
F953
F93F
F8BD
F8B0
F915
F934
F8C8
F85A
F887
F920
F964
F904
F88E
F8A5
F913
F918
F896
F858
F8EB
F99C
F951
F854
F8A1
FBCD
00EF
0530
06A2
05FC
0557
05BA
066B
0665
05C5
056F
05D4
0675
06A9
0667
0621
0606
05D6
0577
0553
05D5
06A5
06D0
05F7
0508
0547
0676
0678
036E
FE14
F973
F7DE
F8C3
F9C5
F98B
F8C5
F89E
F908
F917
F889
F82D
F8A6
F977
F9B1
F93F
F8E8
F929
F98A
F958
F8A8
F84F
F8C5
F965
F925
F834
F869
FB8A
010E
061C
0824
0744
05C4
0566
05D2
05CB
0540
0545
0641
071E
06BE
058D
04E5
053B
05B8
0596
052B
0537
05B2
05E3
058D
056D
0625
06FA
0629
02C0
FDD2
F9BF
F824
F892
F940
F8FC
F844
F84B
F932
F9E3
F99A
F8F7
F903
F9AA
F9E7
F956
F8D8
F948
FA2D
FA58
F9A1
F91E
F979
F9DB
F93A
F83B
F8E0
FC4C
014F
0573
0721
06B9
05C2
056B
05C0
0611
05E5
0575
054E
0593
05CA
0585
0513
051E
05A5
05E0
0560
04DA
0533
0602
0595
02B8
FE31
FA29
F83B
F83E
F8E0
F92D
F935
F970
F9DE
F9F8
F96E
F8B0
F88A
F92C
F9D6
F9C1
F932
F92A
F9EF
FA77
F9BF
F87F
F8D2
FC0B
0119
0566
0732
06E1
0619
05EB
0625
0617
05A4
055F
05BD
066B
069A
05FA
053B
053D
05E9
0644
05D5
056A
05F8
06F4
0668
0305
FDCB
F957
F780
F7ED
F8E7
F934
F8EC
F8C4
F90B
F970
F98C
F96B
F972
F9BF
F9D7
F950
F8A4
F8DB
FA13
FAF2
FA1C
F83C
F7EC
FB18
00BE
05AF
0798
06E9
05C1
0585
05F5
0634
05FC
05BC
05D9
0638
0664
062A
05D4
05C2
05DD
05A6
0504
04AB
0550
0664
0605
02CF
FDA8
F948
F7BD
F898
F9D5
FA11
F991
F942
F969
F988
F939
F8BD
F89B
F8F1
F953
F959
F930
F957
F9E9
FA4B
F9D4
F8EC
F92C
FBFA
00E2
0595
07E4
079F
065F
05C1
0603
065B
0631
05C5
05B1
061A
0688
0688
063F
0625
0659
0666
05F2
0562
057E
062E
05FD
0365
FEB4
FA2C
F7F0
F80D
F8D0
F8D4
F849
F82F
F8DE
F9A2
F9B1
F91C
F8A3
F8C5
F939
F961
F915
F8D0
F90A
F981
F96F
F8B6
F8A0
FAE3
FF9F
04B5
0789
0774
061D
057E
05FC
0694
0686
063A
066C
070A
074B
06CF
061C
05EC
0639
0655
05E1
0569
05C4
06C9
06EC
0490
FFD4
FAE3
F81F
F810
F931
F9BA
F94F
F8E5
F938
F9E1
F9F2
F934
F85B
F823
F880
F8DE
F8F1
F904
F961
F9AD
F93D
F838
F813
FA68
FF20
040F
06CD
06D7
05C7
0562
05E3
0646
05F3
057D
05BC
0691
0713
06BD
060C
05D1
062C
0679
062D
05A1
05AA
066A
06A3
04AB
0034
FB10
F7DC
F7B4
F950
FA82
FA5C
F9B1
F994
F9F6
FA04
F977
F8F5
F90C
F968
F949
F89C
F820
F85E
F8DF
F8CA
F83B
F891
FB30
FFE4
04B2
076A
077B
063B
0575
05C3
065B
0654
05C4
0579
05D7
065F
066A
061B
061E
06A0
06EE
0669
058F
0588
068B
070F
051D
0079
FB3C
F808
F7BB
F8F5
F9CA
F996
F918
F91E
F98A
F9AD
F947
F8CE
F8BB
F8EC
F8EB
F8AF
F8BA
F957
F9F9
F9B9
F8A1
F829
FA0E
FE77
037F
06C0
0760
0683
05E1
061B
0692
068C
0621
05ED
0627
0661
0630
05C8
05B8
061B
0661
0602
055B
0566
0666
0711
0583
014A
FC38
F8E8
F85C
F947
F9BA
F922
F878
F8AC
F970
F9CE
F96D
F8E7
F8DA
F923
F93C
F917
F939
F9E4
FA79
FA09
F8A5
F7DD
F993
FE16
0383
0738
0805
06FD
0607
05F2
061B
05C6
0540
0559
061B
069E
0641
0596
05A5
0684
071D
06A0
05B3
05BA
06F2
07AB
05CE
011C
FBAF
F82E
F78E
F894
F963
F93E
F8C6
F8CB
F94C
F9A2
F972
F90E
F8F4
F92C
F955
F94B
F961
F9E1
FA67
FA25
F906
F854
F9D3
FDF9
031C
06B7
0798
06B8
05EA
05FA
064A
0621
05C6
060B
0702
07BC
075E
0632
0551
055D
05D9
05E3
056F
0555
061D
06DB
05B6
01C3
FC5B
F849
F751
F8A6
F9F6
F9DA
F8F2
F891
F8F8
F94C
F90E
F8D6
F95B
FA3F
FA77
F9BF
F90D
F944
F9EE
F9CB
F896
F7CB
F955
FD99
02D8
0693
0792
06B9
05E6
061F
06DB
0704
066A
05E9
0631
06CF
06CC
060B
0578
05BB
063F
0612
0559
0548
0669
0770
0647
023C
FCEF
F8F1
F7A2
F860
F989
F9F8
F9B1
F95A
F95F
F98E
F97D
F926
F8EA
F8FD
F91A
F8EE
F8B0
F8DB
F96C
F9A7
F91A
F897
F9D7
FDAE
02D8
06D9
081F
0737
05EF
0586
05D0
05FD
05CD
05CB
0668
073E
0778
06E0
0626
05FA
062A
05FE
055C
051B
05DF
06CD
05F8
0259
FD2C
F90F
F7B4
F895
F9CC
F9FD
F949
F8AD
F8C1
F93D
F986
F971
F94E
F95C
F97D
F981
F992
F9FA
FA84
FA68
F94E
F841
F92B
FCF5
0241
0660
07B0
06E5
05FA
0618
06C1
06E1
064D
05D5
0616
06A4
06A3
05F2
0562
05A6
0667
06AE
062E
05BF
063D
0715
0678
032D
FE1A
F9B1
F7CE
F847
F96B
F9C4
F932
F893
F891
F8FD
F93B
F911
F8D9
F8EC
F92A
F934
F918
F958
FA0C
FA64
F996
F85B
F8DA
FC78
01F8
0655
07A2
06BD
05F0
0655
070C
06E0
05F5
0573
05F7
06E5
074C
06EF
0660
062B
0646
0642
05FF
05F2
0687
0734
0669
02F8
FDA5
F909
F761
F86C
F9D5
F9CA
F8BE
F851
F90D
F9D3
F98A
F892
F831
F8DC
F9B8
F9D7
F96A
F952
F9CD
FA13
F97B
F8B0
F967
FCB3
01AD
05ED
078F
06CF
059B
058E
0683
073A
0704
0678
0679
0701
0742
06CF
062F
061A
0671
0678
05EF
0590
0618
0706
06A4
03A1
FEA1
FA08
F7EE
F84B
F94B
F95C
F8A2
F84E
F8E7
F9A9
F9A7
F904
F8A9
F8F7
F958
F937
F8EC
F93D
FA21
FA8F
F9C5
F87A
F893
FB75
0088
056E
07E2
0793
0635
05B7
0672
0730
06E4
05FD
05BA
0677
073A
071D
0674
0632
067E
0692
0606
0591
060A
06F6
0697
03A9
FEE0
FA72
F83A
F856
F96B
F9FF
F99D
F8E5
F8A4
F8F9
F95D
F975
F96D
F98B
F9A1
F95E
F8F9
F917
F9DD
FA69
F9C8
F872
F862
FB35
0050
0525
0774
072B
0614
05DB
0698
072F
06D8
0609
05BE
0634
06BA
06B9
0670
066A
0691
064D
058E
053F
062E
07AC
07B9
04DC
FFB5
FA9E
F7C7
F7A6
F8FA
FA0D
FA13
F98C
F95D
F9AE
F9D4
F96A
F8EF
F917
F9B7
F9EE
F973
F91A
F99C
FA4E
F9D4
F851
F7F6
FAC7
0027
0531
077B
070F
05CB
0559
05EE
06AF
06D5
0667
0600
0611
0664
0667
05F8
05AB
0604
0696
0686
05EE
05F4
0707
0794
0575
0095
FB7E
F8D9
F8E7
F9B9
F9AE
F901
F8D9
F980
FA23
FA0B
F976
F92E
F982
F9F2
F9C9
F906
F889
F90A
F9FB
F9F0
F885
F77C
F957
FE88
0486
0807
0815
0693
05D3
0645
06C4
0682
05F0
05E1
0669
06DC
06BF
065A
0652
06C3
06FF
0672
059C
05B8
0710
07F6
060F
00F2
FB1D
F7D3
F7FF
F99D
FA3F
F975
F883
F863
F8CE
F90E
F900
F8FF
F937
F96C
F960
F932
F93A
F999
F9FE
F9E0
F927
F8BD
FA36
FE4F
039C
075C
0805
06C0
05F3
0695
0784
0767
0678
05FD
067C
0722
070C
0675
0635
0674
067F
05F6
0585
060E
073F
077A
0548
00DC
FC16
F8F4
F818
F89F
F94A
F977
F947
F910
F8FB
F8F5
F8E0
F8C6
F8D9
F92E
F980
F976
F928
F921
F99C
F9F3
F966
F895
F994
FDB1
035B
0743
07C1
066E
05E0
06B0
0780
075E
06E5
06E3
0703
0692
05E4
05E3
0672
0689
060B
0618
06E2
066C
02CF
FD33
F90B
F849
F97C
FA1B
F993
F91D
F956
F97A
F914
F8DB
F952
F9B1
F93B
F8B1
F92A
FA0F
F9CA
F899
F922
FD45
033B
0734
078B
062C
059B
0619
0664
062E
0645
06D2
06F7
0665
0612
06AD
0751
06CE
05BD
05E6
074D
0742
036D
FD29
F87B
F7C4
F97A
FA89
F9F0
F913
F934
F9DC
F9FF
F98D
F931
F91D
F902
F8F3
F955
F9D2
F96A
F840
F881
FC3A
025D
0736
0850
06EE
0601
0683
070D
068A
05D1
060A
06BC
06AB
05F6
05E3
06AA
06FA
0643
05E8
06ED
0789
04D5
FEE2
F962
F7A0
F8E8
FA08
F980
F8AD
F8EF
F99A
F972
F8D9
F900
F9D3
FA22
F9AF
F97C
F9E9
F9D9
F8BE
F86F
FB68
0142
0670
080F
06EE
05F3
0667
072B
0718
0699
0685
06AC
0666
05EB
0607
06A0
06AB
05EB
059E
0696
0755
054F
0039
FAE5
F85C
F8B8
F99B
F951
F86B
F843
F8F7
F98C
F984
F957
F96B
F97B
F953
F960
F9E2
FA1D
F96C
F8ED
FADE
FFC2
0508
0781
06D4
0585
05B2
06D6
073C
0699
0623
0677
06DC
06BD
06A3
0705
073A
069F
0601
0683
0747
05B1
00BA
FAEE
F7EF
F86E
F9D6
F9E5
F914
F8F4
F998
F9E6
F99C
F987
F9DC
F9D1
F917
F8A6
F930
F9BF
F91F
F846
F9D3
FE97
03F9
06C3
06B2
0622
06B2
07A2
07A6
06E2
0669
0683
068C
0645
0634
067C
066E
05CE
05A0
06B3
07C8
0667
01E0
FC7C
F933
F8B7
F959
F978
F914
F8F5
F93B
F974
F997
F9F7
FA6B
FA4B
F997
F946
F9E5
FA79
F9BC
F865
F90E
FD3B
0320
0732
07CE
0688
05D1
0645
06D9
06E0
06C3
06D0
069E
0602
05B2
0634
06CD
067F
05C5
0614
074F
0706
0330
FD33
F8D2
F813
F95E
FA0A
F984
F914
F95D
F9A7
F973
F956
F9C3
FA0E
F988
F8E3
F951
FA63
FA52
F8E7
F8B2
FC29
0235
0703
0839
0725
0677
06F8
077D
0740
06E1
06FB
0707
0662
058E
0577
05EA
05ED
0583
05DB
072B
076B
0457
FE88
F966
F7A8
F8A1
F99F
F939
F85B
F84D
F8EC
F956
F95F
F98B
F9E7
F9EF
F9A0
F9A1
FA0D
F9FA
F910
F8F2
FBD3
016E
068B
0849
0732
0622
069A
0774
0742
067A
0667
06FA
0705
0642
05C8
0636
06AE
065F
0604
0698
06FF
04BC
FF73
FA2D
F816
F8EE
F9EE
F992
F8ED
F947
FA0A
F9F3
F93B
F923
F9CA
F9FD
F961
F926
F9E8
FA49
F91C
F811
FA4C
002D
061B
0862
0740
05EA
0641
071C
06D6
05E0
05B9
067D
06FB
06BF
068F
06CC
06B5
05ED
058E
0693
07A3
05F3
00C5
FAE5
F7D3
F82A
F9A0
FA30
F9E5
F9A4
F983
F923
F8DA
F950
FA2A
FA42
F96F
F905
F9E0
FACF
FA39
F8EC
F9DC
FE7A
045E
07A5
073E
05AB
0597
06E3
07AC
0728
064C
0612
064E
0679
0698
06BF
0680
05AB
0534
0622
077C
0699
0233
FC6D
F8C1
F85A
F966
F9D8
F995
F992
F9DE
F9BE
F934
F926
F9CB
FA26
F999
F911
F997
FA73
FA1D
F8EC
F97B
FD89
0357
073A
0793
062D
059C
0651
06FA
06CE
0652
0625
0629
062C
067A
072B
078B
06FA
062A
0658
073B
069B
02DC
FD5B
F953
F87A
F97B
FA0F
F99F
F93A
F985
F9E2
F9A6
F92F
F92C
F97D
F98A
F95F
F98C
F9F1
F9AE
F8C5
F907
FC43
01AF
0633
079B
06C6
0619
0689
071E
06EE
0676
068B
0703
0720
06DA
06C8
06F4
06C0
063B
0663
0758
073F
041C
FEAD
FA2C
F8E7
F9E1
FA7B
F9B9
F8CE
F8D8
F95A
F96B
F937
F95F
F9AB
F96A
F8DF
F90D
F9F4
FA3A
F947
F8E3
FB6B
0096
0543
06F3
0666
0607
06B4
0745
06DD
0638
065A
06FB
0732
06F6
06F6
072A
06CE
05FC
0604
074F
07D1
0508
FF65
FA59
F8AA
F993
FA55
F9BC
F8F3
F91A
F9A4
F991
F921
F934
F9A1
F977
F8C1
F8AE
F9A4
FA44
F97A
F8B9
FAC1
FFFB
0562
07C8
0736
062C
063A
06B5
069F
0656
06AA
0748
0734
0682
064D
06E3
0734
06A0
062F
06E7
0784
057D
0060
FB02
F880
F8E9
F9CF
F9A4
F928
F97E
FA34
FA2B
F97C
F940
F9B6
F9F3
F987
F940
F9BE
FA1B
F949
F858
F9E5
FEC9
0473
077A
0744
061C
0606
06C0
0710
06CC
06B2
06DC
06A8
0613
05FE
06B5
0730
06A4
05FB
0692
07AC
069F
021D
FC5F
F8F9
F8F7
FA2D
FA4F
F971
F8FC
F950
F991
F95D
F957
F9D7
FA2F
F9D0
F95B
F99C
FA05
F96A
F855
F93F
FD9A
0374
073B
0796
0669
060F
06B6
0712
06AE
065C
0697
06C5
066D
0619
0656
0698
062A
05B3
0676
07EB
076F
033C
FD13
F8CB
F83B
F9A6
FA59
F9C3
F92A
F955
F9B2
F9BA
F9C2
FA19
FA40
F9CA
F961
F9DE
FA98
FA07
F861
F85F
FC3C
028A
0747
0823
069F
05A3
0611
06A8
0688
064E
069E
06E6
0672
05C4
05D7
067F
06B3
065F
0699
0792
074E
03CE
FE0C
F988
F886
F9CA
FA9A
FA0E
F953
F957
F99B
F97B
F95A
F9C7
FA50
FA23
F98C
F996
FA34
FA13
F8E5
F8BE
FBDC
0178
061E
0773
068C
0605
06BB
0769
070F
0659
0647
06A0
0691
0624
060A
0651
065A
062B
06AA
07DE
07E4
04B9
FF04
F9FF
F836
F90E
FA17
F9FD
F964
F93B
F96E
F985
F991
F9DC
FA1A
F9DE
F984
F9D8
FA96
FA6A
F903
F869
FB0B
0095
05C3
07C3
0704
0612
0657
0707
070A
06A3
069C
06CD
067E
05D4
05B5
0649
069B
062A
05E8
06AA
0736
052C
0036
FB11
F8B2
F91B
F9FD
F9DD
F965
F99C
FA25
FA11
F98E
F994
FA2A
FA49
F9AA
F968
FA24
FAA3
F99A
F84F
F9D1
FF1A
0532
0839
0794
060A
05EF
06C5
06E5
0630
05D6
0642
069D
0663
062F
067D
06BB
065B
0620
0704
080C
069C
01B2
FBC4
F85E
F860
F99E
F9F2
F976
F95B
F9CE
FA08
F9E3
FA09
FA81
FA63
F96D
F8D9
F99C
FA96
F9FC
F866
F8F3
FD8C
03FA
0806
0818
0687
0620
06EB
0724
0643
058F
05F7
06C4
06F3
06AA
0698
0696
061A
05A9
065E
07A7
06F4
02AE
FCC4
F8F3
F8AC
F9E8
FA2F
F982
F96E
FA41
FAAB
F9F8
F933
F967
FA02
F9E8
F960
F98C
FA57
FA5E
F963
F981
FCD5
0267
06C1
07BA
068D
05CC
0644
06E1
06CD
0675
065D
0643
05DF
05A6
0619
06BB
06AF
0637
0683
0798
0763
03F2
FE37
F98E
F849
F97F
FA9A
FA59
F9A5
F9A9
FA31
FA47
F9CB
F997
FA23
FAAC
FA23
F8B2
F7FD
F9C1
FE20
0348
06DB
07D4
071F
066D
067D
06BC
066A
05CE
05C4
066C
06D5
065E
05D5
0687
081F
0851
0527
FF79
FA7A
F89A
F95D
FA63
FA2E
F953
F917
F9A4
FA0A
F9AC
F914
F92E
F9F4
FA61
F9B1
F89D
F90E
FC5D
01B5
0661
081E
0731
05EB
060E
070F
073C
063E
0594
0663
07AF
079C
062A
0570
06B2
081F
0699
017C
FBB1
F8A1
F8CA
F9EA
FA01
F94B
F923
F9DE
FA7D
FA32
F96C
F923
F996
F9FE
F997
F8BC
F8F8
FBB1
00A0
05A0
0846
0800
067B
05D0
066F
0717
06C4
05FC
05E4
068B
06E4
0663
05EF
068F
0799
06E8
0338
FDDB
F9A4
F83B
F8D9
F99E
F99B
F94D
F968
F9CE
F9E8
F99D
F981
F9FA
FA8A
FA4D
F938
F8A7
FA5C
FEB6
03F4
0774
07F7
069E
05A2
0614
0710
0738
0682
061B
069A
0726
06B5
05C3
05D0
0718
0791
04EC
FF73
FA32
F7F5
F8A7
F9F0
FA12
F972
F959
FA05
FA7E
FA1B
F975
F98A
FA4B
FA94
F9B5
F8AD
F981
FD2F
026D
0691
07EB
0723
0638
064F
06D1
06AA
05ED
05B3
0674
073C
06DD
05AC
0548
0667
0774
05EF
013F
FBAF
F858
F842
F9C7
FAA9
FA48
F9AC
F9C8
FA49
FA45
F9A1
F940
F9BD
FA73
FA42
F944
F93E
FBF1
00FB
05D6
081E
07BB
0699
0662
06E5
06EF
0625
0584
05EB
06D0
06EA
060B
0583
0659
0782
0696
0282
FD0C
F943
F888
F98B
FA1F
F996
F8F5
F93C
FA15
FA75
FA08
F987
F99D
F9FB
F9DD
F945
F969
FB95
FFBB
0430
06FF
0787
06CD
0649
067E
06D3
069C
060B
05DF
0649
06A7
066A
0607
0659
0727
06C0
03A9
FE98
FA35
F89C
F956
FA2A
F9BA
F8D2
F8F0
FA1B
FADD
FA46
F937
F934
FA45
FAD8
F9E6
F8B6
F9C9
FE0B
0386
072E
07C2
06A2
05EE
0652
06DB
06A5
060D
0610
06D5
076A
0709
063A
0631
0709
0721
04B1
FFED
FB34
F8D8
F8FA
F9CA
F9CF
F959
F990
FA89
FB0A
FA35
F8DC
F895
F9AC
FA9D
FA01
F897
F8E0
FC72
0216
06BC
0852
0770
0648
063F
06E1
0706
067A
061B
067E
070C
06D4
0602
05E1
070E
0820
06B7
0222
FC8A
F902
F89A
F9AD
FA15
F973
F903
F98D
FA48
FA15
F922
F8C0
F98A
FA79
FA2C
F8E7
F8B2
FB4A
0025
04D1
0737
0753
06B1
0694
06EE
0701
069A
064E
0694
070C
06FF
066D
0639
06F9
07CF
06E4
0347
FE2C
FA16
F89B
F927
F9EF
F9E2
F968
F95C
F9C4
F9EA
F980
F925
F983
FA39
FA2F
F921
F881
FA47
FEC7
0400
074D
07C6
06C0
061C
0665
06C9
0696
0635
066A
0714
0739
0672
05B6
063B
079B
07AF
04AD
FF51
FA76
F86C
F8F2
F9F4
F9F8
F962
F95A
FA11
FA9A
FA47
F993
F970
F9EF
FA20
F967
F8A2
F999
FD30
0243
0670
0818
079E
06AE
0672
06AB
0686
05F5
05C8
0667
0707
06A7
059F
057A
06D4
07F5
0645
0151
FBBF
F8BD
F8E0
FA07
FA1F
F94C
F90A
F9D5
FA8F
FA29
F932
F913
FA1B
FAF8
FA64
F8F9
F8EA
FBD3
00F7
05BB
07EC
0786
0650
05F5
068E
0713
06DA
0657
0654
06C8
06EE
067B
0631
06C4
076F
0643
0243
FCE5
F905
F836
F969
FA55
F9F1
F92C
F94C
FA2D
FA8F
F9DC
F8FD
F91B
F9F3
FA20
F925
F8A6
FAE0
FFF6
054F
0804
07AD
0663
0628
06E8
0738
068A
05D9
0629
0709
0733
065F
05C9
0690
07F8
07BD
0463
FEEC
FA1D
F809
F875
F989
F9D3
F970
F951
F9D3
FA4E
FA1A
F984
F96F
FA06
FA57
F993
F894
F982
FD90
034B
0795
0889
0723
05EA
0630
0713
0725
065D
05EC
0667
06F3
069C
05DF
0619
075F
07B6
0514
FFE5
FAFE
F8CB
F919
F9D8
F9AB
F90E
F91A
F9D1
FA3B
F9CF
F938
F965
FA3C
FAAB
F9FE
F901
F983
FCAC
01B0
0631
082B
07A0
0661
061E
06DC
0764
0706
066B
0678
06F8
06F5
064A
060D
06F0
07BB
062F
01A6
FC30
F8BD
F85B
F98B
FA40
F9E6
F95A
F95B
F9A3
F99A
F94E
F95B
F9E6
FA38
F992
F86F
F88B
FB5D
0070
056F
0815
0812
06FF
0689
06E0
0711
0695
060A
063F
06F4
0727
0685
060D
06BF
07EF
076F
03D4
FE4D
F9D5
F862
F930
F9F0
F973
F8A2
F8E1
FA13
FAC1
FA17
F902
F8F6
F9E7
FA4D
F953
F867
F9F7
FEA0
0422
0778
07B5
068A
0619
06BD
0745
06E3
0643
0678
0761
07BB
06DD
05CF
0618
0790
07EE
0512
FF8D
FA6A
F844
F8EB
FA13
FA11
F951
F923
F9C4
FA2A
F9A4
F8E4
F90B
FA02
FA74
F990
F870
F94E
FD2D
0292
06AE
07E5
070F
0642
069E
076F
077B
06A5
05FB
0638
06CB
06B5
060D
0604
0716
07D4
0612
0163
FBF6
F8AE
F878
F9C7
FA7F
FA0B
F965
F981
FA21
FA5E
F9EE
F97A
F9A1
FA0C
F9D7
F907
F927
FBEA
0113
061B
0863
07AA
0610
05A8
0671
06F5
0679
05D6
0610
06CD
06E1
061E
05C3
06B3
07D6
06DA
02CC
FD6A
F995
F89C
F95F
F9F6
F9BD
F97A
F9E2
FA85
FA7E
F9C2
F94D
F9D7
FAB3
FA8B
F937
F881
FA8A
FF73
04D8
07E5
07DD
0673
05C1
0647
06F5
06DD
064B
0621
068D
06DB
0689
061D
066C
072C
06BB
03B2
FEBB
FA56
F89C
F952
FA64
FA42
F959
F915
F9D4
FA80
FA28
F969
F98A
FA92
FB00
F9D9
F880
F9A2
FE2C
03E7
0782
07CE
0687
060B
06D9
079D
0746
0650
05F4
067B
06FF
06B2
05FE
05FD
06EA
0760
057A
00D9
FB74
F815
F7E3
F976
FA72
F9F4
F919
F92D
F9ED
FA11
F947
F8C1
F975
FA83
FA48
F8F1
F901
FC90
0284
074B
0879
0716
05F2
066C
0773
078C
06C6
0653
06B6
0726
06D0
061A
0623
071F
07A4
05E0
0178
FC2F
F896
F7EE
F939
FA53
FA10
F916
F8BF
F960
FA12
FA08
F99C
F9A8
FA26
FA27
F967
F94B
FBAB
0092
05B8
0886
086D
0714
0662
06B7
0723
06EB
0668
065B
06D4
071A
06AF
0618
063C
06EE
0684
0364
FE14
F948
F77A
F889
FA13
FA2B
F933
F8CF
F981
FA23
F9BC
F906
F959
FA90
FAFC
F9C3
F894
FA1D
FEED
0482
07B9
07D4
06AB
064D
0702
07AD
0783
06DE
0685
06AB
06DE
06BF
067D
0688
06CB
065B
041A
FFF4
FB74
F8B8
F890
F9B8
FA42
F99C
F8DE
F911
F9C7
F9D5
F91C
F8C5
F980
FA57
FA00
F904
F9AE
FD6D
02D6
06D0
07AF
06A5
0600
069C
076F
0754
0697
065C
0704
07A9
0755
066A
063D
073B
07D7
05E7
012C
FBFB
F914
F901
F9F6
FA28
F997
F950
F98F
F999
F92C
F90C
F9A0
F9F9
F937
F87A
FA38
FF2F
04E4
0805
07DF
0699
063D
06A2
06AE
065A
0676
06F6
06ED
064B
0650
0782
080B
0574
FFF6
FACE
F8C9
F95F
FA00
F97A
F8E9
F967
FA4B
FA5B
F9C0
F99B
FA01
F9C5
F8A9
F8A7
FBDF
0192
0665
07E2
06E0
05F3
063F
06CB
06A0
063F
0689
0728
071D
0689
06A0
0781
072D
03B8
FE18
F9A1
F87D
F987
FA2D
F998
F904
F966
FA07
F9E8
F970
F99D
FA23
F9C3
F8B1
F949
FD4E
0330
0747
07CA
0670
05E8
06AF
0754
0712
06BD
0701
0732
06A0
0621
06E2
07F6
06A3
01C0
FBC1
F861
F89F
FA1C
FA5A
F971
F8FE
F979
F9DD
F998
F96A
F9D7
F9FA
F8FE
F831
FA28
FF7A
0553
083A
07B3
0649
062D
06FD
0737
06AD
0670
06CD
06DB
0648
063C
076E
0829
05B6
FFF8
FA4D
F815
F912
FA46
F9E8
F903
F925
F9EF
FA08
F97E
F989
FA3E
FA19
F89D
F819
FB40
0160
068B
07F1
06C1
0601
06A4
0730
06AE
061F
0694
0742
06D2
05CF
0616
07AE
07D5
042E
FE16
F973
F86C
F985
FA26
F9BE
F97F
F9F5
FA3A
F9AF
F927
F993
FA46
F9DA
F8AE
F939
FD31
0303
072A
07D4
067F
05C0
0657
070F
06F9
0699
06B2
06F0
06A4
063D
06BA
079F
06A8
026F
FCB8
F906
F8D8
FA41
FAA0
F9B5
F928
F9AA
FA15
F98B
F8EE
F952
FA02
F98A
F887
F9B5
FE71
0459
07A4
0761
0618
0624
0702
06F9
0611
05E1
06D9
077D
06D8
0627
06E3
07EF
0656
012B
FB44
F842
F8A9
F9F6
FA1D
F993
F99F
FA2C
FA2E
F99C
F984
FA30
FA66
F95B
F89D
FAC3
0015
05A3
0838
079F
063E
05F9
0683
06B8
0684
0694
06D8
068F
05D7
05F0
072F
078A
048D
FEB0
F989
F806
F963
FA9D
FA3A
F96A
F98B
FA1B
F9EE
F951
F98B
FA7F
FA8F
F961
F953
FCCC
02B9
0734
07E0
0650
0591
0666
072F
06DD
065F
06B3
072D
06B2
05D5
0613
071B
0668
0252
FC9B
F8D1
F86E
F9B0
FA3C
F9C8
F97B
F9AE
F9A6
F92F
F933
FA1D
FAC5
FA01
F8E1
FA14
FEAB
0458
07B6
07D2
06B5
067F
0717
0734
06A3
066B
06EB
072F
068F
0600
06A9
0794
0624
0150
FB7F
F82E
F838
F96B
F9A5
F921
F935
F9ED
FA28
F9A0
F961
F9EF
FA38
F955
F8A7
FAC0
FFFA
0576
081E
07DA
06ED
06D9
0718
06DB
068C
06D9
0737
06A1
058E
05B4
0758
07FF
0508
FF1B
F9D9
F7FC
F8CB
F9B7
F993
F93A
F980
F9E2
F9AC
F955
F9C5
FA95
FA62
F91C
F8FC
FC2F
01F1
06E4
0882
077F
0666
0688
0713
06FA
0688
068C
06D7
06A0
0617
064D
0731
06BB
031F
FD7D
F929
F81E
F91A
F9A5
F92E
F8FD
F9A9
FA23
F9A7
F927
F9C1
FAAA
FA3C
F8EB
F994
FDFA
0403
07C6
07EF
06C5
06BE
078E
0780
067A
060B
06CB
076D
06E6
0638
06CB
07B5
063C
015F
FBA5
F878
F876
F963
F960
F8DC
F90F
F9D4
FA0D
F98F
F959
F9D0
F9EB
F8F4
F85F
FA99
FFD9
053E
07C0
075D
068B
06E8
07A8
0771
0691
0661
0704
0733
0671
0614
0721
07EB
0586
FFB8
FA06
F7F9
F937
FA78
F9D1
F89B
F8C8
F9F7
FA51
F984
F91D
F9D6
FA51
F976
F8EE
FB85
013D
069A
0869
073B
0615
0688
075E
071E
064A
063A
06E1
0708
0678
0666
072A
06E2
0385
FDEA
F96B
F846
F95E
FA1F
F9AE
F943
F9B8
FA45
FA01
F97D
F9BF
FA52
F9D8
F8A4
F947
FD8F
03AB
07B2
07E8
065D
05EE
06DC
075D
06AD
0605
0660
06E5
0682
05EE
0695
07C5
06AE
01E7
FBD6
F85D
F899
FA16
FA4D
F96E
F920
F9B3
F9F6
F97B
F951
FA16
FAA2
F9C4
F8B1
FA33
FF1B
04BF
07BB
0792
068C
0682
0706
06F3
067C
0698
071C
06E2
05D5
0586
06CF
07CE
05A7
0035
FAC8
F896
F953
FA39
F9BD
F8F2
F932
F9FC
FA09
F982
F9AA
FA8B
FA93
F92D
F890
FB72
0150
0663
07CA
0693
05D7
06BF
07B4
0743
062E
05F8
068D
06A8
0623
0643
0756
0749
03F0
FE2A
F97B
F847
F976
FA57
F9EE
F95F
F998
F9FD
F9C4
F971
F9E4
FA94
FA1A
F8C1
F91F
FD2C
0350
07A7
082A
0699
05D7
0685
0721
06C7
0658
06AB
070F
0690
05E5
0681
07D3
0704
0268
FC30
F86B
F887
FA27
FA75
F966
F8DC
F986
FA24
F9CC
F949
F98A
F9E6
F946
F88C
FA31
FF09
0496
0787
0755
065A
0692
077E
07A4
06F1
0686
06BD
06C3
0647
064B
0761
07F8
05AD
0067
FB0A
F889
F8E6
F9D0
F9B4
F921
F927
F994
F993
F94A
F998
FA5B
FA3B
F8DE
F859
FB36
011A
0687
0878
0779
0660
06AF
075D
0724
067E
0690
0724
070A
0648
0653
078A
07B9
0472
FE7E
F988
F80D
F8E3
F96A
F8FF
F8FD
F9F0
FA91
F9E1
F8E5
F911
F9E1
F991
F841
F8A8
FCC6
02E4
0732
0800
0712
06C4
073E
073C
0683
0635
06D7
0766
0704
0689
073C
085C
0758
02E1
FCFC
F919
F883
F981
F9D5
F936
F8D5
F939
F9A2
F97D
F952
F9A7
F9C9
F8DC
F7DE
F94F
FE2D
0428
07BA
07DB
06AC
067B
0736
0766
06C7
067C
0701
0756
06D2
0681
0774
0863
0696
0163
FB97
F89A
F8D4
F9DC
F9CA
F91C
F91A
F9A4
F9B2
F933
F926
F9BB
F9C6
F8AE
F820
FA88
FFED
0550
07AF
0714
0606
0648
0735
0764
06DD
06B3
0717
0727
06A7
06A8
07A3
07D4
04EA
FF47
FA5B
F8F6
FA31
FAF0
F9F4
F8D2
F907
F9C2
F992
F8D8
F905
F9F1
F9E7
F89F
F891
FC0F
01DE
0637
0718
0626
05E5
0697
06E9
069C
06C2
0794
07CF
06C4
05D0
069B
0855
07FD
03D0
FDAE
F954
F886
F9B7
FA69
F9E6
F93E
F94C
F9AF
F9B6
F982
F9A1
F9DB
F955
F85A
F905
FD0A
0301
0746
07E8
069C
0637
0732
07CB
0714
0633
0659
06DC
0697
0623
06EF
0834
06F8
01F5
FBF6
F8CD
F8F4
F9C1
F95A
F8AB
F917
FA18
FA3C
F994
F97C
FA2B
FA1A
F8A6
F7E2
FA6E
FFF5
0533
0780
073E
0698
06C4
0740
0737
06C8
06AA
06E8
06CE
063D
0634
0743
07E5
05A4
0038
FA9C
F82D
F90C
FA4C
F9CB
F898
F8C6
FA05
FA3C
F918
F89E
F9B1
FA5B
F923
F845
FB3E
01AE
071A
083D
06AE
060E
071F
07B2
06C6
060B
06BC
077B
06DB
0617
070C
089B
077E
02A5
FCCF
F95B
F8DE
F98C
F9E8
F9D6
F99F
F948
F91C
F997
FA3F
F9D3
F873
F86A
FB97
00E1
0561
0779
07B9
0741
06A3
0636
064C
06B8
06D1
0670
0671
075B
07EB
0605
0163
FC52
F947
F896
F917
F9D7
FA5E
FA32
F95F
F8E6
F97E
FA51
F9FD
F8DC
F92F
FC97
01EF
0657
0811
07B4
06C5
0626
060B
066A
06C9
0689
05FF
065B
07AE
07F5
052D
FFFB
FB27
F8C3
F89E
F954
F9ED
FA2C
FA15
F9DE
FA00
FA85
FA7E
F934
F7F6
F963
FE33
03D6
0728
07A3
06FC
0695
067C
066C
066E
066A
061E
05D8
065D
0785
0780
0486
FF3A
FA77
F873
F8C9
F9B7
FA2F
FA18
F99D
F92B
F96C
FA4D
FA97
F997
F8B5
FA50
FEE9
043C
077B
07E7
06E8
0618
05FD
065D
06D6
06E7
065C
05FD
06C9
0800
0726
02F2
FD5D
F9A1
F8D1
F96C
F9CF
F9C7
F9CA
F9DA
F9C4
F9BF
F9F2
F9D0
F904
F8DA
FB60
008A
057F
0795
0715
062E
0619
0677
06B6
06C4
06A5
0662
0672
0730
07A9
05E9
013D
FBBE
F898
F8B2
FA05
FA68
F9D4
F96E
F98E
F9CD
F9F8
F9FD
F980
F8B9
F943
FCB2
0247
0704
088C
0764
05FE
05F3
06C8
0740
06EF
0646
05E8
0653
0755
077B
04ED
FFCA
FAC0
F87A
F8E7
F9E1
F9F1
F972
F943
F97B
F9AE
F9BD
F9B4
F973
F93E
FA5F
FE0D
0356
0757
0832
0703
0629
067A
070A
06FE
067D
061A
0636
06E7
07AC
072B
0422
FF06
FA45
F833
F8C2
F9E1
FA05
F985
F958
F99B
F9DC
F9F4
F9CD
F937
F8CF
FA4A
FEA5
0444
07FE
084A
06AE
05BA
0640
0710
070A
0677
063F
06B1
076B
07B3
0674
02D7
FDA8
F971
F831
F94D
FA71
FA39
F950
F900
F992
FA3D
FA36
F96C
F890
F8DD
FB7F
0063
057D
082A
07C0
0634
05C7
06A4
0765
0734
068B
0642
069F
0742
074C
05A7
01DA
FCF9
F945
F840
F93A
FA22
F9DE
F926
F914
F99F
F9F5
F9AB
F90D
F8C7
F9CC
FCF4
01DA
066A
0868
07A3
061D
05D3
06C8
0785
0725
064D
061E
06DB
07BE
0788
0521
0075
FB30
F7FB
F80D
F9DB
FAC2
F9DA
F88E
F888
F9B2
FA91
FA20
F8E5
F86C
FA0C
FE04
0328
0741
0888
074F
05CC
05D6
0718
07E0
0754
0643
05F8
06C1
07A2
0715
0426
FF4F
FA7F
F7E9
F838
F9E4
FAAF
F9EE
F8EC
F8FF
F9DA
FA28
F95A
F858
F89C
FB0C
FF68
043E
078D
0829
06CB
058A
05D1
0708
0783
06B3
05D7
064F
07CA
0873
06C1
02B9
FDC8
F9D9
F83D
F8D8
FA35
FAB8
FA0A
F930
F937
F9F2
FA3C
F96F
F863
F8C1
FB8E
003E
04FC
07D3
080C
06BB
05CB
062E
071D
074A
0683
05DD
064D
0771
07CA
0602
0205
FD20
F94B
F7F0
F8D6
FA33
FA4B
F92B
F874
F930
FA77
FA9A
F95A
F85E
F97D
FD07
01AE
05A9
07C7
07ED
0705
0666
06BB
0760
0738
063F
05C5
06AD
0802
07B6
04C1
000E
FB9A
F8F4
F86F
F938
F9F9
F9D6
F91C
F8DB
F99A
FA7F
FA40
F8F1
F859
FA32
FE65
0336
06BB
0806
0764
0621
05B1
067E
077D
0763
064A
05B0
068F
07D9
0755
03F8
FEFC
FAA5
F86B
F863
F999
FAA1
FA74
F967
F8E2
F9A1
FA96
FA36
F8BC
F854
FAD3
FFA5
0465
0726
07BF
0725
0659
060A
066C
06F2
06C7
060D
05FC
0729
082A
06CB
029C
FD8B
FA06
F8E5
F945
F9D9
F9FA
F9AD
F958
F977
FA0E
FA59
F98D
F84E
F89B
FBBC
00A6
04F7
0725
075E
06B5
0628
063C
06D0
0733
06D6
0625
0639
0752
07F1
0621
01BA
FCD3
F9AE
F8D2
F94E
FA08
FA4D
F9D3
F907
F8DF
F9AC
FA6A
F9F2
F8DA
F946
FC94
019E
05C3
0770
0736
068E
0659
06A6
071E
0738
069B
05DC
0616
073B
0772
04EF
0033
FBB0
F956
F90C
F980
F9C3
F9B4
F986
F96F
F9AD
FA32
FA45
F961
F88E
F9F0
FE3E
0379
06D5
077E
06CC
064B
0669
06CC
070B
06DF
0654
05FC
0683
0788
0740
0419
FED1
FA36
F86C
F907
FA12
FA4A
F9CC
F946
F941
F9DB
FA7B
FA2C
F8EB
F85D
FA74
FF39
0460
0762
07B8
06D7
064B
066B
06C3
06E4
069B
060D
05F1
06E0
07F6
0706
02FE
FD8E
F9A6
F890
F939
F9F0
FA0C
F9D1
F99F
F9A3
F9F3
FA43
F9E5
F8D1
F89F
FB4D
009C
05A8
07CF
0745
062C
05E2
0637
0690
06B9
06AB
0678
0687
072D
07A1
0618
01BA
FC47
F8CD
F88E
F9ED
FAAD
FA53
F9CA
F9A8
F9C4
F9DD
F9C1
F93A
F8AD
F97B
FCD0
01EB
0645
07E3
0722
05F4
05AC
0612
066A
067B
0667
0650
0685
072E
0760
055D
00B7
FB8A
F8A7
F8BF
FA13
FAB2
FA47
F9AF
F99C
FA00
FA68
FA5B
F9A1
F8DD
F9AF
FD55
02BC
06E8
07DD
069B
0592
05DC
06B3
06FE
068B
05DC
059A
062B
0727
071D
0495
FFC8
FB06
F8B7
F90A
FA13
FA39
F9B5
F988
F9E5
FA47
FA52
F9E5
F915
F8B9
FA65
FEC2
0418
0779
07AB
0640
0596
0639
06E8
06A8
05F8
05D5
067C
0772
07F3
06E7
035B
FE02
F97B
F812
F960
FAE0
FAD3
F9C4
F940
F9C0
FA63
FA3B
F951
F881
F8EA
FB71
0001
04F2
07E0
07DD
0661
058F
05FF
06B4
06C7
065E
0629
068E
074E
0786
0607
0241
FD39
F93D
F805
F90F
FA45
FA42
F98B
F94F
F9C8
FA33
F9FB
F948
F8D4
F9AD
FCAE
0175
0607
0832
079D
0616
05A9
0694
0774
0730
0637
05C4
0664
0760
0754
0510
0097
FB92
F867
F82B
F99D
FA86
F9FE
F902
F8E7
F9C8
FA91
FA51
F944
F8BD
FA26
FDF2
02FB
070A
086A
076E
0614
05F3
06CA
0742
06B9
05E0
05C2
069B
0785
0704
0418
FF40
FA7E
F7FF
F848
F9D1
FA96
FA0D
F94D
F969
FA25
FA71
F9D4
F8F3
F907
FB0C
FF0F
03D6
075A
083F
0710
05BC
05B8
06B2
0747
06C3
05EA
05ED
06E6
078D
0658
02D2
FE11
FA0E
F851
F8CD
FA09
FA84
F9FB
F956
F96F
FA1C
FA70
F9D3
F8E2
F926
FBC8
005C
04ED
0775
0781
0671
05FE
0694
0735
06EB
05FF
0594
0649
0774
07A0
05A7
019C
FCE6
F979
F87F
F975
FA9D
FA8F
F96F
F89C
F91C
FA6C
FB0A
FA2A
F8D8
F92B
FC54
0161
05DF
07DC
075D
060A
058B
0639
0732
0774
06CD
05FE
05F8
06C0
070A
0530
00ED
FC04
F8E0
F878
F99F
FA70
FA29
F97F
F95B
F9C1
F9F9
F98D
F8D8
F8DB
FA9A
FE4D
02DE
066D
07B4
0712
0611
05EC
069C
0739
0711
065B
05EE
0661
073C
0702
0449
FF4C
FA4F
F7E9
F8A2
FA7C
FB22
FA26
F8EA
F8BC
F98A
FA40
FA08
F929
F8F4
FAE3
FF40
046C
07C9
080B
0682
05A5
064F
071D
06B6
05CB
05FC
074F
07BF
057C
00F4
FC5A
F990
F8D2
F928
F98A
F986
F956
F97C
FA10
FA65
F9D8
F922
FA39
FE2A
0374
0736
0806
0713
066E
06BD
0710
06A3
0605
0646
075E
07D5
060A
01C7
FCB1
F929
F86A
F97E
FA43
F9AF
F8BF
F8E9
FA0D
FA8C
F988
F865
F997
FDE7
0367
0729
07E7
06CA
05E5
0630
06FE
0726
0689
063D
0710
0800
06D6
0292
FCFA
F92A
F89D
F9F9
FACD
FA2C
F929
F917
F9D0
FA13
F93F
F85F
F959
FD1F
027C
06C7
0811
06DD
057D
0599
06A5
0706
0664
0616
071F
0856
0745
02F1
FD44
F95A
F8A1
F9DC
FAC7
FA59
F961
F936
FA03
FA8A
F9B4
F849
F8A5
FC55
0228
06EF
0868
0730
05BD
05B0
067B
06AD
0604
05B2
06A7
0804
0796
0405
FE6E
F9BB
F81A
F919
FA60
FA45
F956
F92B
FA23
FADE
FA19
F898
F8B2
FBF1
0156
0622
0833
0798
061F
058B
0620
06CA
06A0
0614
064F
0750
0745
0454
FEFB
FA0E
F81D
F909
FA7D
FA9E
F9C1
F963
FA06
FAA1
FA19
F8E2
F8E3
FBB6
00E2
05E9
0849
07AB
0603
056E
062C
06D7
067C
05DA
063B
0762
0747
0442
FF15
FA7B
F89E
F942
FA65
FA6B
F98B
F926
F9E7
FAD1
FA6F
F8E9
F867
FB08
0077
05DE
0866
07BF
0606
0569
0625
06EB
06C0
0618
0618
06F8
0756
0559
00B1
FB66
F849
F85E
F9F4
FA97
F9AE
F8C4
F944
FA88
FAB2
F94B
F854
FA46
FF47
04BA
07B2
0787
060D
0578
064B
0743
0729
0651
0617
06F7
0789
05CA
0161
FC50
F934
F8EE
FA13
FAA4
FA07
F937
F945
F9FF
FA3A
F965
F89D
F9ED
FE2D
03A9
075C
07C0
062E
0540
0607
0741
0751
065A
05F2
06D9
07AC
0641
0213
FD00
F998
F8E4
F9CB
FA6D
F9F5
F925
F921
F9EA
FA49
F977
F87F
F98D
FDA2
032B
0730
0807
06B5
0599
05FA
0718
077D
06D4
0630
068F
0754
068C
02F8
FDB4
F985
F84C
F94F
FA41
F9CC
F8BE
F8A5
F9AF
FA6E
F9CB
F8B5
F96B
FD1C
0274
06AD
07FB
06FF
05E2
0624
074F
07DD
0732
064A
0660
071B
0699
036D
FE69
FA15
F85D
F8EC
F9E0
F9DA
F922
F8DD
F979
FA23
F9E2
F90D
F965
FC64
0176
0619
0811
076D
0639
0635
0729
0793
06C0
05B8
05DA
06E5
06DE
0412
FF11
FA6A
F85F
F8E5
F9FE
F9F6
F90E
F8CD
F9D7
FAFB
FAB2
F94C
F90B
FBDF
0124
0601
080C
0761
0618
05F1
06C4
0734
068B
0596
059A
0698
06DC
048E
FFCB
FAE8
F867
F8AD
F9EC
FA3C
F98C
F93E
FA15
FB1F
FAE4
F97D
F8EE
FB3A
0036
0566
081F
07C9
0628
0572
0630
0714
06D0
05B8
054E
0635
06F3
0549
00B9
FB75
F86B
F883
FA08
FAB8
FA17
F975
F9F0
FAEE
FAEE
F9A3
F8D0
FAA7
FF5C
049B
0797
078E
0629
0585
061F
06CC
0683
05AC
0586
0662
06E4
053D
0124
FC66
F965
F8FB
F9E1
FA3E
F99F
F928
F9D9
FB0A
FB1F
F9B8
F8B2
FA70
FF36
0486
0767
072B
05BF
0567
067A
0777
070D
05B3
0518
0603
0718
0600
01DD
FC7D
F8DD
F86B
F9D8
FABA
FA1B
F929
F963
FA93
FB0F
F9F9
F8B8
F9D1
FE3A
0401
07E3
0840
066E
0520
05A1
06E4
0733
0654
05AE
0648
072A
062B
024C
FD04
F901
F7C9
F8B3
F9F3
FA5F
FA2C
FA21
FA64
FA49
F961
F897
F9CA
FDDC
0355
074B
080A
06A8
05AE
0652
0771
075E
0621
055E
061D
073D
0673
02AB
FD55
F938
F810
F931
FA73
FA5C
F95D
F8F4
F9AE
FA70
F9FC
F8F6
F9B2
FD9F
0341
075A
080A
0680
0569
0614
0770
07BC
06AD
05A7
05E3
06C9
0649
02FA
FDCE
F983
F829
F93F
FA68
FA0C
F8E7
F8BF
F9F2
FAED
FA41
F8C5
F913
FCC0
026A
06DB
0804
06BF
059A
0627
079F
0812
06C3
0519
04FD
066E
0717
049E
FF4F
FA1C
F7DC
F8B0
FA45
FA7F
F980
F8EB
F996
FA85
FA4C
F921
F90E
FBE4
011A
05F4
07F9
072D
05C3
05B1
06CB
076D
06BA
05B4
05E1
0724
0770
04DC
FFCD
FAD1
F855
F89A
F9EF
FA95
FA43
F9DA
F9EC
FA03
F963
F868
F8AC
FB93
009B
0562
0797
0703
0592
0547
0650
073C
06F1
0607
05F5
0709
0796
0588
00B5
FB66
F862
F875
FA08
FAF3
FA8B
F9C7
F9A3
F9DD
F98C
F8B9
F8D9
FB61
0001
048C
06E0
06CB
05EF
05E9
06C2
0748
06B7
05BB
05A5
06B9
077D
05F7
01B1
FC7A
F8F6
F858
F984
FA6D
FA28
F97D
F980
FA0D
FA0E
F92B
F8BC
FA97
FEF2
03CA
06AC
06F5
0629
0621
0713
07A3
06D3
0568
0526
0694
07F6
06C3
024B
FC9D
F8C4
F815
F955
FA60
FA41
F9A0
F971
F9B0
F99F
F902
F8D5
FA87
FE72
032E
0690
077F
06C6
0621
0670
0711
06F6
062A
05E1
06D5
07ED
06F5
02DA
FD1D
F8C6
F7C7
F95C
FB00
FAF0
F9A9
F8DE
F948
F9E3
F980
F8B7
F9A7
FD8B
02EB
06BE
0766
062B
058A
066D
077A
0723
05BC
0521
065B
0808
077D
0376
FD98
F917
F7F2
F960
FAF1
FAFD
F9ED
F937
F97E
F9F9
F9BB
F931
F9EE
FD00
019E
05A6
076C
071B
0642
0625
0697
0692
05CA
0541
0607
077D
0764
040A
FE69
F998
F7FF
F935
FAC7
FAE7
F9ED
F95C
F9D3
FA72
FA2B
F95B
F9B5
FC89
0132
056D
0754
06FE
0629
063D
06EA
06D8
059F
0492
053A
072A
07D8
0505
FF42
F9CC
F7A9
F8EF
FAF6
FB35
F9BB
F8A4
F95F
FAF6
FB58
FA14
F93A
FB31
FFF4
04E8
0773
0768
06A0
0697
06F7
0694
0556
0497
0585
0765
07DD
0520
FFD2
FAB0
F83A
F8A9
FA19
FA98
F9ED
F956
F9B2
FA6C
FA53
F95A
F912
FB2D
FFA5
0474
074E
0794
069F
061D
0667
068F
05F9
0570
0639
081D
08D5
0613
0024
FA3D
F7B7
F900
FB6D
FC0C
FA6A
F886
F849
F96D
FA16
F94D
F873
F9FB
FEA2
0447
07BB
07B6
05E0
04DB
0598
06D2
0711
068C
06AB
07DB
087F
066C
015F
FBBD
F897
F8E9
FADE
FBBD
FA8B
F8AD
F814
F906
FA01
F9BA
F8EE
F9C5
FD6D
0293
0686
07B5
06E6
0606
061A
0695
068E
0628
0665
07A0
087D
06EE
0266
FCD8
F93B
F8D2
FA24
FAAD
F98F
F835
F85A
F9DA
FADC
FA1D
F8A1
F8E1
FC48
01A8
063F
081D
079A
068B
064C
06B7
06E3
068F
067F
0740
07F9
06D1
02E0
FD86
F980
F879
F999
FA8C
F9EF
F88F
F830
F948
FA5D
F9E1
F86F
F89E
FC41
0223
06EB
085F
0757
0649
0658
06A1
0642
0605
071F
08C0
081B
0382
FCE1
F842
F7BE
F99A
FAA1
F9C4
F8A1
F8CA
F9A4
F9A0
F8EC
F9C1
FD9C
02F7
06A1
0732
065D
0688
07C3
0825
06D8
0590
063A
07E7
074D
02A6
FC35
F81D
F804
F9C6
FA74
F9AA
F91A
F98D
F9B4
F873
F74C
F93C
FF04
0595
08DB
07E8
059D
052C
06B9
07F5
0783
0694
06D0
0789
0629
0182
FBC3
F856
F83C
F957
F966
F8AA
F8DF
FA3A
FAD3
F967
F7C0
F931
FEA5
051E
08A7
084D
068B
05FD
06B4
071C
06B4
06A6
0792
07D2
050E
FF68
FA1A
F848
F9A4
FB09
FA44
F865
F7DA
F90A
F9FB
F962
F8DD
FB2B
007E
05BE
07DE
0716
0617
0680
0746
06DB
05CC
0615
07FA
08C8
05A0
FF16
F91E
F725
F8C0
FABE
FAE8
F9E4
F966
F98E
F920
F809
F867
FC2D
023D
06F0
07D5
0633
053F
0647
07A1
0761
0613
05D4
0717
077F
0492
FEEA
F9DC
F801
F8CB
F9D9
F9F4
F9DD
FA5E
FAAA
F985
F7AC
F7E9
FC1A
02A0
0787
086F
06A7
0543
059B
0679
067D
062C
06D3
07F7
072A
02F2
FD22
F947
F8EF
FA36
FA5C
F90C
F84A
F95C
FAEC
FAD3
F940
F902
FC57
0213
06AF
07EF
06DA
05EF
0624
066F
05FD
05B9
06CA
082F
0718
0236
FBE9
F83A
F8B1
FAF5
FBBA
FA66
F902
F91C
F9D8
F9AD
F918
FA68
FEB0
03F1
0703
06F8
05D4
05D4
06D9
071A
05FE
0518
05E8
0757
067B
0203
FC1C
F85F
F822
F98C
FA36
F9DC
F9D4
FA7E
FA8B
F935
F837
FA57
FFE5
05AD
0816
06DE
050D
054A
070F
07FB
0729
0622
0658
06C0
04EA
003F
FB37
F8C6
F92A
FA0F
F9AD
F8CF
F931
FA99
FAE4
F929
F7B4
F9DB
FFE6
063A
08FD
07F6
0621
05DA
068E
0681
05BE
05F9
07A0
085C
057B
FF6D
F9D7
F7E5
F91D
FA6C
F9E5
F89B
F894
F9DF
FA9F
F9E1
F94F
FB5E
0025
04F1
0733
0724
06E3
0772
07AC
067A
04F8
0543
0749
0808
04C1
FE70
F924
F7BF
F93F
FA81
FA10
F92C
F947
F9C8
F934
F7F3
F89D
FCE4
0302
0727
0779
05DB
0561
06B1
07CD
0731
05FD
0645
07CF
07C6
040D
FE11
F97C
F853
F93A
F9B3
F938
F92D
FA39
FAEB
F9BA
F7AE
F7F4
FC5D
02FA
07C1
0882
06B4
0555
05AB
069F
06EA
06CF
073B
07B7
065C
0230
FCEB
F994
F953
FA5E
FA59
F91E
F87C
F96A
FA8F
FA2E
F8DF
F95E
FD4D
02F4
06E8
0798
068C
060D
067F
06A0
05F2
05AB
06D3
0815
06AB
01A2
FB8D
F82D
F8A2
FA86
FAF2
F9A1
F890
F8F3
F9B8
F979
F8FB
FA9C
FF28
0445
06DC
0680
05A4
0655
07D2
07F6
0671
0559
063C
079C
0652
0162
FB7F
F844
F885
F9FC
FA59
F9AA
F960
F9C2
F990
F84B
F7CF
FA8F
005F
05F3
0813
06DC
0537
0561
06C6
0781
0719
06CE
074F
0735
0496
FFAC
FB17
F934
F9BD
FA86
FA2B
F95E
F968
FA1B
FA14
F8F8
F897
FB25
0070
059B
07E1
0740
0602
05E6
0684
06A4
065A
06C5
07D7
077F
03E9
FE2A
F9B4
F8CE
FA40
FB09
F9E8
F865
F851
F94F
F99D
F8F1
F94A
FC82
01AA
05C1
06EF
0653
0632
071A
0794
06A5
0588
060E
07C1
07BD
03E1
FD9F
F8D5
F7D8
F960
FA7E
FA04
F92F
F93F
F995
F8F5
F7F8
F90F
FD8E
0382
0747
0755
05B2
055F
06E0
081B
076C
05E1
05A4
06C7
06B9
035A
FDDB
F9B0
F8C4
F9A6
F9C9
F8C6
F868
F9AE
FB0D
FA89
F8DA
F92B
FD60
037C
0782
07BB
0623
05A4
06B8
0799
0726
0661
069E
0723
05AC
015E
FC4A
F968
F966
FA39
F9DD
F8AB
F86F
F9A6
FAAE
FA17
F8FD
FA19
FE82
0409
0768
07A2
068C
0633
068E
065D
058C
058E
070E
0836
0645
00DF
FAF7
F7FC
F877
FA04
FA5F
F9AE
F971
FA00
FA1A
F917
F88F
FADA
000C
0548
0795
06EF
05E1
0647
074E
0717
05A4
04F9
0637
0781
05C4
006C
FA81
F794
F829
F9C0
FA1F
F996
F9AD
FA79
FA6D
F8F4
F821
FAB2
0094
0653
0888
0750
05BA
05FA
073A
076E
066A
05F8
06E6
074D
04A7
FF45
FA6C
F8CA
F99D
FA1E
F921
F833
F8F5
FA88
FAB1
F930
F8AB
FBAF
016D
0658
07ED
070A
0642
06A5
0714
068E
05F0
06A8
0821
07B0
0394
FD73
F914
F883
FA28
FAF9
F9F4
F8B8
F8E0
F9C2
F999
F86C
F8A1
FC36
01FE
0688
07B3
06A6
05F3
0676
06DC
0620
0553
061E
07F4
07F3
0411
FDD7
F919
F810
F963
FA49
F9D4
F954
F9C6
FA32
F941
F7DB
F8C5
FD56
0355
0705
0712
05A7
0581
06CA
0792
06D7
05F2
0682
07BB
06F0
02CC
FD3B
F983
F8E0
F9AB
F9CE
F933
F92B
FA05
FA51
F906
F79F
F8FF
FE0E
042C
07AC
0785
05FA
059C
0683
0704
0686
065B
0783
0882
06A7
0174
FBC2
F8F6
F972
FA9D
FA3A
F8DD
F882
F989
FA31
F945
F84D
FA0F
FF16
0495
074B
06E1
05D3
062C
074C
076B
0670
0628
0773
085E
060D
005E
FAA0
F842
F947
FAC3
FA80
F938
F8DF
F9AC
F9FA
F900
F88F
FB1E
007D
0584
075D
067B
05A4
066B
079A
075B
060B
05BB
0711
07C8
0527
FF81
FA3F
F844
F8FF
F9B6
F912
F857
F8FF
FA41
FA18
F86D
F7F4
FB33
013F
0658
07D1
06A7
05D1
06A3
07BB
0773
064C
0616
070D
06FE
03CB
FE4B
F9BE
F85F
F933
F9A6
F8C8
F80E
F8D4
FA3B
FA4E
F901
F8DC
FC23
01E0
0698
07F6
0704
0663
070E
07B7
072C
0642
0689
07A5
0714
0322
FD59
F93D
F8A2
F9F5
FA79
F97D
F89D
F91B
FA0A
F9CD
F8D0
F994
FDAA
0360
073F
07B3
0673
0611
06EE
0760
0683
05A9
0667
07D3
06FD
0268
FC3D
F84B
F80E
F987
FA08
F94C
F90B
F9FB
FAA1
F994
F820
F951
FE4B
046B
07D8
078E
0609
05F5
072A
0799
0687
0599
064C
076E
0623
0172
FBCF
F8A2
F8B0
F9CA
F9C2
F8D6
F8B0
F9AB
FA3F
F95A
F869
FA1C
FF1D
04D0
07D7
077E
060F
05E0
06D9
074F
06B4
065C
073A
07DC
05B2
005B
FABF
F832
F8F7
FA57
FA1B
F8EE
F8D0
F9F2
FA6E
F939
F83B
FA61
FFE1
057C
07E6
0730
0614
0669
074B
0717
0611
05FF
074A
07C5
0502
FF72
FA49
F83A
F8E0
F9D3
F9A5
F915
F957
FA20
FA1E
F928
F911
FBC2
00D4
0594
07AB
074C
0680
06A0
0712
06B2
05C7
05BC
06D6
071D
044D
FECC
F9C6
F7F8
F8E8
F9E6
F979
F8C7
F957
FA81
FA55
F8D0
F8B5
FC60
0277
0708
07D5
0678
05D6
0687
06E8
062B
059F
0651
06B9
0441
FEE2
F9C5
F7D5
F8A3
F994
F960
F90E
F98F
FA06
F976
F910
FB41
0055
0575
07B6
073D
0674
06A5
06DE
0641
05C8
0695
0767
0576
002F
FA92
F80E
F8B8
F9DA
F9B7
F93D
F9B0
FA4A
F9A0
F89D
FA25
FF48
0537
0826
0789
0628
0637
0701
06F2
0665
06D1
07B3
065D
017C
FB8A
F853
F8AF
FA00
F9F8
F931
F956
FA20
F9E5
F8D0
F98E
FDE1
03C1
0758
0762
062C
061D
06E2
06DE
0635
067A
0795
06EC
02AD
FCCA
F924
F908
FA1B
F9E1
F8DB
F8EE
F9F6
F9EF
F88C
F89F
FCA7
02FA
073D
076C
05E4
05C7
0706
075D
064E
05E3
071B
078C
043D
FE05
F924
F857
F9EC
FA96
F9B9
F944
FA07
FA59
F931
F8AF
FBC6
01EB
0705
0820
069D
05CA
0685
0700
064E
05FD
0737
0803
0547
FF2B
F9A2
F7F4
F92F
FA21
F9A3
F948
FA01
FA5D
F91E
F81D
FA91
0098
065D
085E
0743
0642
06BB
072A
066A
05D6
06EA
0818
0617
005D
FA7D
F828
F911
FA17
F9AA
F92E
F9E7
FA91
F985
F815
F99E
FF08
04FF
07AE
070D
0622
0699
071C
0647
0550
0619
07A6
0696
0196
FB9F
F89C
F8F6
F9D7
F962
F8B8
F95A
FA5B
F9DE
F88C
F97E
FE25
03E4
06F1
06B5
05DD
0655
0717
0688
0574
05D9
0756
06D3
0270
FC6A
F8C1
F8A4
F9AD
F994
F8E7
F93B
FA24
F9CF
F85D
F8AF
FCCE
02D6
06D1
0743
0657
0669
0715
06B4
0595
05BA
0753
077F
03B8
FD84
F913
F873
F99D
F9BD
F8D6
F8D9
FA0D
FA76
F92B
F88E
FB93
019E
06B6
080C
06DC
0622
06A8
06E6
0625
05D7
06FB
07B8
0538
FF94
FA4E
F86A
F939
F9F4
F982
F927
F9C0
FA21
F939
F890
FAE0
0055
05AC
07CC
071B
064C
06A0
06EF
064E
05E2
06E3
07E1
05E6
0071
FABD
F83E
F8DD
F9CF
F984
F91D
F9C0
FA5C
F973
F832
F9BC
FF0C
050D
07EB
0751
0621
064E
06DD
065C
05A2
066C
07EC
06EA
01E7
FBAB
F85D
F8C4
FA03
F9BE
F8D5
F91D
FA14
F9B7
F838
F8B9
FD51
03C5
07B4
079D
060D
05CA
068B
0689
05E0
0655
07E6
07AC
036F
FD12
F8D6
F879
F9BA
F9E4
F92C
F94F
FA2D
F9DF
F840
F843
FC63
02E2
0752
07AE
0644
061E
0720
072A
05FF
05C7
075E
0814
04C6
FE55
F92D
F831
F9BF
FA75
F994
F906
F9B2
FA06
F8E2
F83F
FB19
0129
0688
0811
06C5
05D5
066C
0702
068C
0641
073B
07D3
053B
FF83
FA40
F882
F977
FA23
F977
F8F9
F99C
F9F5
F8B9
F7AB
F9FD
FFEC
05BD
07E7
06FA
0625
06C8
075B
06A7
0604
0707
0841
065D
00A7
FAA2
F82E
F92B
FA60
F9EF
F925
F992
FA49
F98A
F830
F961
FE64
0461
0770
0705
05F2
064E
0723
06CB
05E9
0661
07CB
0718
0272
FC31
F881
F8A9
FA20
FA45
F96C
F948
F9C6
F955
F819
F8C1
FD20
0332
0706
073C
061A
0608
06B1
0686
05D4
064B
07B7
0733
02CF
FCAF
F8EE
F8E4
FA17
FA0A
F945
F994
FA9D
FA47
F878
F845
FC3D
02A5
0718
078F
0633
05E4
06A5
06A3
05B4
05AD
071E
077D
041A
FE00
F949
F876
F9E6
FA84
F9B7
F941
F9F1
FA58
F971
F903
FBBB
0155
064F
07D4
06CD
0613
06A0
070A
0676
061D
06FD
076C
04C5
FF34
FA35
F8A3
F992
FA24
F970
F90C
F9D5
FA4A
F92A
F83F
FA9D
0059
05C8
07A5
06AF
05F9
06AF
073E
0687
05E7
06D9
07E5
05F2
0087
FB03
F8C9
F97F
FA2F
F977
F8CA
F97B
FA55
F98D
F825
F960
FE81
0494
079A
0706
05C3
060F
0706
06DC
0601
0652
0797
06DE
0240
FC02
F85F
F89F
FA0D
F9EE
F8CD
F8BC
F9A8
F98B
F831
F891
FD0E
03A0
07A9
0764
05A0
059B
06F6
0749
0654
0648
07BD
07CC
03AA
FCF8
F86A
F843
FA12
FA79
F969
F912
F9DB
F9CE
F84A
F80A
FBE4
0284
075A
07DC
061F
0598
06B9
0756
0697
063D
0768
07F3
04DD
FEA0
F955
F811
F993
FA7B
F9B3
F8F8
F972
F9C9
F8C7
F830
FB05
0121
068E
07FD
0686
059C
066C
070F
0645
05AA
06DA
0804
059D
FF6F
F9B0
F81C
F9A1
FA7D
F976
F8C4
F9DC
FAE4
F9C5
F82E
FA01
FFEC
05DB
07CF
0688
05BB
06CB
079B
0694
0565
063E
07CF
065E
00D3
FABA
F831
F92D
FA55
F9C0
F8D5
F942
FA18
F983
F848
F984
FE81
0479
078E
0733
062B
0685
074D
06E8
0605
0682
07E8
0722
0277
FC5E
F8EC
F916
FA17
F994
F878
F8C4
F9F7
F9CF
F849
F896
FCFB
0340
06FF
06E6
05C1
063C
0786
076E
0639
0636
07A3
0770
033D
FD10
F93F
F93D
FA60
F9F9
F8AD
F8A7
F9D4
FA0F
F8D6
F8D0
FC72
0254
0685
072C
0638
0639
071B
0726
062C
05E4
06ED
0719
03FB
FE66
F9EE
F8CC
F99C
F9C3
F8ED
F8C7
F9D2
FA65
F977
F8F3
FBA7
0142
0617
0760
065E
062D
0769
07EB
069A
055F
061E
073D
0541
FFAE
FA36
F857
F944
F9A5
F865
F7AC
F8EF
FA6C
F9F1
F8C2
FA6B
FFD3
0589
07CA
06E5
0616
06F4
07ED
0763
0658
0694
0746
058E
0081
FAF3
F84F
F8C0
F9A6
F955
F8BC
F923
F9CF
F94F
F865
F9D3
FEBE
0496
07BB
078A
0685
06A6
0730
06B7
05E4
0681
080D
075A
0280
FC02
F852
F8AD
FA21
F9DF
F8A8
F8C3
FA01
FA10
F89A
F8BE
FD12
038C
0779
0721
0580
05D2
0778
07CA
068F
0632
077F
0797
039F
FD23
F8BC
F89B
FA54
FA9F
F97D
F91B
F9DC
F9D1
F85B
F823
FBE5
0250
0701
0789
05E9
0563
0659
06C4
05FF
05D9
074F
080A
04F6
FEB3
F98C
F884
FA0A
FA97
F965
F8C0
F9E5
FAE0
F9BE
F83F
FA2A
000C
05D5
07A3
0647
0583
06BC
07B6
06A9
053F
05D8
0748
05C8
0044
FA73
F867
F9B4
FAB1
F9AC
F890
F92E
FA3E
F9AD
F88B
FA45
FFC6
058D
07B9
0696
0587
063A
070F
0675
05A1
0677
07E1
067E
012C
FB19
F838
F8CB
F9DD
F996
F922
F9EA
FAD5
F9F6
F832
F904
FE13
0482
07FA
0794
063F
0674
0758
06F5
05C3
05EE
0777
0739
02D4
FC48
F809
F7E9
F989
F9FA
F942
F92E
F9EC
F9DD
F8C7
F926
FD11
02FC
071A
07AD
0687
0614
0674
066D
0609
0681
07A0
0703
0305
FD5A
F97B
F8CC
F992
F9B7
F946
F95A
F9D2
F97F
F88F
F92A
FCE4
0245
061B
06F9
0664
065D
06E9
06D7
061C
0610
0710
072E
043B
FEC7
F9F9
F843
F8F4
F9A7
F94C
F8E5
F96F
FA4D
FA47
F971
F912
F9C4
FA91
FA61
F988
F941
F9E3
FA73
FA1E
F961
F93B
F9B7
F9FD
F9A9
F95D
F9B1
FA33
FA09
F93F
F8CF
F94A
FA10
FA3E
F9E8
F9DC
FA5D
FAB9
FA5E
F9BA
F9B2
FA61
FAF7
FAD5
FA5B
FA3F
FA84
FA87
FA0E
F9AE
F9E7
FA43
F9F7
F94F
F9E4
FCF2
01B0
05C7
0782
0748
06C3
06F3
077A
079B
0755
0731
075E
0779
0740
06FE
071B
0777
0790
073D
06E7
06EC
071B
0705
069B
0646
0651
0693
06C0
06D6
06FC
0727
0713
06BB
067A
06A3
0708
0737
0713
06F3
070E
071C
06BB
060F
05AE
05DB
0630
063A
0619
063F
0697
067E
05C2
053E
05E4
072C
0718
0431
FF4B
FAEA
F8E4
F8F2
F98C
F9BA
F9A9
F9CC
FA05
F9EA
F976
F908
F8DF
F8DC
F8D9
F8E7
F91C
F959
F96C
F95B
F95E
F98E
F9C2
F9D8
F9E8
FA17
FA53
FA67
FA51
FA45
FA59
FA55
F9FD
F977
F930
F961
F9C3
F9EE
F9D6
F9CA
F9E9
F9ED
F99C
F953
F9A8
FA95
FB49
FB19
FA67
FA31
FAB3
FAFB
FA3B
F943
FA0B
FD89
026A
0639
07A7
0751
069E
0652
065E
0685
06BE
06FB
0713
0706
0713
0758
079B
07A1
078B
079E
07CB
07BF
0764
070E
0702
0717
06F5
0696
064A
0637
0620
05D4
058E
05AF
0630
069B
0699
0656
063E
067D
06DA
070C
0715
0734
0773
077D
06FF
0639
05E2
0656
0705
06FB
0617
0560
05BE
067E
05B7
025E
FDA8
F9FB
F8A5
F8FB
F982
F989
F96A
F9A1
FA1C
FA78
FA76
FA18
F980
F8EE
F8B6
F8F9
F972
F9B6
F99B
F946
F8EB
F8B4
F8BF
F91C
F9AC
FA24
FA54
FA52
FA52
FA63
FA6C
FA64
FA67
FA7D
FA88
FA6A
FA29
F9D2
F96B
F91B
F920
F969
F98D
F949
F8F1
F905
F97A
F9C6
F9C4
FA04
FAD3
FB63
FAB9
F993
FA52
FE5F
0419
082A
08DC
0778
065A
0661
06C1
06B4
0678
068A
06B9
0691
0633
062C
069B
070B
0728
0729
075A
0798
0786
0724
06DE
0706
0765
077F
0725
0694
0620
05E1
05CF
05F3
0651
06B8
06C5
0645
0596
0577
0632
0726
0775
071D
06E0
071F
0746
06CA
0631
0674
0768
07AD
0693
0560
05A6
06A6
05A4
014A
FBB9
F855
F815
F903
F91D
F882
F876
F938
F9DA
F9DF
F9D9
FA40
FA95
FA48
F9C5
F9DC
FA73
FAA7
FA1C
F97D
F96F
F9AC
F988
F8FE
F8B6
F900
F960
F947
F8DF
F8B8
F8F4
F92E
F930
F941
F9B4
FA64
FACB
FA98
FA15
F9E8
FA5E
FB08
FB3C
FAEC
FAA5
FAAF
FA92
F9D2
F8EC
F8F2
F9FF
FAA7
F9BD
F86A
F95F
FDB1
033B
06D0
077C
06E8
06E5
0789
07DD
0786
0718
0711
074A
0773
0784
0775
071A
0692
0663
06BD
070E
06CC
064D
064B
06C0
06E8
066D
05F4
0636
06EA
0730
06D4
0686
06B8
06FA
06C7
0665
0662
06B2
06D3
06A2
0674
0670
0663
0637
062B
0663
0699
0683
0652
0656
0662
061B
05D2
0634
06C8
05A8
01A6
FC38
F870
F7E4
F953
FA5A
F9FC
F914
F8CC
F949
F9E5
FA24
FA09
F9CB
F998
F980
F963
F922
F8F5
F93A
F9C7
F9E8
F950
F8A7
F8B6
F955
F9BB
F9A8
F9B1
FA29
FA71
F9E8
F91D
F941
FA64
FB39
FAE2
FA11
F9DA
FA1D
FA02
F978
F94D
F9DA
FA6E
FA4F
F9A8
F919
F8D9
F8D9
F950
FA54
FB02
FA51
F915
F9FD
FE82
049A
088F
08E3
076A
06A0
0700
075C
06FF
0678
067A
06DD
070A
06D9
0684
0641
0642
06B6
0755
076A
06C7
063D
068F
074D
0768
06B6
0631
068A
072A
070B
0637
05B6
060F
069E
0699
061B
05B8
05A9
05E0
0661
0704
0743
06D9
064C
0644
069E
06B6
0680
0699
071E
072D
0639
0543
0596
0664
051C
00B1
FB62
F84E
F80A
F8B6
F8D6
F8B3
F908
F99C
F9CF
F9B6
F9D6
FA0D
F9C5
F92A
F934
FA1A
FABD
FA42
F962
F947
F9CC
F9DE
F93C
F8C9
F918
F99D
F996
F92B
F911
F965
F997
F96D
F961
F9C3
FA22
FA13
F9DB
F9F2
FA3A
FA56
FA46
FA38
FA1A
F9EA
FA01
FA83
FAD5
FA49
F95A
F952
FA5A
FAD3
F991
F850
FA3F
FFDD
05AD
0809
071E
05F4
065F
0769
0788
06D9
0682
06E1
074E
0757
0742
0744
0716
06B2
069C
0706
074B
06F2
068D
06CF
0749
0700
05F3
053C
0598
067F
06F6
06C6
0682
068A
06A4
0689
064B
0610
05ED
062B
0708
07EF
07CB
068A
0583
05B9
0679
067F
05E8
05E5
06A4
06DB
05D4
04E3
0579
0664
04B8
FFC5
FA94
F874
F932
FA0C
F985
F8B0
F8E7
F9D5
FA54
FA2A
FA04
FA1E
F9F9
F96A
F910
F955
F9B5
F994
F92F
F91A
F941
F92C
F8DF
F8CC
F90B
F94B
F96B
F9A1
F9F8
FA1F
F9E7
F99F
F9AB
F9E9
F9EF
F9C6
F9E0
FA42
FA5F
F9F4
F978
F94C
F93B
F927
F97A
FA44
FAA7
F9EB
F8E0
F909
FA63
FB17
FA26
F97D
FBF5
0176
067E
081A
070C
0624
069E
0775
0795
0733
06D3
0656
059B
053E
05E4
0709
077E
0700
0685
06AF
06EB
069D
064D
06C8
07A7
07C9
06FB
064C
0685
0727
073D
06AA
062A
0636
0670
0653
05F2
05C4
05FE
067B
06EB
06ED
0651
0585
0550
05DE
067D
069D
068F
06C8
06E3
0633
052E
053F
06AD
0766
04F9
FFAC
FA92
F841
F867
F90D
F935
F944
F991
F9C4
F99F
F971
F974
F95F
F907
F8E0
F956
F9ED
F9C7
F908
F8CA
F97F
FA29
F9DB
F91E
F91B
F9D5
FA3A
F9CB
F93F
F961
F9F1
FA26
F9DA
F99D
F9C2
F9F1
F9DA
F9B3
F9C1
F9DC
F9D6
F9D6
F9F7
F9F4
F9AD
F987
F9D0
FA22
F9F7
F99D
F9C6
FA3D
F9E2
F893
F85F
FB88
0169
0682
0826
072E
064F
06B6
0760
074B
06E6
0709
078E
079C
06FF
066A
0675
06E5
0730
072B
06F9
06A8
0653
063B
0671
069B
0681
0664
0686
06A1
065D
05F9
0604
0680
06C8
0680
061C
0630
0690
06AA
0689
06B9
0729
070D
0633
058B
05D1
066E
066E
05F7
05E1
062D
0601
0550
0550
067A
06E8
041B
FE69
F941
F77A
F86F
F987
F98E
F958
F9A3
F9E8
F986
F8E3
F8CE
F948
F9A5
F9A3
F9AB
F9EC
F9F6
F981
F912
F940
F9D0
FA16
F9EA
F9A9
F987
F96B
F94C
F94D
F97E
F9C6
FA0F
FA38
FA0E
F982
F8FC
F912
F9C3
FA3C
F9D9
F929
F93B
F9FD
FA40
F992
F907
F997
FA9F
FAE0
FA63
FA31
FA71
FA22
F928
F96E
FCDF
0277
06CF
07C8
069D
05CE
061C
068E
0682
066A
069D
06B6
0668
0625
0674
0718
0763
0739
0729
0779
07B7
0771
06EB
06AE
06C8
06F2
0705
06EA
0671
05B6
054E
05A7
0654
0680
0601
0580
0598
0619
0679
0699
06BA
06E3
06DD
06CC
0712
077B
0751
0689
0621
06A0
0719
0675
0550
054C
0675
066B
030C
FD5B
F8C7
F784
F887
F965
F934
F8D3
F90D
F997
F9D1
F9A8
F977
F975
F992
F9A1
F98C
F95E
F93C
F93D
F942
F913
F8BE
F8A7
F90A
F982
F97D
F921
F934
F9EE
FA93
FA7F
FA0F
F9FC
FA44
FA5A
FA25
FA12
FA26
F9D0
F92A
F9B1
FCD3
01C5
05C9
0702
064E
05CA
063D
06C4
069F
062D
060E
062B
0617
05F5
064D
071D
079B
0732
064B
05D2
0616
0699
06C8
069A
0669
0678
06AE
06AA
0641
05C7
05BF
062D
068A
067B
0640
0638
063A
05EE
05A3
061E
0723
06D2
0369
FDC7
F91F
F7C7
F8DD
F9C1
F93F
F867
F88C
F970
F9F1
F9B5
F96B
F995
F9D7
F9B0
F954
F944
F983
F9A3
F985
F973
F996
F9AB
F973
F918
F8FE
F942
F990
F988
F933
F905
F952
F9DD
FA1E
F9FA
F9EA
FA4A
FAA3
FA24
F919
F965
FCB9
023A
06D0
082A
0709
05F7
0647
0714
0716
0674
0643
06C6
071F
06B0
060A
060A
06A1
06FF
06C5
065B
0636
0644
063E
062A
0644
0687
069A
064B
05EF
0606
0695
0700
06C7
0631
05F4
0648
068F
063D
05C5
0623
0734
071A
03FD
FE7A
F983
F786
F827
F935
F94C
F8DD
F8CB
F915
F926
F8F6
F90C
F985
F9CD
F98C
F940
F98A
FA2C
FA59
F9D5
F944
F943
F9A5
F9C5
F96A
F903
F914
F97F
F9AD
F95A
F8F8
F91B
F9A6
F9EC
F9A7
F96D
F9D3
FA64
FA0B
F8DF
F8DB
FBF2
0175
0641
07E0
06F2
05F2
063A
0700
070F
0673
0618
0658
06A3
067D
062D
0633
0681
06A6
067D
0651
065D
068A
069E
0685
065E
065C
068C
06A9
066B
0601
05F0
065A
06C2
06BA
0684
069C
06D9
0698
05E2
05B7
068B
06D9
046B
FF41
FA2E
F7F1
F85E
F92A
F8EB
F84B
F864
F91C
F988
F956
F915
F92E
F958
F93D
F917
F94D
F9C2
FA04
F9E9
F9A4
F962
F93B
F942
F96F
F991
F997
F9A5
F9C4
F9BB
F972
F930
F934
F94F
F93C
F942
F9E1
FAC4
FAB8
F970
F8DF
FB7B
00FD
060F
07E4
0724
0677
0702
07A2
073C
0669
0649
06C9
06E9
0665
060C
065F
06C2
0689
0610
061E
06AF
070A
06D4
0664
062A
063D
0678
0699
0679
063F
064E
06B3
06ED
0690
05F0
05BF
0610
062A
05C6
05BF
06A7
070C
0490
FF29
F9F7
F7EE
F8AA
F989
F937
F8B0
F914
F9DC
F9DE
F92B
F8DC
F95B
F9E1
F9C8
F977
F98A
F9CC
F9C0
F985
F986
F9AE
F9A7
F986
F9AB
FA0A
FA37
FA08
F9BB
F987
F96F
F972
F998
F9C6
F9C1
F99E
F9CE
FA44
FA14
F8D0
F81D
FA80
000C
0582
07AF
06DE
05D5
0631
0703
06F3
0648
0630
06DC
075D
0725
06B4
0690
0682
0643
0623
066D
06B8
0682
0612
05F6
061D
0613
05D4
05D0
0624
067A
0697
06A1
06C1
06D3
06B5
068D
067D
064B
05ED
0601
06DE
0723
049F
FF3E
F9F6
F7C8
F887
F99C
F964
F898
F888
F932
F9A9
F990
F95E
F964
F96E
F96D
F9B5
FA33
FA33
F976
F8D9
F928
F9F4
FA2B
F990
F8D8
F8A2
F8ED
F963
F9AB
F984
F905
F8B8
F918
F9E0
FA3C
F9E3
F98D
F9D6
FA20
F995
F92C
FB29
0010
0547
07CD
077D
0696
0699
0703
06E0
0662
0653
06C1
0702
06CE
068B
0683
0675
063A
0629
0666
067A
061B
05C6
05FE
0670
0681
0635
05FE
0602
0623
0664
06C9
06FC
06B6
065B
0693
072E
071D
0610
0562
0649
0755
0575
FFFD
FA30
F7AD
F878
F9B3
F983
F8A8
F87C
F8FA
F93E
F909
F8E8
F924
F964
F96D
F981
F9CA
F9F3
F9BF
F983
F990
F9B0
F9A9
F9A2
F99F
F94C
F8C6
F8CF
F9A1
FA3E
F9C0
F8C9
F8BB
F9AA
FA38
F9A4
F8FF
F979
FA50
F9F7
F91A
FA96
FF9C
0578
087B
0814
06AD
064A
06C0
070D
06EE
06B5
068A
0669
0674
06AF
06B1
062E
05AD
0601
06E8
072B
065B
0593
05CF
068A
06C0
066A
0621
05FB
05BC
059A
05F0
0665
0657
05ED
05FA
0690
06A5
05BB
051A
0607
0722
0568
0043
FAE5
F892
F8FE
F9A7
F975
F947
F99A
F9A2
F8F3
F883
F935
FA4B
FA5F
F971
F8EA
F97E
FA32
FA09
F978
F973
F9E5
FA13
F9D8
F990
F95D
F94B
F9A7
FA63
FABD
FA33
F978
F98D
FA36
FA3D
F96D
F91E
FA15
FAD4
F9AA
F812
F9B3
FF75
0589
07D1
06B1
05B7
0695
07A7
072F
05F0
05B5
06A4
0746
06CF
0614
0608
0671
069D
0688
068C
0693
066A
064B
0666
066B
062A
060D
064F
0665
05EB
058D
061A
0708
06F7
05C2
04FF
05D4
072C
0736
0635
0611
06E1
05F6
0178
FB84
F807
F830
F9A4
F9EF
F91B
F89F
F907
F98D
F981
F91C
F8E7
F902
F949
F995
F9A1
F931
F8A8
F8D4
F9AF
FA23
F98B
F8C7
F8F9
F9DB
FA40
F9C7
F93D
F942
F97F
F95F
F901
F8EC
F929
F955
F960
F989
F9A0
F94D
F94D
FB4C
FFB3
047D
073B
07A4
074E
074E
0747
06C8
065F
06B8
0762
0758
068E
0613
0673
06ED
06AC
0612
05FE
066A
068E
0630
05F3
064F
06E9
0713
069C
0604
05EA
0673
071F
074E
06EA
0687
06B0
0718
06DF
05EA
0570
065E
0758
059A
0069
FA9C
F7BC
F834
F95B
F919
F828
F85D
F9B8
FA73
F99A
F869
F880
F9B3
FA73
F9FF
F929
F8F9
F95B
F98B
F944
F903
F92D
F974
F94C
F8D4
F8D8
F9BE
FAC2
FABA
F995
F89C
F8F7
FA3C
FAEC
FA59
F977
F976
FA11
FA18
F99E
FA87
FE3A
0371
072A
07D4
06B6
0614
0696
0726
06E9
0674
06B2
0767
0773
067B
0580
059B
0698
073A
06BD
05B8
0550
05E2
06B1
06E7
0687
0634
0647
0676
066B
0647
0657
068B
068A
0641
0608
061E
0646
0638
0625
0665
0681
052A
0195
FCBD
F8D6
F770
F83D
F9AA
FA5F
FA1C
F96E
F8F6
F8F5
F948
F98F
F988
F954
F95C
F9CD
FA47
FA43
F9BA
F939
F935
F98D
F9BE
F991
F94D
F94B
F985
F9A8
F991
F96E
F96F
F977
F952
F922
F951
F9F4
FA74
FA18
F91B
F8E8
FAEA
FEFB
0352
061D
0705
06FF
06ED
06D4
0676
061B
064A
06ED
073A
06C1
060E
05FC
068F
0704
06DE
0683
068D
06E2
06EA
067D
0637
0694
0724
06FF
0605
052C
0560
0659
06E6
065F
0574
0550
0624
06F4
06ED
0672
066F
06B0
05A4
021B
FD01
F8DE
F77D
F861
F9A2
F9EC
F967
F8E9
F8DA
F91D
F981
F9D9
F9D6
F949
F887
F84B
F8F4
F9FF
FA77
F9E6
F8E1
F870
F905
F9FF
FA59
F9C5
F905
F903
F9AA
F9FE
F98D
F97F
FB94
0000
04C5
078D
07CE
06D0
0603
05D5
060E
0684
0718
075A
06E0
05FF
05A6
0644
072A
074D
0680
0592
0566
061D
0706
073D
0682
0595
0586
066E
0733
06DB
05E4
05A4
063C
05D2
0291
FD2E
F8A4
F72F
F838
F989
F9D3
F958
F8CB
F877
F884
F923
FA17
FA93
FA09
F903
F8AC
F971
FA77
FAA3
F9E0
F917
F923
F9F3
FAA6
FA5C
F92D
F84E
F8CE
FA1F
FA7F
F953
F87E
FA94
FFC1
0537
07F9
07B2
0667
05D1
05F3
062A
0667
06D2
06F7
0658
057D
0586
06AD
07D1
07C2
0696
0587
0596
0685
072F
06C7
05B9
053A
0603
0761
07D7
06D3
058E
059B
06A0
0651
030B
FDE3
F994
F7DF
F867
F9BA
FAA2
FA8D
F984
F841
F7DC
F8C3
FA0B
FA43
F926
F7F6
F7F8
F90E
FA10
FA2E
F98E
F8E7
F8E9
F9B6
FA9E
FA9E
F991
F898
F8D0
F9D3
FA24
F952
F90A
FB62
003C
051A
07A6
07C6
06F2
064D
0605
0607
0651
06AF
06B7
064A
05C3
0597
05EF
068B
06F0
06B7
05EC
053B
0560
0649
06EE
0692
05DE
0614
0729
0798
0697
0572
05C9
06FC
0678
02C3
FD6C
F974
F854
F90B
F9CC
F9D0
F960
F8E3
F890
F8A7
F94A
FA0D
FA37
F999
F8D9
F8CA
F97F
FA25
F9CF
F89A
F7CE
F890
FA63
FB69
FA7F
F8C2
F864
FA00
FBA4
FB20
F8EA
F804
FABE
002A
0525
076D
073D
0638
059C
05A2
05FC
065B
0688
0653
05CA
0561
05A8
069C
076D
0740
063B
0581
05F5
071E
0797
06B1
055F
051A
0617
0717
0709
065C
063B
06E8
0747
05F4
028A
FDF1
F9CF
F793
F79C
F909
FA5C
FA93
F9C9
F8E0
F8A1
F925
F9E9
FA3F
F9CC
F8ED
F890
F942
FA5D
FA97
F9AF
F8E0
F952
FA77
FAB2
F980
F83A
F866
F9BD
FA75
F97C
F7F7
F837
FB64
005C
04C6
0700
0729
069C
0676
06B3
06B2
065B
0640
069E
06E5
0699
061D
0622
0697
06C3
0670
064B
06D3
0767
0705
05D6
0537
05EF
070F
0716
05E7
04EB
0561
06E9
07C1
0648
025F
FD9A
FA04
F88C
F89F
F92E
F9AE
FA04
F9FF
F973
F8D5
F8FC
F9F4
FA84
F999
F7F8
F788
F8BF
F9E5
F96B
F81D
F803
F98C
FB04
FACC
F94B
F842
F8B3
F9E6
FA6C
F9AB
F874
F861
FA9E
FEE9
038D
06A9
07B7
078F
070B
0657
05B5
05D8
06D2
0785
06FC
05E6
05C2
06BE
0761
06A7
0587
05A0
06DD
0785
06B6
05A8
05D4
06E9
0767
06C2
05E4
05D8
06AA
0792
078C
05DB
0287
FE81
FB0C
F8DF
F7F5
F803
F8CD
F9D3
FA3A
F99A
F8C5
F8EB
F9E9
FA52
F980
F8A0
F8FC
FA0F
FA58
F98F
F8FB
F98B
FA8C
FAA9
F9A7
F899
F888
F95C
FA2E
FA3B
F975
F894
F8E2
FB54
FF77
0392
062F
0725
070F
066B
05B7
05A6
066F
0735
06FC
0608
05A4
0661
073D
0702
05FD
05A2
067E
0771
0742
062B
0558
0569
060E
06A2
069E
05E4
0523
0571
06DE
07D0
066B
02A2
FE4F
FB30
F97C
F893
F85F
F91A
FA1E
FA25
F919
F877
F941
FA86
FABE
F9F3
F96D
F9BE
FA2D
F9FE
F978
F94F
F99F
F9ED
F9DB
F97F
F91E
F8F9
F950
FA08
FA60
F9AF
F8AF
F932
FC14
0027
03A6
05F2
0745
078A
069B
0556
0532
066C
0785
071E
05CD
0548
0604
06AE
0637
0560
057C
0682
0735
06E3
0610
059D
05DC
0677
06BB
0622
04F5
0452
0515
06B4
076F
05ED
0280
FE97
FB56
F91B
F822
F89E
F9EA
FA9D
FA0E
F928
F91A
F9C1
FA13
F9B6
F950
F966
F9A7
F99F
F97D
F9B0
FA1D
FA34
F9D2
F972
F965
F972
F976
F9BF
FA56
FA90
F9F4
F929
F974
FB6C
FEB0
0274
05D5
07D2
07CC
0657
0519
0543
065A
06EF
067B
05D5
05CB
061A
062A
0614
0643
0695
0696
0644
0606
0600
0605
0623
069A
0729
0702
05F2
0517
05B3
0745
07B2
05A8
01FF
FE6E
FB9E
F957
F7CF
F7B4
F8E2
FA13
FA38
F996
F932
F972
F9D8
F9F8
F9F8
FA07
F9ED
F988
F941
F979
F9EC
FA0E
F9C9
F96E
F926
F8F2
F904
F996
FA50
FA67
F9A1
F8EA
F988
FBCD
FEFE
025A
0577
07A1
07EB
067B
0508
052F
0693
0772
06EA
05F1
05CD
0664
06AF
0663
0645
06CB
0750
070F
0648
05D0
05EB
062F
0648
0637
0604
05B6
0597
0603
06C6
06FA
05C4
031A
FF9F
FC15
F92C
F7B2
F81A
F9AC
FAD7
FABC
F9F6
F985
F98F
F9AE
F9CF
FA19
FA3C
F9B7
F8CD
F87D
F92D
F9F8
F9CB
F8E7
F88C
F929
F9D8
F9DC
F9A3
F9C4
F9DB
F94C
F8A0
F919
FB3F
FE74
01E1
0504
074C
0802
071D
05CE
057D
0646
0703
06F7
068A
0649
0616
05D1
05E7
0685
06F1
0687
05CD
05B1
062E
0678
0662
0690
0728
073A
0637
0546
05FA
07D7
087C
0696
0348
001C
FD0F
F9C4
F761
F771
F96C
FAE3
FA61
F8F1
F86D
F91F
F9DF
F9F2
F9B6
F993
F958
F904
F91B
F9A3
F9CE
F94C
F8FC
F97F
FA00
F98A
F8B7
F8DB
F9E5
FA5C
F993
F8BB
F94C
FB42
FDBD
00B0
047C
0804
0906
071D
04E2
04E2
068B
076F
06B2
05AB
059B
063A
06B6
06E6
06FD
06D3
0644
05D5
062E
06F1
0712
066F
0615
0685
06E4
0686
0628
069D
0738
06BD
0523
0340
010F
FDC1
F9B1
F707
F76E
F9D5
FB5E
FAA2
F8EA
F824
F8A7
F990
FA2B
FA35
F98D
F8A3
F88D
F9AE
FAD7
FA9F
F947
F855
F88C
F929
F956
F966
F9F1
FA73
F9EB
F8AA
F84B
F992
FB94
FD94
004A
0438
07D0
08D9
0747
0569
052F
0645
071D
06EF
0632
05A0
057F
05D8
0694
0728
06EF
0612
058B
05CC
0648
0693
070D
07C5
07C5
067E
0528
057A
0735
082E
0708
04C6
02EB
011A
FDDD
F99C
F6FC
F7A3
F9F0
FB07
FA36
F90D
F8D3
F939
F97A
F97F
F993
F9B1
F9A3
F977
F961
F959
F93A
F928
F95F
F994
F946
F8C6
F903
FA09
FA9B
F9E8
F8DC
F8DD
F9FC
FB6A
FD3A
005F
04A8
07FA
0874
06D2
05A2
0627
072B
0722
0654
0603
066C
06B9
0680
0648
0681
06E0
06EE
06AA
066A
065D
0683
06D0
0710
06DA
060A
0543
055B
0635
06CB
068A
05BF
0471
01BF
FD55
F8DA
F6B3
F769
F919
F9BF
F944
F8E3
F92A
F974
F941
F904
F934
F977
F951
F90D
F941
F9CB
FA04
F9C3
F973
F951
F92D
F8F0
F909
FA14
FC4F
FF84
0329
0651
07DE
0778
0645
05F2
06CE
0792
0745
068B
066A
06B3
0689
0604
061E
070B
07A6
06F6
05A8
0538
05FD
06E8
072E
0735
0758
06C2
045A
0062
FC53
F977
F822
F80F
F8BD
F97A
F9B4
F971
F929
F91C
F91D
F90E
F93A
F9CB
FA32
F9D7
F92C
F938
F9EB
FA00
F8F5
F807
F863
F954
F979
F94D
FAFE
FF70
0491
0775
0787
06AC
0678
0697
0637
05C3
062F
073C
07A5
06DA
05AA
0536
05C4
06AC
070B
068B
05B9
0581
062E
0705
0723
069C
0646
0625
04BC
00D7
FBB1
F83D
F7E3
F91A
F9B3
F980
F9A8
FA42
FA24
F8F2
F808
F8AE
FA36
FAD1
F9EE
F8DC
F8DF
F98C
F9AC
F90C
F89F
F8FD
F99D
F9A8
F932
F972
FBC0
0024
04CF
0779
077A
064D
05C7
0636
06AA
06A4
06BE
0764
07D6
0725
05DA
0586
0685
0752
06AC
0572
0564
069C
0770
06CB
05A8
05A7
06BF
06FC
0495
FFE8
FB2E
F87F
F830
F907
F9A0
F98D
F949
F93E
F924
F8A0
F823
F877
F960
F9A0
F8B6
F7D9
F869
F9E5
FA7D
F992
F8A2
F933
FA8E
FAAD
F940
F8A2
FB32
0061
0538
076E
0744
067C
064E
06A6
06DF
06BF
069B
06C2
06FB
06DC
0670
0646
06B0
0735
071F
067C
062E
06A9
0724
069E
0592
0594
06F5
0790
04F9
FF81
FA43
F7FF
F88B
F9AD
F9CE
F93D
F8F0
F90D
F90E
F8E0
F900
F982
F9B4
F907
F7FF
F7BD
F89E
F9AD
F9C4
F8FF
F89C
F954
FA3B
F9EC
F8A9
F8A4
FBB0
00F8
0591
075B
06E3
0636
066C
06E2
06B1
061F
0613
06A6
06F9
0687
05FB
0648
0741
07BF
072B
065F
068B
0783
07D8
06CC
058B
05BD
070B
06F9
03A1
FE22
F9B8
F86D
F94A
F9F0
F964
F8A3
F8CC
F98D
F9CB
F944
F8D0
F913
F9A0
F9AE
F946
F928
F996
F9D4
F92E
F82A
F81E
F966
FA9F
FA36
F8AA
F882
FBA8
0121
05DF
07BE
0747
0681
0692
0700
0703
06B4
06AF
06FC
0702
067F
05FF
061C
06AB
06F4
06B5
0682
06F0
0799
076D
0632
052A
05AB
0714
06E9
0374
FDF4
F9A1
F86C
F94C
F9DE
F93B
F877
F8A3
F94B
F960
F8D5
F891
F903
F996
F9A5
F95E
F95E
F9A8
F995
F8D5
F81B
F873
F9D4
FAE3
FA68
F907
F91F
FC7F
0232
06F0
0839
06D2
05A5
0650
07A2
07B5
068E
05D0
0654
0732
0746
06C3
069C
06E9
06D7
0625
05BE
065A
0732
06EA
0584
0490
053C
06AA
0688
0359
FE18
F994
F7F2
F8D2
F9FC
F9D5
F8DD
F894
F95C
FA06
F985
F860
F7F6
F8A4
F976
F9A3
F97A
F97C
F96A
F8E9
F886
F91C
FA4D
FA9B
F95E
F81E
F94B
FD9A
0311
06D4
07B8
06E0
0634
068A
0742
0749
0673
05B8
0613
073F
07FF
07A7
06CC
064E
0643
064E
0677
06F0
0745
06AA
055E
04F8
067D
0867
07A9
030B
FCDB
F8AF
F7E4
F8EB
F987
F90B
F861
F891
F993
FA66
FA26
F90E
F83C
F872
F93F
F993
F912
F877
F88D
F92A
F99A
F9B8
F9DF
F9E2
F928
F839
F923
FD4B
0333
077A
0848
06F4
0616
0697
0733
069F
0548
04AE
0585
0703
07CF
0749
0603
0542
05D6
0742
082C
07D0
06B7
05F3
0601
06A9
077C
07C7
065A
0257
FCB0
F837
F740
F924
FAE3
FA78
F8DC
F853
F96B
FA96
FA68
F94B
F8B1
F941
FA3E
FA8D
F9E6
F8EB
F865
F89E
F954
FA01
FA2A
F9A3
F8C3
F86F
F9CA
FD72
0294
06F6
0892
0787
05FA
05CC
06BA
0729
0675
05B3
060A
070C
074F
065F
0561
0592
06BA
0796
0761
0677
059C
0540
057F
0656
0765
07A0
05C1
0173
FC28
F85E
F7A4
F92D
FA99
FA47
F8D6
F82D
F91D
FA70
FA77
F930
F831
F899
F9BB
FA3D
F9CC
F937
F925
F96A
F9A4
F9D5
FA05
F9D8
F91B
F8B6
FA44
FE56
036F
0728
0845
077D
0679
064F
06E3
0757
070C
064C
05F0
065A
06F2
06DF
0626
05B5
063C
073D
07AC
073F
069C
0654
064C
0653
0682
0681
0516
0160
FC69
F8B3
F7CB
F8C1
F970
F8F5
F84B
F891
F97F
F9F4
F973
F897
F846
F8DC
F9FE
FACF
FA8C
F951
F82A
F822
F92B
FA39
FA5E
F9A5
F8D7
F8E1
FA91
FE59
0387
07F1
0961
07DE
05DA
0592
06CE
07B8
076E
06C4
06B5
0706
06DE
0628
05A3
05D1
0667
06EA
0734
072A
0699
05C5
0596
0686
07A9
0753
04B2
007D
FC3F
F953
F84A
F8C6
F9A4
F9C7
F90B
F857
F881
F943
F99F
F945
F8E2
F906
F95F
F967
F93B
F93A
F94E
F941
F95F
FA00
FA99
FA19
F89F
F822
FAA2
FFC3
04D8
0778
0792
06BE
063F
0636
0650
065F
0656
063E
063A
0668
06AF
06E0
06EA
06D4
069A
0650
064F
06DA
078D
0784
0689
05A9
05E4
0654
04B3
0030
FAF8
F81D
F85F
F9CF
FA6D
FA1D
F9EF
FA43
FA70
F9EF
F928
F8D5
F917
F989
F9DB
F9F8
F9C8
F941
F89E
F848
F877
F90C
F997
F985
F8C4
F865
FA2A
FEC3
047F
085E
08C3
06EE
0579
059F
0679
06B8
0645
05E7
05F5
0629
0653
0689
06B2
0681
060A
05E7
0679
073B
0745
067F
05E5
066D
07AE
07F5
05C0
012C
FC12
F8BB
F827
F961
FA82
FA82
F9D9
F975
F985
F98E
F958
F932
F954
F97A
F965
F959
F9B8
FA31
FA09
F93E
F8CE
F95E
FA1C
F9A1
F809
F76F
F9E7
FF24
0472
0729
06EE
059C
0525
05D5
069B
0697
0609
05C7
0620
069B
06B7
068F
068A
06A2
067C
062B
0647
06F9
0771
06E0
05CA
05B3
070F
0812
063F
013C
FBA1
F88F
F8BC
FA38
FACC
FA22
F974
F9AF
FA6C
FAA8
FA1D
F973
F94E
F988
F997
F969
F972
F9E8
FA54
FA3A
F9D7
F9D7
FA32
F9F9
F8C1
F7E5
F99D
FE70
041A
077C
0799
0636
0597
0625
0699
0600
04FC
04D3
05C9
06D9
0701
0661
05E3
060B
0671
0665
05D9
055C
0555
0591
05C2
0613
06B3
06DC
0512
00D6
FBD8
F8C1
F8A2
F9F8
FA7A
F998
F8B4
F916
FA51
FAF0
FA4B
F91F
F889
F8E0
F9AB
FA4B
FA83
FA6C
FA39
FA09
F9E8
F9D4
F9BD
F996
F994
FA50
FC7C
0035
046A
0750
07D2
06A9
05A8
05E1
06BC
0711
06A0
061D
060A
062B
0629
0629
0673
06CF
06B2
060F
057E
0574
05B3
05DE
0619
06A8
070C
0617
0327
FF0E
FB8E
F9D6
F98D
F960
F882
F78C
F7B6
F946
FB02
FB67
FA50
F914
F8E3
F96F
F998
F923
F8FB
F9AE
FA80
FA85
FA04
F9F6
FA61
FA3B
F936
F8E4
FB47
0043
0543
07AD
0754
0628
05EF
06BA
076C
072B
063F
05A0
05E5
0694
06C0
0641
05F6
0694
0785
0788
065E
0542
053F
0586
042D
00A4
FCA4
FA43
F9AA
F964
F885
F7B8
F7F8
F90E
F9CA
F986
F8ED
F911
FA09
FACD
FA7E
F970
F8CB
F92A
F9DF
F9CC
F8FB
F90B
FB9D
0055
04E4
0733
0738
0674
061F
0644
066D
068B
06D2
072A
072C
06C1
065E
0677
06E8
071B
06B4
0601
05B4
0639
0714
06F1
049F
004D
FBB2
F8B5
F7E6
F860
F8F5
F933
F953
F98A
F9B9
F9B4
F987
F95F
F956
F968
F984
F98E
F97A
F96D
F980
F97F
F935
F937
FADA
FECB
03C4
0749
07F0
06AE
05AC
05F7
06C9
0704
06A9
0698
0729
07BD
079E
06E8
0652
0641
0664
0642
0602
065D
077F
0827
066A
01B0
FBD4
F7DE
F754
F8F9
FA57
FA49
F9A8
F996
F9EA
F9B0
F8C1
F819
F883
F987
FA0B
F9BF
F977
F9F4
FABD
FA93
F92B
F813
F979
FDE6
035B
06F1
076D
0628
0560
05DC
0696
067C
05E1
05E5
06CE
07A8
078F
06D5
0675
06B4
06C6
0609
0520
055A
06DC
07E6
0641
0193
FC05
F87B
F814
F970
FA69
FA35
F9AE
F9BD
FA24
FA0F
F966
F8F8
F959
FA0A
FA25
F9A1
F963
F9FA
FAA8
FA2B
F871
F73D
F8B9
FD60
034A
0797
08C1
079C
0637
05DB
0636
0659
060F
05F3
066A
0703
0713
06A1
0649
0645
0613
055D
04D1
0584
0754
086B
06B3
01FF
FC7F
F8F6
F873
F9B8
FABD
FA8E
F9C8
F96C
F9A3
F9C2
F94F
F8AE
F89B
F926
F9A7
F9A9
F995
FA17
FAF5
FB0D
F9D2
F882
F962
FD73
0314
0741
0838
06D6
0560
0537
05F8
068A
0689
066B
0694
06CB
06BA
068D
06AC
06F6
06BC
05BD
04DC
0554
071D
085F
06EE
0269
FCDA
F906
F828
F930
FA21
F9F8
F943
F90E
F990
FA12
F9EC
F952
F8F7
F920
F969
F977
F988
F9FC
FA86
FA49
F90E
F81D
F95B
FD61
0296
0670
07A2
06F5
062E
0653
070C
077B
0746
06C1
064D
05E5
056A
051D
0571
065D
071A
06EB
0619
05CE
06AB
07A3
06A4
02B7
FD4A
F91E
F7E4
F8F0
FA37
FA57
F98B
F8E5
F8F5
F962
F992
F964
F930
F93D
F97A
F9BA
FA0A
FA7D
FABF
FA2B
F8B3
F79B
F8CA
FCF7
028A
06BA
07F3
070F
0624
0651
0707
0740
06E9
06BB
070B
0755
0706
065F
062F
06B4
0733
06D0
05BB
051C
05BB
06D0
0679
0388
FED4
FAA6
F8C1
F8FB
F9C1
F9C6
F913
F87D
F87F
F8D6
F91A
F949
F990
F9CF
F99B
F8E8
F851
F87D
F93D
F99E
F915
F882
F9AA
FD6D
0296
06A2
07E3
06DA
0572
0515
05B1
0666
06BA
06DD
070A
0721
06EF
06A1
0695
06D6
06FE
06BD
0655
0666
0722
07C8
06FA
03D9
FF05
FA7A
F824
F852
F98F
FA25
F9B0
F90D
F909
F96D
F989
F93F
F91C
F969
F9AE
F95D
F8BA
F898
F938
F9D9
F9A9
F901
F968
FC24
00CE
055D
07CA
07B3
0674
05BD
0619
06CC
06FC
06AC
0679
06A8
06DB
06BF
0699
06D8
0749
0738
0677
05DA
0648
0755
0734
0467
FF74
FAB1
F84B
F87C
F9B8
FA57
F9FF
F96F
F94C
F962
F928
F8A2
F869
F8D2
F973
F9AF
F98D
F9A6
FA2A
FA64
F9A5
F884
F8CD
FBCE
00C8
0560
07A2
0784
0683
05FB
0624
066B
0671
0663
067A
068B
064C
05DC
05C1
063C
06E1
0701
0684
0611
0643
06BD
063F
03CD
FFC1
FBB1
F935
F8BC
F964
F9F1
F9D6
F970
F94C
F97D
F9A4
F996
F990
F9C7
F9FF
F9E0
F992
F9A0
FA21
FA4B
F961
F80C
F839
FB4C
0084
056D
07F4
07F4
06D1
05F9
05D7
0602
0609
05ED
05F7
0655
06D2
070C
06D9
067B
064F
0650
0638
060C
063A
06CB
06BC
04B2
0091
FC0F
F949
F8C3
F92B
F914
F87C
F860
F92C
FA26
FA71
FA23
F9F9
FA36
FA4E
F9C2
F8FE
F8E9
F9B8
FA7F
FA3F
F94C
F956
FBD7
0072
0500
075D
073C
0623
05BE
064B
06D0
0690
05F2
05D9
0667
06D3
0674
05A9
055C
05D1
0655
0647
0605
066A
0751
072C
0479
FF9D
FAEF
F8A5
F8D8
F9C5
F9D9
F92E
F8F1
F9A6
FA84
FA86
F9B6
F918
F958
FA05
FA3C
F9D5
F983
F9C8
FA25
F9C2
F8D2
F8E1
FB67
0007
0489
06CD
06AB
05CA
05BC
0678
06DD
064B
0565
0531
05D2
067E
0692
0655
0673
06F7
072A
0696
05CC
05C9
068D
069C
0457
FFE0
FB66
F93A
F9A4
FACA
FAD8
F9D7
F941
F9EA
FAF2
FAF1
F9CE
F8DA
F91C
FA10
FA6E
F9D8
F936
F95A
F9DC
F9BB
F8FD
F91C
FB95
0020
04A5
0703
06DB
059E
0500
0578
062E
0635
05A3
0553
05C2
067A
06B9
066F
063F
067D
06A9
0633
0588
05B8
06DB
074D
052A
008F
FBDD
F981
F9A5
FA68
FA2D
F939
F8E2
F9A7
FA9E
FAB2
F9F5
F960
F98F
FA17
FA3C
F9EF
F9C8
FA20
FA78
FA07
F8E6
F871
FA40
FE8B
0393
06EA
0775
0646
055B
05A9
0675
0698
05FF
059A
0603
06B1
06CB
0652
060A
064E
0687
0623
05A5
061A
0771
07E7
0598
00A7
FB73
F88B
F888
F9E7
FABD
FA63
F98C
F927
F95E
F9B3
F9C0
F9A7
F9B8
F9E5
F9C9
F948
F8EF
F952
FA22
FA5B
F99C
F922
FAD0
FF13
0403
06F9
0707
05AE
0516
05E9
0711
0753
06AE
0610
0613
0669
0683
0664
0687
06FC
071C
0657
0532
04EE
05F7
06E7
058E
0144
FBF3
F88C
F857
F9F9
FB1B
FABE
F9BA
F946
F98D
F9D2
F99B
F93E
F93E
F985
F998
F961
F970
FA25
FAEA
FAA3
F923
F7F4
F943
FDB7
036B
0758
07F9
067E
0558
05CF
0717
07B4
073C
068B
066B
06A0
0677
05E5
059F
060F
06A8
06A2
062A
0644
074F
07FD
0656
01D5
FC59
F89B
F7D6
F8EA
F9D4
F99F
F8E3
F8AB
F939
F9F1
FA36
FA0A
F9D6
F9BE
F978
F8DC
F862
F8B3
F9B3
FA49
F9A0
F897
F96F
FD82
035D
07BA
0891
06F5
059E
05F6
0703
0728
0636
056A
05B6
06B2
0763
0772
074E
074B
072B
069D
05E1
05A6
062E
06A4
0589
020C
FD27
F92C
F7E0
F8ED
FA51
FA71
F98F
F909
F96A
F9D9
F982
F8CF
F8C6
F97B
F9ED
F979
F8D8
F917
FA09
FA65
F99F
F8FA
FA58
FE17
0296
05C1
06D0
0689
061E
062E
069A
06F3
06FC
06CA
0699
067B
0642
05DD
05AA
0616
06E2
072F
0691
05D8
0629
0734
06EF
03B5
FE75
FA1B
F8A9
F969
FA2F
F9EB
F94B
F935
F97F
F983
F94A
F972
FA10
FA76
FA27
F97C
F8F9
F8AB
F898
F984
FC58
00B6
04C9
06E8
071E
06AA
0661
061D
05B6
0593
05F6
0669
0665
062A
0646
0688
0647
05B7
0604
076E
07FF
0557
FFCF
FAAC
F8BA
F972
FA36
F9B7
F901
F956
FA4B
FA95
F9F5
F94D
F929
F932
F929
F96B
F9FE
FA0B
F937
F8F9
FB58
0032
04C6
0693
05FE
0568
0615
0710
0715
0663
05FF
0615
060E
05E9
063A
06EB
0705
0643
05E2
06C8
0777
053A
FFC5
FA4B
F828
F936
FA87
FA3C
F941
F92C
F9C4
F9C2
F915
F902
FA01
FAE9
FAB2
F9ED
F99D
F97C
F8C0
F841
FA31
FF2C
04A6
076A
0728
0650
06A3
074D
06E3
05CA
0586
0650
06DD
0676
05EA
0602
0629
05A6
0547
064C
07C9
06C5
01E5
FBC0
F84B
F880
F9D9
F9EF
F912
F8D5
F95C
F985
F91D
F942
FA55
FB03
FA3D
F8FD
F8E5
F9C1
F9F3
F962
FA53
FE69
03E8
074B
075E
063D
062D
06E5
06DF
061B
05FD
06E5
0776
06B7
0596
0570
060A
0635
05F3
0668
0753
0649
01AF
FB85
F7BD
F7DE
F9AD
FA57
F9A2
F927
F977
F99A
F91E
F8FC
F9D4
FA9F
FA37
F944
F94C
FA29
FA28
F8F8
F90A
FCBA
02D0
0768
0852
0726
0696
070D
071D
0654
05E0
0671
070C
06A4
05CE
05CD
0684
06BD
064D
0667
0741
06C6
030B
FD5B
F949
F8A8
F9BC
F9E7
F8EA
F86C
F90E
F99A
F92E
F8AE
F931
FA22
FA31
F975
F935
F9AF
F99C
F897
F8B1
FC2F
0223
06D5
07DD
069C
05E3
066C
06D6
066E
0638
06FE
07CE
0763
0630
05BB
064A
06A0
062F
060F
06EB
070D
0429
FEB3
F9FB
F886
F968
FA08
F97E
F8FE
F952
F99B
F901
F84A
F8A2
F9A7
F9F8
F96A
F93D
F9F4
FA50
F970
F8EC
FB54
0099
0583
0749
0692
05FB
0687
06F8
0667
05C6
0640
073B
0745
0653
05CC
064B
06BF
0653
05F1
06A7
074E
0562
0063
FB11
F887
F8EC
F9EA
F9DB
F940
F917
F935
F90A
F8EF
F990
FA70
FA61
F969
F900
F9D9
FA92
F9B9
F881
F9E7
FEDC
048F
0770
070F
05E7
05DE
066F
0661
05DF
05EE
0692
06D2
0663
0624
0689
06C5
0632
05B5
0665
0748
05D3
0126
FBB4
F8C9
F902
FA1F
FA27
F967
F925
F990
F9EC
FA0B
FA54
FA94
FA07
F8CD
F849
F944
FA6C
FA0A
F8D7
F9C7
FE52
0421
0774
0749
05F0
05CA
06BB
0746
06F5
0692
067D
0633
058F
055F
060F
06C0
0691
062B
06B9
0782
05FC
0105
FB0C
F7D4
F867
FA46
FABD
F9C6
F902
F919
F94A
F924
F93F
F9F0
FA79
FA38
F9CE
FA24
FAB0
FA1D
F8D2
F960
FD79
0348
0715
0759
0608
05AB
0671
06DD
0671
0639
06D4
0766
0709
0642
060A
0630
05D4
0539
05A3
06FB
06DD
032C
FD27
F898
F7BF
F92D
FA13
F9A3
F924
F96F
F9D8
F99F
F938
F966
F9E1
F9E0
F98A
F9BC
FA5C
FA2E
F900
F8EB
FC1D
01C5
0671
07C1
06C2
060E
068A
070E
06BB
0649
0695
071E
06E5
0614
05B8
0611
064C
0612
0636
0711
0710
042C
FECD
FA06
F857
F920
F9E4
F974
F8C1
F8E4
F98F
F9E4
F9D2
F9D6
F9DE
F975
F8E7
F921
FA17
FA64
F95A
F8BA
FB19
008A
05F6
084C
0795
0641
0609
0686
06AE
067E
0678
0681
062B
05BE
05F4
06B5
070F
06B4
0697
0743
0749
048D
FF3D
FA4E
F870
F938
FA25
F9C8
F8F0
F8D3
F94E
F98C
F978
F9A5
FA09
F9FC
F981
F975
FA15
FA35
F909
F814
F9FD
FF3F
0504
07FE
07C0
068C
064C
06CF
070F
06E3
06BD
068E
0605
0590
05FB
0702
0748
0649
056D
0618
0731
05E7
0141
FBD0
F8EA
F908
F9D6
F97D
F888
F85A
F900
F975
F962
F968
F9C2
F9D2
F959
F92E
F9DE
FA73
F9C7
F8C7
FA07
FE92
041E
074A
0740
0619
05ED
06A0
0704
06E4
06E2
070A
06BB
0602
05DE
06AD
074C
06B2
05B4
05FD
073B
06C2
02C4
FCFC
F90B
F889
F9C3
FA54
F9CE
F942
F930
F913
F8B0
F897
F901
F941
F8EA
F8B5
F962
FA2F
F9BA
F876
F8F5
FCEC
02A8
0690
0707
05CE
0566
0635
06F4
06FA
06D8
06FD
06F8
0689
065E
070C
07E4
07CC
0706
06F2
07AE
072C
038B
FDDD
F964
F825
F919
F9FC
F9F3
F9AB
F99E
F96E
F8EF
F8AD
F8F2
F916
F88B
F800
F875
F977
F97E
F860
F862
FBBF
0199
0679
07FF
071B
0646
0678
06CE
068A
062D
065D
06D7
0703
06FE
073C
0781
072C
0687
06B7
07C5
07B5
0487
FEF3
FA14
F833
F8B2
F96D
F963
F929
F94D
F96C
F929
F8F9
F950
F9AC
F95A
F8BE
F8E6
F9C5
F9FF
F905
F89A
FB20
0074
0594
07C4
073B
0639
0625
0694
06C2
06CF
071E
0760
0710
0666
061A
0638
0624
05DA
063F
077B
07D5
0541
0015
FB2D
F8FE
F93A
F9C5
F975
F8E9
F8F3
F950
F961
F941
F964
F999
F958
F8EA
F933
FA24
FA59
F90C
F7E5
F99A
FEA5
0442
0744
073F
063F
0602
066B
06A9
06A7
06C6
06EA
06AA
0643
0664
0700
072D
069D
0652
0712
079E
05B0
00E2
FBAF
F8F3
F8FE
F9D5
F9E2
F978
F97E
F9DA
F9D2
F95B
F913
F922
F913
F8E3
F941
FA43
FAAA
F97B
F80E
F940
FE18
0415
0799
079F
0636
05AD
063E
06C5
06BA
068B
0687
0674
0650
068A
0720
073D
0674
05BB
0639
0728
061E
01E3
FC62
F8DD
F889
F9B1
FA29
F9A5
F934
F954
F984
F967
F953
F984
F99E
F962
F94A
F9BC
FA11
F964
F86D
F97B
FDD1
0397
0761
07AD
0628
055D
0609
070A
0753
06F8
067C
0607
05B5
05DE
0681
06DF
0668
05C9
062E
0740
06D6
0351
FDDE
F993
F847
F8FC
F998
F95A
F907
F93D
F9A8
F9C5
F9AA
F99F
F990
F95F
F967
F9F4
FA65
F9C5
F884
F8CD
FC46
01CC
063D
0799
06B6
05CC
05EF
068F
06E6
06ED
06DC
069E
0635
0618
0688
06E5
067F
05CE
060D
0731
072D
0411
FEAA
FA15
F88C
F94F
FA11
F9C0
F917
F8F0
F91B
F916
F90D
F96B
F9F1
F9F7
F986
F957
F99C
F997
F903
F934
FBD8
00A3
0519
0711
06D2
0642
0681
070E
0723
06E3
06D0
06D1
068A
062F
0646
06A1
0678
05C7
05AE
06BE
0765
053C
0013
FACB
F874
F917
FA30
F9E8
F8DA
F884
F8FE
F92F
F8B2
F872
F932
FA4E
FA95
F9DA
F903
F8C4
F921
FA2F
FC82
0045
044E
06DE
0756
06BD
0667
06A2
06F5
0720
0744
0749
06D2
05F4
0568
05AA
064A
0692
0695
06DA
06EB
0524
00AD
FB3D
F7E9
F801
F9BB
FA60
F94D
F824
F854
F959
F9C6
F95F
F933
F9E2
FA96
FA3B
F942
F982
FC42
00C6
04FC
074E
07B5
0733
06BB
06A4
06D1
070B
072A
0713
06B6
0627
05B8
05D1
0673
06C1
055D
01A4
FCB6
F8F5
F807
F954
FAA8
FA72
F92B
F85D
F8B5
F963
F96B
F8FD
F905
F9A8
F9F7
F968
F926
FB24
FFC4
04DD
07A4
0767
0605
05A4
067B
071E
06AD
05EB
060B
06F4
0767
06C0
05ED
062B
071A
06BD
0398
FE90
FA40
F894
F92E
FA30
FA40
F99B
F946
F9A5
FA17
F9E7
F934
F8C9
F90A
F966
F926
F8B7
F9BA
FD5A
029E
06D5
0802
06B4
053F
052B
05ED
0628
05AD
058B
0650
0715
06CC
05F7
0630
07C4
089A
0636
00B2
FB1A
F885
F924
FA99
FACA
F9E0
F964
FA06
FAE0
FACB
F9D6
F90C
F901
F91F
F896
F7D1
F878
FBCE
0104
0586
072F
0636
04CD
04CB
05FE
06D8
0680
05B9
05A5
0647
06B0
0690
06BB
07BE
086D
06AD
01F6
FC78
F936
F920
FA69
FACC
F9ED
F930
F991
FA62
FA59
F95D
F8A5
F91A
FA09
FA00
F8C9
F82C
FA42
FF28
047F
0783
0782
0631
05A1
0632
06B6
0651
05A1
05C8
06C0
0756
06D0
0608
0641
0725
06A4
033C
FE03
F9D8
F890
F95C
FA1D
F9D4
F93F
F956
F9DC
F9E2
F93E
F8DD
F96F
FA43
FA04
F892
F7B9
F9A9
FEA7
046C
07FB
0832
0687
0560
05C5
06D3
0733
06C2
066E
06B5
06F1
0664
0593
05C9
071E
0795
04F9
FF88
FA31
F7D0
F873
F9C8
F9E9
F929
F8EB
F983
F9E7
F959
F88D
F8AB
F99C
FA11
F950
F882
F9B9
FDAC
02C6
0681
07A3
0706
0666
06A1
0731
0736
069E
0630
0674
06FD
06FD
0680
0676
074D
07BE
05BB
00CE
FB2D
F7E5
F7E8
F95F
F9EC
F924
F869
F8B2
F957
F93E
F897
F89B
F9AE
FA88
F9D1
F82F
F815
FB44
00CB
05C4
07F1
0781
0655
05FA
0677
06F4
06FB
06E8
0727
077B
074A
0694
0635
06D2
0798
0697
02BF
FD6C
F970
F86F
F96C
FA28
F9A4
F8D6
F8ED
F99F
F9B4
F8E4
F84D
F8E0
F9DF
F9B8
F84C
F7AA
FA06
FF2F
0474
0727
06FC
05D5
058F
065A
0725
072F
06D0
06C3
0714
0727
06AE
064C
06D1
07DC
07A6
049D
FF52
FA64
F839
F8D6
FA25
FA54
F981
F8F4
F930
F966
F8E4
F846
F8A7
F9DB
FA57
F933
F7D3
F8D9
FD3C
02F0
06C2
0763
0650
05C6
0664
0718
06EF
065B
066A
0737
07B6
071B
0610
05F3
0700
0790
0596
00E6
FBAF
F89A
F86C
F9A7
FA52
F9DF
F92C
F905
F92C
F8F9
F886
F8A0
F980
FA1F
F96A
F805
F847
FBE7
01D3
06C1
0836
06CA
0535
0559
06A4
075D
06F3
066F
06BA
074A
0704
0607
05CC
0717
0858
06E4
01EE
FBD0
F801
F7D1
F987
FA8C
FA05
F915
F8F7
F98A
F9DA
F991
F950
F995
F9E2
F95F
F84F
F85D
FB13
000E
04F3
077B
0769
067A
0659
06FA
071D
0633
0537
056D
069E
0748
0694
0595
05E6
0746
0744
03DF
FE1A
F95B
F810
F96C
FAB3
FA55
F933
F8ED
F9B7
FA5A
FA10
F980
F9A1
FA36
FA0C
F8D1
F813
F9EA
FEA2
040C
075A
0791
0624
0531
0581
0645
0682
0647
0648
06A8
06B5
0605
0561
05F5
0775
07B7
04B8
FF11
F9DD
F7E2
F8F9
FA94
FAA6
F992
F90C
F9B9
FA7D
FA25
F918
F8C5
F9B1
FAAF
FA6B
F962
F9B8
FCF2
0212
0653
07BF
06DC
05BB
05B1
0651
0688
0632
061F
06AE
071A
0686
056D
0544
0679
074B
055D
0078
FB2F
F875
F8C7
FA1D
FA72
F9BF
F951
F9B6
FA17
F99E
F8CA
F8CA
F9C6
FA79
F9CB
F880
F8D1
FC32
019E
0647
080A
0723
05A0
0546
061E
06EA
06D5
064C
063A
06B9
0705
06AA
0651
06C6
076F
065E
0266
FCDF
F8C3
F7DA
F91F
FA32
F9F5
F942
F93C
F9B1
F9A1
F8F3
F8BA
F9A0
FAA5
FA34
F866
F78A
F9ED
FF4D
04D2
07B8
07AD
0691
0627
0685
06B7
065F
0631
06CB
07A5
079A
0677
0581
0603
0776
0792
0489
FF17
FA15
F7E8
F880
F9E0
FA5A
F9E5
F970
F95F
F938
F8A4
F824
F874
F962
F9CF
F924
F874
F9B9
FDBB
02EC
06A5
078B
069B
05CB
0602
0698
06B6
0691
06E7
07A8
07CB
06C2
0591
05C9
075A
0806
058D
003F
FB04
F893
F902
FA30
FA4A
F972
F8E6
F92E
F996
F957
F8B1
F88A
F923
F9AE
F959
F899
F919
FC1F
0111
05A5
07CB
0768
062C
05C0
0648
06BE
0684
0622
065B
06FE
0724
069C
065E
0725
07E5
0676
0208
FC84
F8EB
F86B
F97F
F9F5
F956
F8D4
F945
F9F6
F9C5
F8DB
F88E
F986
FAA1
FA44
F894
F7DE
FA60
FFCF
0552
080D
0799
05F6
0550
060C
0706
0741
06EC
06C0
06DC
06B8
0629
05E3
068B
076A
06A7
0321
FDEE
F9A7
F818
F8C8
F9D1
F9EC
F966
F932
F985
F9BF
F96F
F90B
F942
F9EC
FA10
F944
F8AE
FA3B
FE8D
03E4
077B
0808
06CE
0605
0683
073C
06FC
0611
05CB
0697
0756
06E2
05BA
0579
068E
0724
04E6
FFC9
FA7C
F7E1
F855
F9C0
FA18
F950
F8BB
F916
F9BA
F9BF
F946
F933
F9C8
FA26
F987
F8AD
F994
FD5D
02C2
06F9
083A
073F
062F
063B
06C4
06AF
0612
0600
06DE
07A4
0729
05D8
055D
066E
076C
05D4
0112
FB74
F805
F7BC
F8FB
F9AE
F95E
F90F
F97D
FA24
FA19
F962
F8F7
F96B
FA16
F9E6
F8FF
F913
FBC8
00C6
05A7
080C
07B4
066C
0604
069A
0703
068E
05DC
05E4
068D
06D4
064B
05D4
066B
076A
06B6
02F4
FD6B
F919
F7E7
F8F7
F9F1
F99E
F8D4
F8E3
F9C0
FA32
F9A9
F915
F994
FAB0
FABE
F929
F7D0
F967
FE74
045D
07CE
07DB
066E
05D1
0662
06E9
06A1
062A
0665
0708
06FC
0604
054F
0609
0794
07B3
04BC
FF73
FA8C
F849
F8AC
F9E0
FA3F
F9AB
F91D
F932
F983
F970
F919
F930
F9D0
FA14
F943
F846
F936
FD2B
02A3
06A7
079A
0691
05C7
062A
06D5
06C0
0637
0639
06EB
0756
06CC
0600
062C
0746
0793
0547
007F
FB6B
F875
F848
F992
FA81
FA58
F9AE
F95C
F96E
F956
F8DF
F896
F900
F9B3
F9C6
F93B
F98D
FC47
010B
058A
079D
0740
062C
05D2
0627
066D
0679
06BF
0755
079C
0714
0632
05EA
0675
06CB
057E
020A
FD72
F995
F7E4
F855
F989
FA0B
F991
F8F7
F8FE
F963
F96F
F92A
F94A
F9E9
FA11
F936
F8B8
FADE
0003
057D
081E
077F
0613
0602
06F7
075B
06CF
0660
06A6
06E8
0681
0612
065C
0675
0460
FFBD
FACF
F832
F826
F8E3
F925
F945
F9CD
FA2C
F9AD
F8EA
F914
F9FA
FA1C
F92B
F949
FC94
020E
0642
072D
064E
063C
0741
079A
068C
058D
05EC
06C2
0675
0573
05AA
0739
0748
0361
FD02
F86E
F7F7
F9C3
FAAA
F9F7
F947
F992
F9F7
F9A0
F940
F9C2
FA6D
F9DC
F8A3
F96D
FDC0
0396
074D
079F
0681
0631
06A9
069B
05E6
05AF
0651
06AE
0605
056A
062C
0757
0637
01B0
FC14
F8C8
F8A9
F9B5
F9EF
F97C
F977
F9E2
F9D3
F937
F919
F9DA
FA4F
F980
F8B1
FA63
FF23
0468
072B
070F
062A
0623
0696
0680
060D
061C
0699
0696
0605
0624
076C
0800
0568
FFDC
FAA1
F8A5
F974
FA5A
F9E8
F927
F95C
FA08
F9EF
F936
F922
F9D7
F9E5
F8B0
F839
FB16
00E1
0606
079D
0670
056B
05DF
0695
0655
05CA
0622
06F7
06F7
0639
064D
0787
0792
0413
FE15
F971
F88D
F9F1
FAA5
F9E6
F94D
F9D5
FA6D
F9E7
F8F8
F8FD
F9AA
F975
F86F
F90E
FD29
030D
06ED
0728
05C3
0570
0655
06C1
0621
05B5
064F
06FB
06A8
0613
06A2
07AD
068B
01F5
FC3E
F8FF
F91B
FA39
FA18
F918
F8DC
F99C
FA12
F9B1
F96F
F9F0
FA39
F94A
F861
FA16
FF02
0469
0708
0697
0590
05DF
06F1
0742
06B5
0653
0677
066E
05FD
0608
06F7
0747
04E9
FFFF
FB38
F902
F91E
F993
F95E
F931
F9A8
FA11
F99D
F8E1
F913
FA05
FA2D
F915
F8BE
FB7B
00CF
058E
074F
06D6
0673
06EC
0719
0644
057B
05EC
06FC
072B
066F
0653
0750
074E
03F6
FE0A
F91F
F7C6
F8F4
F9DF
F979
F900
F986
FA51
FA3F
F99A
F96B
F999
F90B
F7FE
F8B6
FCE6
02FE
0759
0824
0701
0678
06E1
06D5
05E4
0559
060B
06EA
06AC
05FD
067A
07B8
06E5
0248
FC08
F834
F83E
F9C5
FA04
F910
F8CE
F9BA
FA59
F9C1
F90E
F97D
FA4C
F9EB
F8EA
FA05
FEA4
0475
07C0
0781
0612
05D7
069E
06E0
065B
062B
06AB
06DA
062C
05B9
0677
0710
04FD
FFE7
FAB0
F86C
F90E
FA11
F9DC
F93A
F960
F9E6
F9AB
F8EB
F8F3
F9ED
FA56
F967
F8F1
FB8A
0106
061C
07E6
06E9
05CE
0600
0694
0671
0608
0648
06E8
06DD
063C
0645
072C
06F5
03A7
FE21
F99F
F849
F928
F9DE
F99A
F953
F9B2
FA03
F998
F911
F94F
F9D0
F954
F837
F8DD
FCF3
02E6
0727
07F1
06CA
0627
068C
06C9
0650
05FD
0671
06E9
0686
05F1
0676
0792
06C2
027C
FC8F
F891
F815
F962
FA00
F97F
F919
F968
F9B7
F981
F95A
F9BE
F9EA
F90B
F82D
F9BA
FE84
042C
0768
0771
065D
0639
06DC
0707
0690
0665
06C4
06D5
063D
060E
0714
07E6
05F5
00D0
FB43
F881
F8CB
F9C0
F995
F8D6
F8CF
F96D
F99E
F938
F92B
F9B9
F9C8
F8BB
F832
FA9D
0005
056A
07D1
074E
064B
065E
06E7
06CA
0644
0643
06BE
06D3
0678
06B2
07B2
07A7
0495
FF17
FA3F
F862
F8DA
F972
F941
F922
F9AF
FA22
F9AD
F8EE
F905
F9B0
F985
F866
F879
FBCC
016F
0612
078B
06D6
0642
068B
06B4
0634
05E9
0685
073B
06EA
060D
0631
0758
0728
0397
FDD3
F961
F85E
F986
FA4B
F9DF
F95C
F988
F9C9
F97C
F923
F970
F9D7
F950
F877
F999
FDE7
036F
06DE
0711
05EC
05A7
0651
0698
062A
0600
068F
06F0
0677
0608
06BD
079E
0621
015E
FBC3
F8AF
F8D8
FA02
FA16
F95E
F942
F9E1
FA1E
F99D
F95D
F9EB
FA39
F942
F841
F9E1
FEDC
048A
0789
074D
0620
05FF
069A
06B4
0643
0630
0689
0669
05BC
05C9
0722
07E8
057E
FFF7
FA97
F864
F910
F9FE
F9B6
F91E
F95E
FA06
FA05
F986
F989
F9FE
F9A7
F85D
F842
FB82
014A
0627
07A4
06B3
05EF
0652
06B8
0630
057E
05BC
0694
06D7
0678
069E
0775
071C
03B5
FE26
F9A8
F861
F94E
FA0A
F9CC
F9A3
FA37
FAA8
FA19
F93C
F936
F9B3
F956
F847
F8E2
FCED
02D2
06E8
077B
0653
05F3
068F
06AC
05DF
0567
0604
06BF
068C
061B
06B3
07A2
065C
01C4
FC2A
F8FF
F911
FA24
FA21
F950
F917
F9A3
F9F3
F9B1
F9A9
FA2E
FA3B
F91D
F849
FA38
FF3A
047F
0702
06B4
05F0
0646
06F1
06B7
05F5
05EF
06A6
06CE
05FF
059F
06AF
078D
0575
002B
FAD0
F876
F8E1
F993
F952
F920
F9DA
FA89
F9FB
F8EE
F911
FA3F
FA6C
F8EC
F83F
FB3C
0129
062C
07A6
06C0
062C
06AA
06EC
0645
05BD
0638
06E4
0695
05DB
063C
0780
072A
0366
FDAA
F96D
F875
F95C
F9D3
F95A
F917
F994
F9F6
F98F
F919
F983
FA38
F9D7
F8AB
F925
FD18
0306
074E
0807
06B9
0602
066F
06AE
0628
05E1
068C
0732
06BD
05EC
0643
074D
0666
01FE
FC13
F84B
F801
F947
F9CF
F985
F99A
FA2B
FA33
F970
F8F3
F95F
F9C9
F933
F894
FA42
FF06
04A2
07E6
07E8
0684
05D9
062A
0674
0647
0627
0666
0690
0656
064C
06F1
073F
0539
0069
FB22
F85D
F89A
F9B6
F9DB
F95C
F961
F9CA
F9A0
F8FD
F91D
FA37
FAAF
F97E
F886
FACC
0067
05BE
079B
06B0
05F6
0699
0724
0678
05A8
0618
071E
0703
05DB
0594
06DC
0765
0495
FF10
FA46
F88E
F906
F97A
F933
F906
F964
F9AF
F981
F981
FA32
FAAD
F9BE
F821
F87E
FC68
021F
062A
070B
0660
065E
0726
0756
0690
060C
068D
070B
0660
0572
0617
07E1
07AF
0368
FD08
F8BC
F844
F990
F9F2
F941
F8FE
F984
F9AE
F90A
F8BB
F970
F9F9
F914
F7FB
F972
FE42
03DE
071F
0778
06C9
0694
069D
0641
05EF
066E
075E
0796
06F0
06A3
075E
07C3
05A3
00B2
FB49
F837
F814
F92E
F9C2
F9AA
F99A
F9A5
F94A
F8AB
F891
F918
F935
F86E
F853
FB23
00BC
05F9
07E9
06F6
05F9
067F
0761
072F
0674
0684
072E
0722
0656
0650
077C
079E
0446
FE55
F98B
F856
F95B
F9D1
F90E
F890
F923
F9C1
F97A
F903
F96A
FA1A
F997
F825
F85B
FC37
023F
06B3
0791
0669
05F6
06D2
0781
070B
0645
0647
06B6
0691
0613
0675
0798
0728
0345
FD62
F922
F850
F93D
F987
F913
F942
FA19
FA1B
F8D8
F80B
F90E
FA7E
FA11
F85E
F8E0
FD80
03BD
0774
078F
0668
062B
068E
066E
05FF
063D
06F8
0700
0632
05FD
0712
07BE
05A5
00C3
FBAD
F8E1
F8A9
F990
FA29
FA05
F97D
F92C
F971
FA0E
FA38
F97C
F8B4
F9A3
FD2F
0225
062A
07C1
0750
064E
05E0
0621
066C
0628
0587
0566
0653
078F
0757
0471
FF8B
FAE8
F882
F889
F99D
FA42
FA01
F96A
F94A
F9DC
FA85
FA63
F95D
F8A8
F9F7
FDE2
030E
0704
082D
070A
0591
0553
062E
06D4
0662
0562
0524
0622
0733
067E
0341
FEA0
FAAC
F8C1
F8B8
F96F
F9D9
F9B2
F96F
F99F
FA40
FAAB
FA41
F958
F953
FB82
FFC5
0456
0725
0784
0683
05CA
0612
06C4
06D5
05FF
0511
051E
0636
0702
05BE
01E5
FCE6
F922
F805
F8F3
FA19
FA2F
F96F
F8FB
F97B
FA6E
FAC3
FA0E
F923
F990
FC56
00F0
057A
0802
0808
06BE
05D9
0609
069D
0698
05E8
0577
0601
070F
0723
04FF
00D1
FC32
F905
F81B
F8BD
F987
F9B1
F984
F99E
FA0D
FA3F
F9C0
F8D4
F875
F9B8
FD0F
01BB
05F6
0805
079B
0638
05B8
0678
0730
06C3
05B1
0569
0678
07BD
0772
04A9
0005
FB50
F869
F812
F951
FA36
F9B3
F8A7
F8B7
FA17
FB18
FA46
F85F
F7B0
F9C4
FE1A
02DF
065C
07CA
077C
0698
0646
06B7
0707
066F
057D
058A
06E9
0819
0730
03B9
FEF7
FAB9
F859
F82F
F95D
FA4A
F9F7
F8FE
F8C9
F9B2
FA6E
F9AE
F819
F7F4
FAC1
FFA6
0459
071D
07A5
06CC
05EC
0604
06D8
072C
065D
0568
05CA
0769
0841
066D
0220
FD58
F9F2
F87E
F894
F96A
F9F8
F984
F898
F8A2
F9FA
FB01
FA1A
F826
F802
FB60
00DE
0577
0766
073D
068E
0653
0693
06E3
06CA
0625
0594
0606
0754
07CD
05BA
014E
FC92
F98F
F8C2
F93A
F9AE
F980
F908
F907
F9BB
FA66
F9FF
F895
F7C5
F956
FD51
01E7
053A
06C7
070B
069E
061C
0630
06E9
0760
06DD
060B
0649
0795
07EE
0558
0043
FB50
F8C0
F89E
F972
F9F8
F9D3
F941
F8CE
F8F9
F98B
F992
F8A2
F7E3
F942
FD5C
0299
067A
07B0
06F6
0612
062C
06FE
0768
06C5
05C3
05D7
0772
08F1
07E8
03BD
FE78
FAB3
F948
F950
F9A0
F9AB
F95D
F8F6
F8F1
F97B
F9E4
F93D
F7DA
F7AB
FA62
FF59
03FA
0659
06C0
0682
0655
0649
067D
06F2
0722
06B9
0664
06FC
07DF
06FF
032D
FDD4
F9D6
F8B9
F97E
FA33
F9F5
F92D
F89E
F8B9
F96B
F9FD
F996
F87C
F873
FB1C
0004
04CD
074B
073E
061B
0585
060E
0717
078E
06FB
0613
061E
075B
0812
060B
012F
FC08
F936
F901
F9CC
FA2A
F9DC
F946
F8DE
F902
F99F
F9E9
F920
F7F9
F89D
FC7C
0231
067E
078A
067E
05AB
05FA
06B2
0704
06D3
0666
0630
06A3
078B
0788
050B
0025
FB07
F82F
F831
F97A
FA29
F9C2
F905
F8D2
F966
FA34
FA30
F8EF
F7C3
F909
FD99
035F
0731
07DA
06D6
0636
0696
0728
0725
0695
0603
0600
06C7
07C3
075B
042C
FEEB
FA50
F881
F8F9
F99C
F947
F89B
F890
F92D
F9C3
F9CA
F939
F887
F8AC
FACE
FF21
0411
0736
0789
0657
05AA
0638
072A
077C
0700
0655
064D
072D
07FF
06EF
02F8
FD59
F8F0
F7C3
F936
FADC
FAE1
F98A
F864
F881
F989
FA34
F97E
F7E5
F792
FA98
0084
062F
0889
0777
0580
04F7
05F9
0715
0737
0697
062F
06AF
07D0
0840
0655
019E
FBF6
F857
F817
F9AA
FA97
FA13
F93E
F932
F9BD
F9EB
F93B
F81B
F7A2
F8FD
FCB0
01D4
0639
07FA
0734
05DC
05A5
0672
070B
06CD
0633
0609
06A3
078B
0782
0538
009C
FB84
F877
F864
F9CC
FA6E
F99A
F887
F87F
F961
FA15
F9E2
F90C
F899
F9D5
FD73
0284
069A
07C7
068F
055D
05E7
0777
081B
071A
05B5
0588
06B0
07B7
06F6
03C5
FEF6
FA87
F86A
F8E9
FA4E
FA8D
F95A
F834
F879
F9C6
FA7C
F9AF
F848
F83F
FAE0
FFA7
048F
076B
0783
061B
054A
05ED
070A
0739
0666
05C6
0646
076B
07B3
05E1
01EE
FD2C
F983
F841
F91D
FA6B
FA9C
F9B5
F900
F948
F9E4
F9BA
F8C7
F841
F964
FC7E
00D1
04F7
077B
07B3
0666
0550
0594
06B1
073E
06B4
0605
0649
073F
0767
056A
0142
FC54
F8AF
F7B8
F909
FAA5
FABE
F967
F852
F8BD
F9F8
FA4F
F93B
F838
F94E
FD16
0234
066F
082B
076C
05D2
054F
0657
0787
0765
0638
05AD
06A7
07F1
0761
0417
FF47
FB05
F8AB
F855
F927
F9E3
F9B8
F8F9
F8BE
F975
FA25
F9AB
F866
F81E
FA40
FE84
033F
06B5
080F
0793
0666
05E1
0681
0761
073C
0621
0596
0694
07F5
0773
03FF
FEC5
FA16
F7BC
F7F9
F988
FA90
FA17
F8D4
F860
F949
FA46
F9C4
F826
F7C4
FA70
FF76
0466
0748
07CA
06DF
05EF
05F4
06C2
073C
06B4
05F5
0659
07D7
0885
067F
0205
FD4A
FA3E
F924
F92C
F996
F9E2
F9B4
F934
F912
F986
F9BE
F8F9
F7F7
F88C
FBAE
0062
049C
06EE
073A
0655
056B
0572
067F
0785
0761
0665
0624
0738
0806
065B
01F3
FCC1
F921
F828
F945
FAD4
FB33
FA04
F88D
F868
F990
FA3A
F91A
F781
F845
FC78
020B
0607
0751
06D6
05F7
059A
0614
06F3
0732
0670
05CA
0698
084B
0862
0516
FF96
FAF6
F911
F932
F9AF
F9C6
F995
F942
F90A
F950
F9D3
F989
F82A
F761
F95F
FE3F
039B
06DF
077E
06C4
061F
0618
0689
070A
0715
0695
0672
0797
0910
0843
03DF
FDD6
F978
F830
F8D5
F9AA
F9F1
F9BD
F94A
F8F0
F901
F938
F8BE
F782
F73D
FA09
FFA0
0513
07B5
0796
069A
0611
061F
0693
072F
076F
0719
06E0
0780
083D
070A
02D8
FD3E
F92C
F811
F8E2
F9CE
FA01
F999
F8EA
F87A
F8CB
F977
F94D
F83A
F837
FB43
00B2
058F
07A2
074E
0676
0649
06A3
06FC
0713
06CE
065A
066A
0763
07FF
0600
0103
FBA9
F8E6
F8F3
F9B8
F9AE
F917
F8D0
F90C
F97E
F9DA
F9C9
F905
F830
F918
FD01
0293
06A4
077C
067A
05EE
066B
06FF
070C
06BE
0651
05FB
063B
071E
0747
04DA
FFCA
FA96
F806
F869
F9B6
FA29
F9CC
F96D
F948
F94B
F98F
F9CA
F95A
F8B4
F9D8
FE12
03C2
07A1
0825
06C3
05C9
05E6
0646
064E
0639
0650
0681
06DB
0753
06C8
03A4
FE3E
F977
F7DB
F8E0
FA0E
FA16
F9A5
F997
F9C9
F9CA
F9AD
F993
F945
F91A
FAA5
FF11
04D1
085C
0803
05D4
04E4
05C7
06D0
06D2
0641
0601
0657
06FD
0732
05B2
01AB
FC4D
F891
F86E
FA7C
FB80
FA51
F8EB
F942
FA70
FA4C
F8BE
F80E
FA1E
FE8B
035B
06AF
07BA
06F5
05C4
0565
05D8
060B
057D
0533
0650
07D7
0710
02B3
FCD0
F8B9
F7B4
F879
F958
F9C9
FA1B
FA89
FAE2
FAB6
F9D2
F8D5
F942
FC62
01A3
0676
087C
07D3
06B1
069C
06F0
0672
0569
0531
062C
070C
061F
02D9
FE38
FA20
F82A
F878
F995
F9D7
F90F
F895
F957
FA67
FA2A
F8EC
F921
FC9B
0219
0674
07CE
06F6
05FD
0617
06EB
0765
06FA
063E
0633
06DB
06A4
03CA
FE8D
F9A5
F7CF
F8FD
FA87
FA4E
F8EE
F85F
F92E
F9FF
F996
F896
F8F5
FBFB
00F1
0590
07C6
075B
05FA
0588
065D
072D
06DA
05FD
0616
073C
0769
049E
FF5F
FA77
F851
F8E7
FA39
FA73
F987
F8CD
F948
FA5A
FA7A
F93E
F869
FA65
FF86
0527
0807
077E
05D8
0584
0685
071D
0662
055E
0591
06E1
0763
0531
0065
FB4B
F87B
F89A
F9F3
FA5A
F96A
F8A5
F956
FABF
FAF3
F97A
F865
FA42
FF38
04AF
07C6
07D7
0685
05CE
0632
06BB
067B
05C7
05C2
06BB
074B
0578
00E7
FBA5
F872
F829
F93C
F9AD
F931
F8F7
F9B7
FAA8
FA78
F91D
F84E
FA0B
FEA1
0415
07AD
0841
070D
0634
068E
0717
069D
0585
055C
069A
0785
05D2
0142
FC18
F8F2
F86E
F913
F939
F8B4
F888
F956
FA64
FA6B
F948
F88F
FA3A
FE9C
03C5
071F
07BB
06DF
0669
06DF
075B
0705
0638
0602
06AD
0711
0585
018E
FCA2
F90B
F7F9
F89C
F93A
F8FF
F8A0
F90F
FA08
FA43
F946
F86E
F9CC
FDF1
0327
06ED
0810
076A
06B8
06E2
0760
0732
0649
05B3
0648
0740
0686
02D7
FD6D
F926
F7CC
F887
F930
F8D0
F856
F8EA
FA27
FA81
F952
F80C
F903
FD13
0290
06AD
07EB
072B
067B
06EB
07B5
078B
066A
05BB
067B
07A9
0703
035B
FE02
F9AD
F815
F8A9
F97F
F960
F8BC
F8B3
F97B
F9FF
F943
F804
F881
FC36
01EE
067F
07C8
069F
05A1
0647
079E
07DD
06BB
05B5
0627
076E
075A
0459
FF2D
FA66
F832
F899
F9C3
F9F0
F924
F8AE
F941
F9F2
F97D
F841
F856
FB71
00D0
05A9
07B5
0725
0614
062C
072A
0794
06B4
0589
05A6
0724
07FA
05D3
0093
FADA
F7AF
F7C9
F94C
FA01
F985
F90F
F981
FA35
F9E8
F89A
F813
FA48
FF45
04B9
07D8
07D6
067B
061C
0717
07C2
06CC
052D
050E
06E7
085B
0689
0139
FB55
F81B
F82B
F97E
F9EB
F933
F8A1
F91D
FA02
FA01
F8EB
F863
FA64
FF0B
041C
06F6
0707
060F
0608
0711
07B4
06FE
05CD
05BA
06F8
07BE
05F6
0166
FC22
F8CF
F863
F98C
FA38
F9A5
F8CD
F8DF
F9AD
F9F7
F935
F8AC
FA48
FE72
0354
067D
071D
0675
063C
06DA
0753
06C2
05A3
055A
0671
0782
064C
0212
FCB7
F923
F893
F9A4
FA22
F96D
F8C1
F94A
FA7C
FAC4
F9A8
F8B3
FA00
FE04
02EF
0648
0719
0685
064A
06E2
0748
068A
0536
04D8
0610
0765
0679
0272
FD0D
F926
F82C
F91F
F9EE
F994
F8D5
F8F9
FA18
FAE5
FA4A
F90D
F971
FCEA
0253
06BB
0821
0737
064E
06B4
078F
0751
05F1
050E
05E2
076D
0722
037F
FDCB
F923
F7A4
F8A8
F9C5
F972
F85E
F836
F960
FA72
FA04
F8B7
F8EB
FC42
01B0
064B
0807
076B
0692
06CC
0785
0771
0670
05C9
0682
07C2
0751
03CE
FE5B
F9C8
F818
F8D5
F9DB
F9A7
F8A7
F84F
F921
FA08
F9BF
F89F
F8B1
FBA7
00E5
05C3
07EC
0767
063C
062B
0707
076C
06B8
05E6
063C
076C
076C
047E
FF3F
FA66
F84D
F8D5
F9D9
F9A6
F8A4
F86D
F988
FAA3
FA3C
F8C3
F88A
FB61
008A
0547
0773
074C
06B6
06FB
079D
075B
060E
050D
059B
071C
0756
04A7
FFC9
FB3D
F8ED
F8A8
F8DD
F88B
F821
F87D
F992
FA52
F9F2
F900
F91A
FB85
FFE9
0460
0701
076C
06E9
06DD
075F
0775
06A5
05CB
0617
0757
07AF
0558
0080
FB51
F82C
F7D3
F91C
FA23
F9F8
F937
F90C
F9A8
F9F8
F92A
F83F
F981
FE0B
041B
0858
08E9
070A
0569
056D
064F
06B1
065F
064B
0703
0791
0625
01FC
FC8E
F898
F7BD
F923
FA83
FA83
F9C9
F9A3
FA18
F9ED
F8AA
F7DF
F9BA
FE79
03C8
06DC
0705
05F1
059D
0653
06C8
0611
0505
0552
0741
08C2
072C
0213
FC1D
F8B7
F8E8
FA9F
FB28
F9FC
F8CE
F92C
FA90
FB0C
F9B7
F80B
F8AA
FCB7
0271
06A5
078B
0635
0524
05A8
06CD
06EF
05E6
053A
061B
079B
0751
03DE
FE7E
FA0C
F882
F965
FA92
FA77
F970
F8EB
F97E
FA2A
F9BF
F8AB
F8ED
FBFF
00FF
0547
06F0
0676
05CF
0627
06E4
06E0
0615
05BE
06B9
0813
0790
03ED
FE75
FA1D
F8D1
F9CD
FAAC
FA0A
F8B6
F85B
F948
FA13
F972
F81F
F868
FBD3
0154
0609
07C5
06E6
05AB
05D3
06FE
078F
06DE
061B
06AD
0812
07EB
046F
FE95
F984
F7B2
F8C6
FA51
FA62
F934
F85B
F8B4
F972
F946
F84A
F85B
FB48
00A1
05C7
0844
07FE
06DD
0684
06D7
06C8
0625
05FD
071F
0897
0833
04A6
FF0C
FA29
F80C
F870
F954
F932
F86D
F872
F9A7
FAB2
FA18
F854
F7C7
FA6C
FFBF
0510
07EC
0814
072F
06D9
072F
0738
066F
05A0
05FD
0767
07F3
0594
006A
FB0D
F842
F870
F998
F9AB
F898
F7EC
F8B1
FA19
FA75
F958
F870
FA08
FEA6
0434
07BF
0815
06AD
05E0
0677
0746
071C
0667
0673
075C
0777
0505
0048
FB89
F907
F90A
F9F1
FA0F
F937
F88C
F8F5
F9EB
FA12
F903
F847
FA13
FED4
0456
07A5
07C0
0640
0567
05EB
06C6
06D6
064E
0646
071B
0789
05B6
0139
FBF4
F8A6
F870
F9D7
FA7A
F99D
F8AF
F92C
FA8B
FAE2
F96B
F7E1
F8F7
FD89
0388
07B6
087C
06FF
05A8
05BF
0689
06A4
05EC
05A8
06B6
07E1
06C6
027D
FCEC
F90E
F81E
F8D5
F94F
F914
F90E
F9DA
FABE
FA72
F8D2
F777
F888
FCC8
02A2
073A
08B1
079E
0637
0607
06AA
06E2
0673
065E
0749
0834
0723
0335
FDC5
F96C
F7CE
F866
F95D
F973
F8F2
F8E8
F98D
F9D1
F8C9
F761
F801
FC1D
024C
0744
08C7
0776
05D4
05BA
06DE
07B2
0762
06AD
06C4
0787
0730
0410
FEAA
F9B5
F7AF
F876
F9AE
F983
F880
F854
F95A
FA1C
F95C
F7F7
F849
FBBF
0144
061D
083D
07C9
069A
066D
0761
0821
0795
0648
05CB
0694
06F2
04B3
FFC7
FAAD
F80E
F827
F8F7
F8C0
F7E4
F7F1
F94A
FA66
F9C2
F813
F809
FB8A
016F
065C
07FF
072D
0681
0736
0820
07C2
0690
063F
072A
075E
04BB
FFA2
FAC3
F85A
F836
F89E
F894
F882
F8EE
F959
F8F3
F81B
F892
FBC6
0102
05B2
07B7
074D
066D
0674
06F3
06EE
069E
0711
081E
07B0
03FF
FE26
F994
F881
F9B6
FA60
F976
F879
F8DD
F9EB
F9E3
F8BB
F8BC
FBEF
017B
063C
07E2
0707
05FC
0612
06A3
0695
061F
0658
0730
06BD
0348
FDBC
F938
F7F1
F911
FA22
F9F7
F97A
F9A5
F9EA
F94A
F877
F9A9
FDEC
0362
06F8
078E
06BD
0684
0706
06FF
0609
0565
0632
076B
067A
0229
FC66
F88F
F80E
F934
F994
F8DA
F899
F99F
FA8F
F9E1
F898
F9A4
FE51
0438
07A4
0789
0634
0627
0747
07BC
06D9
0607
0682
0731
05A2
0118
FBC9
F8B0
F890
F991
F9AD
F8E0
F894
F952
F9E4
F93C
F87C
FA28
FF08
04AF
07D1
07AA
066F
0652
0717
0726
0644
05FE
071A
07CA
057C
0029
FAD0
F85C
F8C0
F99E
F955
F894
F8C7
F9C8
FA09
F901
F88A
FAFF
0047
0571
07A3
06FD
0605
067C
0788
076E
0650
0603
0728
079A
04C4
FF0D
F9E1
F81A
F923
FA2F
F9B2
F8B7
F8C4
F989
F97E
F879
F87D
FB89
00FD
05E5
07D8
0730
062D
0646
06E1
06D1
064A
0683
0788
0763
0432
FEBC
FA11
F868
F8FA
F973
F8F3
F8A6
F96D
FA36
F985
F80F
F887
FC77
0221
0629
0718
067F
0692
077E
07BD
06AB
05B4
0667
07F1
0780
036C
FD75
F93B
F887
F9B2
F9FF
F8E3
F825
F8F5
FA13
F9A4
F835
F8A2
FCB8
02B4
06E9
07A0
0686
0631
0720
07C6
072A
0644
0672
073C
067C
02D3
FD8E
F987
F858
F8FD
F963
F8DE
F876
F8F9
F9AA
F966
F8BA
F9D4
FDE8
034A
06E0
076A
0693
0684
0757
079B
06DD
0667
0729
07D1
05EF
010E
FBB2
F8D9
F8E9
F9B4
F959
F84F
F833
F93E
F9D8
F8EA
F7E8
F995
FEB6
04A5
07DD
079D
0653
0666
0788
07CB
06BC
0619
0722
083B
0661
00EB
FAD8
F7C9
F84D
F9D4
F9F0
F8CB
F818
F880
F8F5
F89A
F87A
FA98
FF65
04B3
07AD
07A4
0672
0631
070B
07B1
077C
0741
07B5
07BB
0551
003F
FAFD
F852
F889
F98C
F99D
F903
F8D7
F909
F892
F779
F7AC
FAFF
00AC
059E
076E
06AB
05D0
0659
0771
0799
06DF
06BC
07A7
07C8
04DB
FF40
FA2E
F86D
F970
FA57
F987
F844
F86F
F9A4
F9D6
F88D
F83A
FB71
0172
068B
0803
06C0
05AC
0630
0726
071B
0679
06B3
07AE
072D
0368
FD9B
F92F
F83D
F989
FA49
F97B
F89E
F920
FA2D
F9EF
F89A
F8E2
FCC3
02B3
0701
07CB
06B4
0656
0711
073E
061C
0533
061D
07C7
0722
02AD
FC88
F869
F7DF
F935
F9DF
F954
F8F1
F989
FA17
F963
F859
F98E
FE23
03F1
077B
0799
065C
063D
0731
0762
0640
0587
06A1
0817
06CD
01CB
FBC5
F855
F846
F95B
F970
F8D5
F91B
FA53
FAB2
F934
F7AD
F936
FE8D
04C8
081D
07B7
0624
0602
071F
0774
065F
0595
067A
079F
060E
010B
FB69
F892
F8E7
F9DF
F97F
F888
F8C1
FA15
FA91
F956
F850
FA3F
FF62
04D7
0790
0753
065C
0667
06ED
069D
05B2
05C8
0749
080A
0569
FFAC
FA41
F844
F949
FA51
F99E
F876
F8C9
FA36
FA8D
F922
F84F
FAD6
0066
0596
0792
06E4
0636
06E0
07AC
0715
05AE
0571
06CF
0784
04F2
FF62
FA1B
F80A
F8DE
F9EF
F99E
F8DA
F91C
FA00
F9E2
F8A3
F898
FBEB
01A0
0639
076A
065F
05D9
06BE
0789
06E8
05C7
05F6
0753
075A
03FB
FE4F
F9BA
F869
F94F
F9E2
F93B
F8AF
F969
FA76
FA07
F860
F84E
FC0F
024B
070F
07F4
0667
057F
0646
0720
06AA
05CE
0642
078E
06FA
02CF
FCE0
F8E3
F888
F9F8
FA6A
F967
F8B5
F972
FA66
F9D9
F877
F926
FD9A
03D1
07D7
07F5
0637
0598
0683
070C
062D
0563
065F
07F4
06D9
01AF
FB35
F79C
F815
FA06
FA81
F97B
F8F3
F9B9
FA58
F983
F881
FA11
FEFD
04B1
07CC
0797
064C
061D
06D8
06E4
05F2
058B
06A2
0795
05A8
006D
FACE
F817
F893
F9C7
F9BE
F911
F94B
FA42
FA3B
F8B4
F7E4
FA7A
0036
05BA
07F9
0730
0614
0669
0759
0736
061B
05D0
0716
07FB
05C3
0041
FA8B
F7E2
F86E
F997
F95C
F871
F8A7
F9F7
FA6F
F91F
F80B
FA2F
FFC5
0593
083E
07AA
067A
06A3
0778
0759
0659
0623
0746
07C3
051A
FF81
FA27
F7F6
F8AA
F99F
F935
F866
F8C8
F9EA
F9E2
F861
F7F1
FB2A
0144
067E
081A
0719
0668
071A
07A2
06B7
0594
063F
0837
0849
043A
FDBE
F8E8
F7EA
F924
F9AF
F8DA
F856
F946
FA66
F9D9
F82E
F863
FC78
02BD
074A
0813
06BD
0636
072D
07DA
06F9
05BB
0606
0766
0707
0306
FD07
F8B8
F7FB
F93F
F9D6
F915
F87F
F929
FA16
F9C2
F8AD
F959
FD62
0330
074A
07EC
06A5
0620
06FB
0797
06D7
05DF
0657
0790
06BB
024D
FC55
F88F
F85C
F99D
F9B4
F8A0
F84E
F970
FA5A
F988
F83A
F970
FE3D
041E
077E
0777
064F
0660
0772
07B3
06A1
05D6
06A0
07AC
062B
0144
FB8C
F871
F8A3
F9CB
F9AC
F8A3
F87B
F985
FA1D
F92F
F849
FA1D
FF29
04B5
0795
0763
0665
0688
0759
074D
0648
05D4
06C8
078D
0596
0087
FB14
F852
F890
F983
F94D
F886
F8CD
FA15
FA91
F96A
F889
FAAF
0003
0570
07DF
075B
0664
06A1
0741
06D4
05B6
059E
06E5
0760
04A6
FF20
FA01
F802
F8C5
F9D2
F9AF
F92B
F98C
FA6A
FA3D
F8EC
F8B5
FBCF
0181
0670
080E
0710
0612
065D
06DE
0657
0571
05C5
0728
0723
03B2
FDFB
F975
F84B
F95C
FA0B
F96C
F8D2
F971
FA72
FA3B
F90F
F965
FD0A
029A
06A5
074E
0614
05A8
06AF
0776
06B8
0588
05B7
06EB
0678
0293
FCE6
F910
F8C4
FA34
FA96
F972
F8A6
F972
FA9F
FA4F
F8F6
F960
FD66
034D
074C
0783
05C4
0513
0625
071E
068D
0581
05DE
0738
06B3
0277
FC6A
F883
F884
FA55
FADD
F9AD
F8DA
F9A3
FAA1
F9FE
F88E
F95A
FDDA
03B8
0729
0704
059A
0585
06A9
0711
0619
0564
0654
0794
0646
018D
FC07
F91B
F966
FA87
FA4C
F920
F8DF
F9EF
FA9E
F9A8
F86D
F9BB
FE68
03F8
0716
06FE
05D7
05D7
06D0
0716
0636
05AF
069F
07A1
05FB
0102
FB6B
F89E
F921
FA70
FA4D
F938
F906
F9DC
F9F2
F886
F7C0
FA6A
0034
057E
0745
064C
058D
064F
0722
06B4
060D
06C3
07E4
0673
014B
FB3A
F826
F8BA
FA2C
FA15
F911
F8F1
F9B2
F9C2
F907
F9C6
FDC0
0363
0730
07A3
067E
0611
0680
069B
0647
0691
074F
065F
0245
FCAD
F8FC
F88E
F992
F9D5
F969
F98D
FA19
F9A5
F860
F8EB
FD33
0361
0767
0793
061D
05CE
0697
06A9
05DC
05FA
0766
077B
03AA
FD58
F8CF
F84E
F9C6
FA1F
F934
F910
FA1D
FA65
F905
F87C
FBC1
01EB
06B3
0777
0613
05D1
0708
077A
065C
05A5
06AB
074D
0464
FE65
F97C
F89E
FA29
FA9D
F945
F86A
F93F
FA04
F924
F875
FB37
014B
068C
079F
05DB
0501
0642
076F
06EC
0625
06E1
07B2
0558
FF78
F9E4
F83B
F9BB
FAD2
F9F6
F8F0
F958
FA03
F93D
F840
FA2F
FFA0
0523
072F
063C
057C
0658
072B
068B
05CA
06AC
07EA
062F
00B8
FB08
F8E7
F9F6
FACD
F9C6
F8A8
F940
FA52
F9AB
F820
F939
FE6D
0497
0771
0694
054E
05E8
0721
06EF
05EF
063E
0795
06D6
0232
FC22
F8C4
F914
FA53
FA1B
F927
F945
FA18
F9C5
F875
F904
FD53
0345
06E2
06EF
05D5
05F5
06C9
06A0
05C3
060C
077C
0746
0347
FD4D
F957
F902
FA23
FA2D
F95B
F95F
FA2C
F9F9
F88A
F885
FC3F
023C
0677
06FC
05CB
05A3
0686
06AB
05E3
0605
0799
0800
0475
FE1E
F94F
F89B
FA28
FAA9
F99C
F916
F9E9
FA48
F8EA
F7E8
FA8D
00BB
065B
07F3
0670
0547
05E8
06B4
064D
05DA
06CF
07D0
05CD
003A
FA79
F826
F91B
FA50
FA09
F96A
F9C8
FA3F
F960
F845
F9E7
FF21
04E4
077E
06C8
05AE
0613
06DA
0674
05A9
0636
0772
0653
0173
FB8A
F88F
F930
FA84
FA33
F91B
F925
FA04
F9DD
F8C6
F986
FDEE
03D9
074F
071C
05C7
05D4
06C5
06C6
05F4
0616
0737
06A6
0269
FC78
F8DC
F8F1
FA31
F9F9
F8DD
F8F7
FA37
FA6C
F910
F8F7
FCC9
02FF
0735
075A
05CF
05C3
0717
0764
061F
056F
0678
06DE
03A4
FDA0
F90E
F887
FA1C
FA6C
F916
F86D
F970
FA46
F987
F91F
FC10
01F1
06BE
0799
060C
0581
06B6
077F
06AB
05DF
06A5
0745
049C
FEB0
F96D
F81C
F9A8
FA96
F9AA
F8C2
F94A
F9F8
F93E
F883
FAD4
0085
0601
07DA
06A9
05A3
0638
06E9
066E
05F6
06E9
07DA
05B5
0011
FA77
F86B
F96E
FA4B
F991
F8DC
F993
FA63
F97A
F815
F99F
FF14
050E
0791
06A2
058A
0636
0735
06BD
05BC
0636
0787
0674
017F
FB7C
F87D
F91A
FA61
FA12
F919
F93A
F9F2
F97F
F852
F95C
FE29
0431
0777
071B
05DB
0611
06FF
06DD
0609
065A
07A4
0702
0287
FC59
F89C
F8AC
FA07
FA03
F901
F8EB
F9C7
F9BF
F886
F8BA
FCAF
02E2
073B
07B2
063E
05C8
0694
06F0
0665
065F
0756
0724
038F
FDB1
F944
F86D
F999
FA0F
F964
F920
F9B8
F9C2
F8AB
F88D
FBD8
01BB
0677
078F
0658
05B5
065D
06CB
0648
0625
0733
0791
049B
FEBC
F9A6
F83D
F987
FA7D
F9FB
F96C
F9D1
FA0C
F910
F86F
FAEE
009F
0604
07DF
06B5
058D
05E2
0673
060D
05AD
069C
078C
0586
FFF9
FA31
F7DE
F8F5
FA61
FA33
F97D
F9C3
FA56
F9AE
F89F
FA18
FF3A
0531
081E
076F
05EF
05D7
0675
0649
05C9
066A
0784
063D
0143
FB3A
F80D
F880
F9DD
F9DA
F92E
F97C
FA47
F9C8
F863
F928
FDEB
043B
07D3
0780
060D
0628
072C
0706
05E0
05DD
0741
0716
02E1
FC75
F850
F856
F9FF
FA1E
F8DD
F88C
F9A0
FA16
F910
F8FD
FC97
02C3
074A
07C5
0628
05B2
06C5
0755
0698
062B
06FB
0701
03A1
FDAD
F90E
F848
F9BA
FA42
F945
F8A4
F942
F9AD
F8E4
F8C2
FBE3
01C0
0695
07B4
0669
05C6
0699
0733
06AB
065C
0747
079C
04A4
FEC2
F9BC
F86C
F99E
FA34
F94F
F8B8
F971
F9F3
F8E9
F81A
FAA6
0098
0619
07C8
0682
05A3
0676
073F
06A3
05F9
06E0
07F2
05F0
0040
FA6B
F82C
F934
FA42
F9A7
F8D9
F95D
FA1E
F952
F801
F972
FECD
04F2
07DE
0732
05F2
0638
06FE
06A8
05ED
0693
07F3
06EC
01F7
FBC0
F859
F8A2
F9E2
F9C9
F90F
F958
FA25
F9A6
F82E
F8C3
FD49
038A
076D
079D
0676
0662
06FC
06B5
05DF
0638
07A0
074B
032D
FD1F
F90E
F889
F980
F993
F8FB
F936
FA0F
F9D1
F870
F895
FC6E
026A
06A7
075B
066E
065B
070F
06EE
05F9
05F9
0759
078F
0417
FE15
F982
F89C
F9AE
F9E8
F90C
F8EA
F9F1
FA52
F91B
F87F
FB66
014F
0655
07A7
0684
05FC
06D4
0749
0670
05D1
06B9
0779
0511
FF6B
FA1B
F858
F96D
FA3F
F97F
F8BB
F947
FA11
F994
F8E6
FAD7
0009
056D
07A3
06CC
05CD
0650
0720
06C6
0608
066E
072F
0584
0074
FAD1
F838
F8F3
FA25
F9CE
F8ED
F92A
F9F6
F9A6
F8BD
FA0D
FEF0
04D1
07D2
0741
05E9
061A
070B
06F4
062E
0678
078C
0691
01D7
FBB5
F843
F8A0
FA1D
FA1E
F928
F924
F9F9
F9D2
F899
F918
FD73
03BE
07B8
07B1
061C
05EC
06F5
072B
0644
061E
074A
073A
035B
FD06
F882
F811
F9A5
FA1A
F933
F8EC
F9C7
F9F9
F8BF
F888
FC20
027A
074E
0807
067F
05F8
06E0
0736
0650
05FD
073A
07BB
047E
FE32
F915
F80D
F98D
FA3A
F957
F8DC
F9BD
FA4B
F938
F873
FB1D
0117
0678
0804
06BB
05E2
069A
072D
0677
05E1
06D3
07AE
0556
FF95
FA19
F843
F95B
FA28
F969
F8CE
F997
FA59
F96E
F849
FA3B
FFE0
05A2
07D4
06E1
0603
06B8
0766
06A9
05CC
0696
07D1
062F
00CA
FAF1
F866
F918
F9F7
F957
F899
F934
FA14
F96E
F82E
F97D
FE8F
047D
0775
070D
0616
067F
0740
06D2
05FB
0686
07DC
06ED
022E
FC26
F8CC
F8FF
FA18
F9D3
F8F2
F92C
FA0A
F9B1
F85B
F8FC
FD76
038C
0726
070F
05D8
0600
06F1
06D3
05E5
0619
0784
0747
0328
FD00
F8ED
F898
F9CA
F9E4
F919
F92A
FA15
FA12
F8C5
F8B6
FC4C
0249
06CE
07B8
06A7
063D
06CB
06D4
0612
0606
0737
0776
043F
FE5A
F985
F849
F95D
F9E8
F943
F903
F9D2
FA2C
F90F
F868
FB1C
00F4
0638
07DB
06C7
0605
069F
0705
064B
05DB
06E3
07A3
052A
FF77
FA20
F843
F929
F9EB
F969
F904
F9AB
FA21
F938
F86A
FA7A
FFBD
0528
079F
0720
0613
061D
06BD
06D5
0666
0634
066D
0687
0647
0619
064C
0693
0685
063D
0626
0653
066E
0645
0617
062B
0662
066C
063B
0610
0613
0625
061C
0604
0602
0616
061E
0609
05F1
05EF
05FF
0605
05F9
05EF
05FD
0617
0623
0611
05ED
05D4
05D7
05E6
05E7
05D4
05C2
05C7
05D7
05CF
05A9
0585
0587
05AA
05C5
05BF
05A8
05A3
05B2
05BC
05B2
05A4
05A6
05B1
05AE
059A
0588
0586
0586
0578
0561
0552
0550
054F
0549
0548
0551
0559
0551
0542
0545
0559
0564
0555
0542
0544
0558
055E
054D
053A
0536
053C
0539
0530
0532
053F
053D
0521
0501
04FA
050B
051A
0516
0508
04FC
04EF
04E0
04D8
04E1
04F4
04FD
04F5
04EB
04EE
04FB
04FC
04ED
04D9
04CF
04CF
04D2
04D3
04D3
04D6
04D6
04CA
04B3
04A0
049E
04AC
04B6
04B0
04A1
0499
049C
049F
0498
048F
0492
049A
0490
0474
045C
045F
0471
047D
047D
047C
047E
0473
0457
043E
0445
0465
047C
0476
0462
0459
045A
0455
044D
0451
0462
046B
045B
043F
042F
0433
0438
0431
0426
0425
0429
0425
0414
0407
040D
0421
042E
0427
0410
0400
03FF
0406
0405
03FC
03FA
0404
0409
03F4
03CD
03B8
03CB
03F1
0402
03F3
03DD
03D7
03D7
03CE
03C6
03D3
03F1
03FC
03E1
03BB
03B1
03C6
03D7
03CE
03BC
03B6
03BA
03B0
0397
0384
0387
0394
039C
039D
03A0
03A7
03A4
0397
038E
0395
03A5
03AE
03AB
03A3
039B
038C
0377
0366
0364
036C
036F
0363
0350
0345
0348
0353
035F
036A
0373
0373
036B
0363
0362
0366
0367
0361
035A
0359
0357
0349
0333
0326
032E
033C
0337
031F
030E
0314
0322
0322
0318
031A
0331
0343
0333
030D
02F3
02F9
0310
031E
031F
031D
0317
0305
02EF
02E7
02F1
02FD
02F8
02EA
02E4
02E8
02E9
02E3
02E6
02F8
0305
02F9
02DE
02D2
02E0
02ED
02E3
02CA
02BD
02C2
02C8
02C0
02B6
02B8
02C4
02C4
02B5
02A9
02B0
02C1
02C5
02B5
02A1
029D
02A9
02B1
02AA
029E
029B
02A2
02A3
0298
028A
028D
029F
02AA
02A0
028E
0289
0295
029B
028F
0280
0281
028C
028B
0272
0259
0255
0261
0266
025C
0257
0264
0275
0272
0259
0243
0247
025C
026B
0271
0276
027E
027C
0265
0246
0236
023A
0240
023A
022D
0225
0222
021C
020F
0207
020F
021F
022A
022C
022F
0234
0232
0224
0216
0218
0224
0226
0214
01FD
01F6
0201
020A
0206
01FC
01FA
01FF
01FF
01F5
01EA
01E6
01EB
01EE
01EE
01F0
01F5
01F8
01F1
01E2
01D8
01DC
01EA
01F6
01F5
01E7
01D7
01CE
01CB
01CA
01C8
01CA
01D2
01D8
01D1
01BC
01A8
01A3
01B0
01C1
01CD
01CF
01C9
01BD
01AE
01A5
01A7
01B3
01BE
01C0
01B7
01A8
0198
0189
0184
018D
01A0
01AC
01A4
0190
0184
0188
0193
0197
0196
0198
019D
019B
018D
017F
017F
0189
018C
0182
0178
017B
0186
0189
0180
0172
0169
0163
015E
015E
0167
0170
016F
0163
015A
015A
015D
0156
014E
0153
0163
016B
0161
0152
0152
015E
0161
0153
0145
0148
0157
015A
0149
0138
0138
0144
0147
013D
0135
013B
0147
0145
0133
0124
0128
0136
013A
012D
011E
011A
011F
0122
0120
0122
012C
0136
0136
012A
0121
0121
0127
012B
012A
0127
0122
011D
011C
0121
0126
0120
0112
0108
010C
0118
011B
0111
0105
00FE
00F9
00F1
00EB
00ED
00F7
00FC
00F7
00ED
00E9
00EB
00F0
00F9
0103
010A
0104
00F2
00E2
00DF
00E6
00EC
00EB
00EA
00EA
00E5
00DA
00CF
00CC
00D3
00DA
00DD
00DC
00DC
00DC
00D7
00CD
00C7
00CA
00D3
00DA
00D9
00CF
00C4
00BD
00BD
00BF
00C0
00C1
00C0
00BC
00B2
00A7
00A2
00A6
00AC
00A9
00A0
009B
009D
00A1
00A0
009B
009B
00A2
00AC
00B2
00B0
00AB
00A3
009B
0096
0097
009B
009D
0099
0092
008B
0085
007F
007B
007E
0086
008C
008B
0086
0080
007E
0080
0084
0089
008B
0088
0082
007D
0078
0074
0071
006F
006F
006F
006C
0067
0065
0066
0067
0067
0068
006A
006C
0069
0062
005D
005B
005B
0059
0058
0058
005A
0059
0055
0051
004F
0050
0051
0052
0053
0052
004E
0048
0043
0040
0040
0041
0042
0043
0041
003D
0039
0039
003D
0040
003F
003E
003D
003D
003B
0038
0036
0036
0036
0033
002E
002C
002D
002E
002E
002B
0029
002A
002C
002E
002E
002B
0025
0020
001D
001C
001C
001C
001A
0019
001A
001C
001D
001E
001E
001E
001D
001B
0018
0018
001A
001B
0016
000E
0008
0009
000A
0008
0002
FFFF
0004
000A
0009
0003
FFFE
0001
0007
0006
FFFE
FFF8
FFFA
FFFE
FFFE
FFF8
FFF3
FFF4
FFF6
FFF6
FFF3
FFF4
FFF8
FFF9
FFF6
FFF2
FFF0
FFF0
FFED
FFE9
FFE9
FFEE
FFF2
FFF1
FFEB
FFE6
FFE5
FFE4
FFE1
FFDF
FFDF
FFE1
FFE0
FFDE
FFDE
FFDF
FFE1
FFDF
FFDC
FFD9
FFDA
FFDB
FFD9
FFD5
FFD1
FFD1
FFD3
FFD5
FFD4
FFD4
FFD4
FFD4
FFD3
FFCF
FFCB
FFCA
FFCB
FFCC
FFCA
FFC6
FFC5
FFC5
FFC4
FFC1
FFBF
FFBF
FFBF
FFBD
FFBA
FFB9
FFBB
FFBB
FFB7
FFB2
FFB1
FFB4
FFB7
FFB7
FFB7
FFBA
FFBC
FFB7
FFAC
FFA3
FFA1
FFA6
FFAA
FFAB
FFAB
FFAA
FFA7
FFA1
FF9C
FF9E
FFA4
FFA8
FFA4
FF9B
FF97
FF9A
FF9F
FFA0
FF9F
FF9D
FF9E
FF9E
FF9A
FF93
FF8D
FF8C
FF8D
FF90
FF92
FF95
FF95
FF91
FF8B
FF87
FF88
FF8D
FF8F
FF8A
FF83
FF7E
FF7E
FF80
FF82
FF83
FF84
FF84
FF80
FF7B
FF79
FF7C
FF80
FF81
FF7F
FF7F
FF80
FF80
FF7C
FF78
FF77
FF79
FF7A
FF77
FF73
FF71
FF6F
FF6D
FF69
FF69
FF6B
FF6F
FF70
FF6D
FF6A
FF68
FF67
FF67
FF69
FF6C
FF6F
FF6D
FF68
FF63
FF63
FF66
FF68
FF67
FF63
FF5E
FF5B
FF5A
FF5B
FF5E
FF63
FF65
FF63
FF5D
FF59
FF58
FF58
FF54
FF50
FF4F
FF53
FF58
FF57
FF50
FF4B
FF4B
FF50
FF53
FF53
FF50
FF4E
FF4B
FF48
FF47
FF4B
FF52
FF56
FF53
FF4C
FF46
FF44
FF43
FF41
FF3E
FF3F
FF43
FF44
FF42
FF3F
FF3F
FF41
FF42
FF3E
FF3B
FF3C
FF3F
FF3F
FF3C
FF39
FF39
FF3A
FF39
FF37
FF36
FF37
FF38
FF35
FF31
FF2E
FF2E
FF2D
FF2B
FF29
FF2A
FF2D
FF2E
FF2D
FF2A
FF29
FF2A
FF2B
FF2A
FF28
FF26
FF25
FF26
FF26
FF27
FF27
FF26
FF24
FF23
FF23
FF24
FF24
FF20
FF1B
FF19
FF1A
FF1E
FF1F
FF1D
FF1B
FF1B
FF1B
FF1A
FF17
FF15
FF15
FF14
FF13
FF13
FF15
FF16
FF15
FF11
FF11
FF14
FF17
FF14
FF0F
FF0C
FF10
FF14
FF12
FF0D
FF0B
FF0D
FF10
FF10
FF0E
FF0D
FF10
FF11
FF0F
FF0B
FF08
FF07
FF06
FF06
FF05
FF04
FF03
FF01
FEFE
FEFB
FEFB
FEFD
FEFE
FEFF
FF00
FF01
FF02
FF02
FF02
FF00
FEFE
FEFC
FEFA
FEF9
FEF9
FEF8
FEF6
FEF5
FEF5
FEF7
FEF9
FEF9
FEF6
FEF5
FEF5
FEF5
FEF3
FEF1
FEF1
FEF2
FEF1
FEEE
FEEC
FEED
FEF0
FEF0
FEED
FEEB
FEEC
FEED
FEEC
FEEC
FEED
FEF0
FEF0
FEEC
FEE9
FEE8
FEE9
FEE9
FEE6
FEE4
FEE5
FEE6
FEE6
FEE3
FEE3
FEE4
FEE7
FEE7
FEE6
FEE5
FEE6
FEE6
FEE4
FEE3
FEE1
FEE0
FEDF
FEDF
FEE0
FEE1
FEE2
FEE1
FEE0
FEDE
FEDD
FEDD
FEDD
FEDC
FEDB
FEDA
FEDA
FED9
FED7
FED6
FED8
FEDB
FEDB
FED7
FED4
FED4
FED6
FED7
FED7
FED7
FED6
FED5
FED2
FED0
FECF
FED2
FED4
FED3
FED1
FED0
FECE
FECB
FEC7
FEC7
FEC9
FECC
FECC
FECC
FECD
FECF
FECE
FECB
FEC9
FECB
FECE
FECF
FECD
FECA
FEC9
FECA
FECA
FEC9
FEC8
FEC7
FEC7
FEC6
FEC4
FEC2
FEC3
FEC6
FEC8
FEC7
FEC3
FEC0
FEC0
FEC2
FEC3
FEC2
FEC2
FEC2
FEC3
FEC1
FEBF
FEBF
FEBF
FEBE
FEBC
FEBC
FEBE
FEC0
FEBF
FEBC
FEBA
FEBA
FEBB
FEBA
FEB8
FEB8
FEB9
FEBA
FEBA
FEBA
FEBA
FEBA
FEB9
FEB9
FEB9
FEBA
FEB9
FEB7
FEB6
FEB7
FEB8
FEB8
FEB7
FEB6
FEB5
FEB5
FEB3
FEB1
FEB1
FEB2
FEB4
FEB5
FEB4
FEB3
FEB1
FEAF
FEAE
FEAE
FEAF
FEB0
FEB1
FEB1
FEAF
FEAE
FEAC
FEAB
FEAC
FEAE
FEB0
FEB0
FEAE
FEAC
FEAB
FEAC
FEAC
FEAD
FEAD
FEAE
FEAE
FEAD
FEAB
FEAA
FEAA
FEAA
FEA9
FEA8
FEA7
FEA8
FEA8
FEA8
FEA7
FEA7
FEA8
FEA9
FEA9
FEA8
FEA7
FEA6
FEA5
FEA5
FEA5
FEA5
FEA4
FEA3
FEA5
FEA6
FEA6
FEA5
FEA3
FEA2
FEA1
FEA1
FEA1
FEA0
FEA0
FEA0
FE9F
FE9F
FE9F
FE9F
FE9F
FE9F
FE9F
FE9F
FEA0
FE9F
FE9F
FE9E
FE9E
FE9E
FE9E
FE9E
FE9E
FE9E
FE9E
FE9D
FE9C
FE9C
FE9B
FE9B
FE9B
FE9B
FE9B
FE9B
FE9A
FE9A
FE9A
FE9A
FE9A
FE9A
FE9A
FE9B
FE9B
FE9A
FE97
FE96
FE97
FE99
FE99
FE98
FE97
FE98
FE98
FE98
FE97
FE96
FE96
FE96
FE95
FE94
FE95
FE97
FE96
FE95
FE95
FE95
FE96
FE94
FE93
FE93
FE94
FE94
FE94
FE94
FE93
FE93
FE92
FE92
FE92
FE93
FE92
FE92
FE92
FE92
FE92
FE90
FE90
FE90
FE91
FE91
FE91
FE91
FE90
FE90
FE90
FE8F
FE8F
FE8F
FE8F
FE8E
FE8E
FE8E
FE8E
FE8D
FE8D
FE8D
FE8E
FE8E
FE8E
FE8D
FE8D
FE8C
FE8C
FE8D
FE8E
FE8D
FE8D
FE8C
FE8C
FE8C
FE8C
FE8B
FE8B
FE8B
FE8B
FE8A
FE8A
FE8A
FE8A
FE8A
FE8A
FE89
FE8A
FE8A
FE8A
FE8A
FE89
FE89
FE89
FE89
FE89
FE88
FE89
FE89
FE8A
FE8A
FE89
FE89
FE89
FE89
FE89
FE88
FE88
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE88
FE87
FE86
FE85
FE86
FE86
FE86
FE86
FE86
FE86
FE85
FE84
FE84
FE85
FE86
FE85
FE85
FE85
FE85
FE84
FE83
FE83
FE84
FE84
FE84
FE83
FE83
FE84
FE84
FE84
FE83
FE84
FE84
FE83
FE82
FE82
FE83
FE83
FE82
FE82
FE81
FE82
FE82
FE82
FE82
FE82
FE82
FE81
FE80
FE81
FE81
FE81
FE81
FE81
FE81
FE81
FE80
FE7F
FE80
FE81
FE80
FE80
FE80
FE80
FE80
FE80
FE80
FE7F
FE7F
FE7F
FE7F
FE7F
FE7E
FE7E
FE7E
FE7F
FE80
FE80
FE7F
FE7E
FE7F
FE7F
FE7F
FE7F
FE7E
FE7E
FE7F
FE7E
FE7E
FE7D
FE7D
FE7D
FE7E
FE7E
FE7F
FE7E
FE7D
FE7D
FE7D
FE7E
FE7E
FE7E
FE7E
FE7F
FE7F
FE7E
FE7E
FE7D
FE7E
FE7E
FE7D
FE7D
FE7C
FE7D
FE7E
FE7E
FE7D
FE7D
FE7D
FE7D
FE7E
FE7F
FE7E
FE7D
FE7C
FE7D
FE7D
FE7D
FE7D
FE7D
FE7C
FE7D
FE7D
FE7D
FE7C
FE7C
FE7C
FE7C
FE7D
FE7C
FE7B
FE7B
FE7B
FE7C
FE7C
FE7B
FE7B
FE7C
FE7C
FE7C
FE7C
FE7C
FE7C
FE7C
FE7C
FE7B
FE7C
FE7C
FE7D
FE7C
FE7C
FE7C
FE7D
FE7E
FE7E
FE7E
FE7D
FE7D
FE7E
FE7E
FE7E
FE7D
FE7D
FE7D
FE7E
FE7E
FE7E
FE7E
FE7D
FE7D
FE7D
FE7E
FE7E
FE7D
FE7D
FE7D
FE7E
FE7E
FE7D
FE7C
FE7C
FE7D
FE7D
FE7C
FE7C
FE7C
FE7D
FE7E
FE7E
FE7D
FE7D
FE7D
FE7C
FE7C
FE7D
FE7D
FE7D
FE7D
FE7D
FE7D
FE7D
FE7D
FE7D
FE7D
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7D
FE7C
FE7C
FE7D
FE7D
FE7C
FE7D
FE7D
FE7E
FE7D
FE7C
FE7C
FE7D
FE7D
FE7D
FE7D
FE7E
FE7E
FE7E
FE7E
FE7D
FE7E
FE7E
FE7E
FE7D
FE7E
FE7E
FE7E
FE7E
FE7D
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7F
FE7F
FE7F
FE7E
FE7F
FE7F
FE7F
FE7E
FE7E
FE7E
FE7E
FE7E
FE7E
FE7F
FE7F
FE7F
FE7E
FE7F
FE80
FE80
FE7F
FE7E
FE7F
FE80
FE80
FE80
FE7F
FE7E
FE7F
FE80
FE80
FE81
FE81
FE82
FE82
FE81
FE80
FE80
FE7F
FE7F
FE80
FE81
FE81
FE80
FE80
FE80
FE80
FE80
FE80
FE81
FE81
FE81
FE81
FE81
FE81
FE81
FE80
FE80
FE81
FE81
FE81
FE81
FE80
FE80
FE80
FE81
FE82
FE81
FE81
FE81
FE81
FE82
FE83
FE82
FE81
FE80
FE81
FE83
FE83
FE82
FE81
FE82
FE82
FE82
FE82
FE82
FE82
FE83
FE83
FE83
FE83
FE83
FE84
FE84
FE84
FE83
FE82
FE82
FE83
FE84
FE85
FE84
FE84
FE84
FE84
FE84
FE84
FE83
FE84
FE85
FE85
FE84
FE84
FE84
FE84
FE85
FE86
FE87
FE86
FE86
FE86
FE86
FE86
FE86
FE86
FE86
FE86
FE86
FE87
FE86
FE86
FE86
FE86
FE86
FE87
FE88
FE88
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE87
FE88
FE88
FE88
FE88
FE88
FE89
FE8A
FE8A
FE89
FE88
FE87
FE88
FE88
FE88
FE87
FE86
FE87
FE89
FE89
FE89
FE89
FE89
FE8A
FE8B
FE8B
FE8A
FE8A
FE8A
FE8A
FE8A
FE8A
FE8A
FE8B
FE8B
FE8C
FE8C
FE8C
FE8C
FE8C
FE8C
FE8C
FE8B
FE8B
FE8C
FE8C
FE8C
FE8C
FE8C
FE8B
FE8C
FE8E
FE8E
FE8E
FE8D
FE8C
FE8C
FE8D
FE8D
FE8D
FE8D
FE8E
FE8E
FE8E
FE8E
FE8E
FE8E
FE8E
FE8E
FE8F
FE8F
FE8E
FE8E
FE8E
FE8E
FE8F
FE8E
FE8E
FE90
FE92
FE93
FE93
FE91
FE91
FE91
FE91
FE91
FE91
FE91
FE91
FE92
FE91
FE90
FE90
FE91
FE92
FE93
FE92
FE92
FE91
FE92
FE92
FE93
FE92
FE92
FE92
FE93
FE94
FE94
FE94
FE94
FE94
FE94
FE95
FE95
FE95
FE95
FE94
FE94
FE95
FE95
FE95
FE94
FE95
FE95
FE96
FE96
FE97
FE97
FE97
FE97
FE97
FE97
FE98
FE98
FE97
FE97
FE98
FE98
FE99
FE99
FE98
FE98
FE99
FE99
FE99
FE99
FE98
FE98
FE99
FE99
FE99
FE99
FE99
FE99
FE9A
FE9B
FE9B
FE9A
FE9A
FE9A
FE9B
FE9B
FE9B
FE9B
FE9B
FE9C
FE9C
FE9C
FE9C
FE9C
FE9C
FE9C
FE9C
FE9C
FE9C
FE9C
FE9D
FE9D
FE9D
FE9D
FE9D
FE9D
FE9D
FE9E
FE9F
FE9F
FE9F
FE9F
FE9F
FEA0
FEA0
FEA1
FEA0
FEA0
FEA0
FEA1
FEA1
FEA1
FEA0
FEA0
FEA1
FEA1
FEA1
FEA1
FEA1
FEA2
FEA2
FEA2
FEA2
FEA2
FEA1
FEA2
FEA2
FEA3
FEA3
FEA3
FEA4
FEA4
FEA4
FEA4
FEA4
FEA4
FEA4
FEA4
FEA4
FEA5
FEA5
FEA5
FEA5
FEA4
FEA4
FEA4
FEA4
FEA4
FEA4
FEA5
FEA5
FEA6
FEA6
FEA5
FEA5
FEA5
FEA5
FEA6
FEA7
FEA7
FEA7
FEA7
FEA7
FEA8
FEA7
FEA7
FEA6
FEA6
FEA7
FEA7
FEA8
FEA9
FEA9
FEA8
FEA8
FEA8
FEA9
FEAA
FEAA
FEAA
FEAB
FEAB
FEAB
FEAA
FEAA
FEAB
FEAC
FEAD
FEAC
FEAC
FEAC
FEAD
FEAD
FEAC
FEAD
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAE
FEAF
FEB0
FEB0
FEB0
FEAF
FEB0
FEB0
FEB1
FEB1
FEB1
FEB2
FEB1
FEB1
FEB0
FEB0
FEB1
FEB1
FEB2
FEB2
FEB2
FEB2
FEB3
FEB3
FEB3
FEB3
FEB3
FEB3
FEB3
FEB3
FEB3
FEB4
FEB5
FEB6
FEB6
FEB5
FEB5
FEB5
FEB5
FEB5
FEB5
FEB5
FEB5
FEB5
FEB6
FEB6
FEB6
FEB7
FEB7
FEB7
FEB7
FEB7
FEB7
FEB7
FEB8
FEB9
FEB9
FEB9
FEBA
FEBA
FEB9
FEB9
FEB9
FEB9
FEBA
FEBA
FEBA
FEBA
FEBB
FEBB
FEBC
FEBC
FEBC
FEBC
FEBC
FEBB
FEBC
FEBD
FEBE
FEBE
FEBD
FEBD
FEBE
FEBE
FEBD
FEBD
FEBD
FEBE
FEBF
FEBE
FEBE
FEBF
FEC0
FEC0
FEBF
FEBF
FEC0
FEC0
FEC0
FEC0
FEC0
FEC1
FEC1
FEC0
FEC0
FEC1
FEC2
FEC2
FEC2
FEC2
FEC2
FEC3
FEC3
FEC2
FEC2
FEC3
FEC3
FEC4
FEC4
FEC4
FEC4
FEC4
FEC4
FEC5
FEC5
FEC5
FEC5
FEC5
FEC5
FEC5
FEC5
FEC6
FEC7
FEC7
FEC7
FEC7
FEC7
FEC7
FEC8
FEC8
FEC9
FECA
FECA
FEC9
FEC8
FEC8
FECA
FECB
FECA
FEC9
FECA
FECB
FECC
FECB
FECA
FECA
FECB
FECB
FECC
FECC
FECC
FECC
FECC
FECD
FECE
FECE
FECD
FECD
FECD
FECE
FED0
FED1
FED0
FED0
FECF
FECF
FECF
FECF
FED0
FED0
FED0
FED0
FED0
FED1
FED2
FED1
FED0
FED0
FED1
FED2
FED3
FED2
FED2
FED3
FED3
FED3
FED3
FED3
FED3
FED4
FED5
FED5
FED5
FED5
FED5
FED4
FED5
FED5
FED6
FED6
FED6
FED6
FED7
FED7
FED8
FED7
FED7
FED8
FED8
FED9
FED8
FED7
FED7
FED8
FED9
FED9
FEDA
FEDA
FEDA
FEDA
FEDB
FEDB
FEDA
FED9
FED9
FEDA
FEDC
FEDC
FEDB
FEDB
FEDC
FEDC
FEDD
FEDD
FEDD
FEDD
FEDD
FEDD
FEDD
FEDD
FEDD
FEDE
FEDF
FEDF
FEE0
FEDF
FEDE
FEDE
FEDF
FEE1
FEE1
FEE0
FEE0
FEE0
FEE0
FEE1
FEE1
FEE1
FEE1
FEE1
FEE2
FEE2
FEE3
FEE2
FEE2
FEE2
FEE3
FEE4
FEE4
FEE4
FEE4
FEE4
FEE4
FEE5
FEE4
FEE4
FEE4
FEE5
FEE5
FEE5
FEE5
FEE6
FEE6
FEE7
FEE6
FEE6
FEE7
FEE8
FEE8
FEE8
FEE7
FEE7
FEE8
FEE8
FEE8
FEE7
FEE8
FEE9
FEEA
FEE9
FEE8
FEE8
FEE9
FEEA
FEEA
FEEA
FEEA
FEEB
FEEB
FEEB
FEEB
FEEB
FEEB
FEEC
FEEC
FEEC
FEEC
FEED
FEEE
FEEE
FEED
FEED
FEED
FEEE
FEF0
FEF0
FEEF
FEEE
FEEF
FEF0
FEF0
FEEF
FEEF
FEEF
FEF0
FEF0
FEF0
FEF0
FEF0
FEF1
FEF1
FEF1
FEF1
FEF2
FEF3
FEF3
FEF3
FEF3
FEF3
FEF3
FEF4
FEF4
FEF5
FEF4
FEF4
FEF3
FEF4
FEF5
FEF6
FEF5
FEF5
FEF5
FEF6
FEF7
FEF7
FEF6
FEF6
FEF7
FEF7
FEF8
FEF7
FEF6
FEF6
FEF7
FEF8
FEF9
FEF9
FEF9
FEF9
FEFA
FEFA
FEFA
FEFA
FEFA
FEFB
FEFB
FEFC
FEFC
FEFB
FEFB
FEFB
FEFC
FEFC
FEFC
FEFB
FEFB
FEFD
FEFE
FEFD
FEFC
FEFC
FEFD
FEFE
FEFF
FEFE
FEFE
FEFF
FF01
FF02
FF02
FF01
FF01
FF01
FF02
FF02
FF02
FF02
FF02
FF02
FF02
FF02
FF03
FF03
FF03
FF04
FF04
FF04
FF05
FF05
FF06
FF06
FF06
FF06
FF06
FF06
FF05
FF06
FF06
FF07
FF07
FF07
FF07
FF07
FF07
FF07
FF07
FF07
FF08
FF08
FF08
FF08
FF08
FF09
FF09
FF09
FF09
FF0A
FF0A
FF0B
FF0B
FF0B
FF0B
FF0B
FF0C
FF0C
FF0B
FF0B
FF0C
FF0D
FF0D
FF0D
FF0D
FF0D
FF0D
FF0D
FF0D
FF0D
FF0E
FF0E
FF0E
FF0E
FF0F
FF10
FF10
FF10
FF0F
FF0F
FF10
FF11
FF11
FF11
FF11
FF11
FF11
FF12
FF13
FF13
FF12
FF11
FF11
FF12
FF13
FF13
FF13
FF13
FF14
FF14
FF14
FF14
FF15
FF15
FF15
FF14
FF14
FF15
FF16
FF16
FF15
FF15
FF16
FF18
FF18
FF17
FF16
FF17
FF18
FF18
FF18
FF17
FF18
FF19
FF19
FF19
FF19
FF1A
FF1A
FF1A
FF1A
FF1A
FF1B
FF1B
FF1C
FF1C
FF1C
FF1C
FF1C
FF1C
FF1D
FF1E
FF1E
FF1E
FF1D
FF1D
FF1D
FF1E
FF1E
FF1E
FF1E
FF1F
FF20
FF20
FF1F
FF1F
FF1F
FF1F
FF1F
FF20
FF20
FF21
FF21
FF20
FF20
FF21
FF21
FF22
FF22
FF22
FF22
FF22
FF22
FF22
FF22
FF23
FF23
FF24
FF24
FF24
FF24
FF24
FF24
FF25
FF25
FF25
FF24
FF25
FF26
FF26
FF26
FF26
FF26
FF26
FF26
FF27
FF27
FF26
FF26
FF27
FF27
FF28
FF28
FF28
FF27
FF27
FF28
FF29
FF29
FF29
FF2A
FF2A
FF2B
FF2B
FF2B
FF2B
FF2C
FF2B
FF2B
FF2B
FF2C
FF2D
FF2D
FF2D
FF2D
FF2C
FF2D
FF2D
FF2D
FF2D
FF2E
FF2E
FF2F
FF2F
FF2F
FF2F
FF2F
FF2F
FF2F
FF30
FF30
FF30
FF30
FF31
FF31
FF31
FF31
FF31
FF31
FF31
FF31
FF32
FF32
FF32
FF32
FF32
FF31
FF31
FF31
FF32
FF32
FF33
FF32
FF32
FF32
FF33
FF35
FF36
FF36
FF36
FF36
FF36
FF36
FF36
FF37
FF37
FF37
FF37
FF37
FF37
FF38
FF38
FF38
FF37
FF38
FF38
FF39
FF39
FF39
FF3A
FF3A
FF3A
FF3A
FF3A
FF3A
FF3B
FF3B
FF3B
FF3B
FF3C
FF3D
FF3C
FF3C
FF3C
FF3D
FF3D
FF3E
FF3D
FF3D
FF3D
FF3D
FF3D
FF3D
FF3E
FF3F
FF3F
FF3F
FF3F
FF3F
FF3F
FF3F
FF3F
FF40
FF40
FF40
FF40
FF41
FF43
FF44
FF44
FF42
FF41
FF41
FF42
FF42
FF42
FF42
FF42
FF43
FF43
FF43
FF44
FF44
FF44
FF44
FF45
FF45
FF45
FF44
FF44
FF45
FF46
FF46
FF46
FF46
FF47
FF47
FF47
FF47
FF47
FF47
FF48
FF47
FF47
FF47
FF48
FF48
FF48
FF48
FF49
FF4A
FF4A
FF4A
FF4B
FF4B
FF4B
FF4A
FF4A
FF4A
FF4B
FF4C
FF4C
FF4B
FF4A
FF4B
FF4C
FF4C
FF4C
FF4C
FF4D
FF4D
FF4D
FF4E
FF4E
FF4F
FF4F
FF4F
FF4F
FF4F
FF4F
FF4F
FF4F
FF4F
FF50
FF50
FF50
FF4F
FF4F
FF50
FF51
FF52
FF52
FF51
FF51
FF52
FF52
FF52
FF53
FF53
FF53
FF53
FF53
FF54
FF55
FF55
FF56
FF55
FF54
FF54
FF53
FF54
FF55
FF56
FF57
FF57
FF56
FF56
FF56
FF56
FF57
FF57
FF56
FF57
FF57
FF58
FF58
FF58
FF58
FF58
FF59
FF58
FF58
FF58
FF5A
FF5A
FF5A
FF59
FF59
FF5B
FF5C
FF5B
FF5B
FF5B
FF5C
FF5D
FF5C
FF5C
FF5C
FF5D
FF5D
FF5E
FF5D
FF5E
FF5E
FF5E
FF5E
FF5D
FF5E
FF5F
FF5E
FF5E
FF5D
FF5D
FF5D
FF5E
FF5E
FF5E
FF5E
FF5E
FF5D
FF5E
FF5E
FF5F
FF5F
FF5F
FF5F
FF60
FF61
FF61
FF60
FF60
FF60
FF61
FF61
FF62
FF62
FF61
FF61
FF62
FF62
FF63
FF64
FF63
FF63
FF64
FF64
FF65
FF65
FF65
FF65
FF65
FF65
FF65
FF65
FF66
FF66
FF66
FF66
FF67
FF67
FF67
FF67
FF68
FF69
FF69
FF69
FF68
FF68
FF68
FF69
FF69
FF69
FF69
FF69
FF69
FF69
FF69
FF6A
FF6B
FF6B
FF6C
FF6C
FF6C
FF6C
FF6C
FF6C
FF6C
FF6C
FF6C
FF6C
FF6C
FF6D
FF6C
FF6C
FF6C
FF6D
FF6E
FF6E
FF6E
FF6E
FF6E
FF6F
FF6F
FF6F
FF6F
FF70
FF70
FF70
FF70
FF70
FF71
FF71
FF70
FF70
FF70
FF71
FF71
FF72
FF71
FF72
FF72
FF72
FF73
FF73
FF73
FF74
FF74
FF74
FF75
FF75
FF75
FF75
FF75
FF75
FF76
FF76
FF76
FF76
FF76
FF77
FF77
FF77
FF77
FF77
FF78
FF78
FF78
FF78
FF78
FF79
FF7A
FF7A
FF79
FF78
FF78
FF79
FF7A
FF7A
FF7A
FF7A
FF7B
FF7B
FF7B
FF7A
FF7A
FF7B
FF7C
FF7C
FF7C
FF7C
FF7C
FF7C
FF7C
FF7C
FF7C
FF7D
FF7D
FF7D
FF7D
FF7D
FF7D
FF7D
FF7E
FF7E
FF7F
FF7F
FF7E
FF7E
FF7F
FF80
FF80
FF80
FF7F
FF7F
FF7F
FF7F
FF80
FF81
FF81
FF81
FF81
FF81
FF81
FF82
FF83
FF82
FF83
FF83
FF84
FF85
FF84
FF83
FF83
FF83
FF84
FF85
FF85
FF84
FF84
FF85
FF86
FF86
FF86
FF85
FF86
FF87
FF88
FF88
FF87
FF87
FF87
FF88
FF88
FF88
FF88
FF88
FF88
FF88
FF88
FF88
FF88
FF89
FF89
FF89
FF8A
FF8A
FF8B
FF8B
FF8B
FF8B
FF8A
FF8B
FF8C
FF8C
FF8D
FF8C
FF8C
FF8C
FF8C
FF8D
FF8D
FF8D
FF8E
FF8E
FF8D
FF8D
FF8D
FF8D
FF8D
FF8D
FF8C
FF8D
FF8D
FF8E
FF8E
FF8F
FF8F
FF8F
FF8E
FF8E
FF8F
FF8F
FF90
FF90
FF90
FF90
FF91
FF91
FF91
FF91
FF91
FF91
FF92
FF92
FF93
FF93
FF92
FF91
FF92
FF93
FF93
FF93
FF92
FF93
FF94
FF95
FF94
FF94
FF94
FF95
FF95
FF95
FF95
FF94
FF94
FF95
FF96
FF97
FF98
FF98
FF97
FF97
FF97
FF97
FF97
FF97
FF97
FF98
FF99
FF99
FF99
FF99
FF99
FF99
FF99
FF99
FF99
FF9A
FF9B
FF9B
FF9A
FF9A
FF9A
FF9A
FF9A
FF9B
FF9B
FF9C
FF9C
FF9C
FF9C
FF9B
FF9B
FF9C
FF9D
FF9D
FF9D
FF9C
FF9C
FF9C
FF9D
FF9E
FF9E
FF9E
FF9E
FF9E
FF9F
FF9F
FF9F
FF9F
FF9E
FF9E
FF9F
FF9F
FF9F
FF9F
FF9F
FFA0
FFA1
FFA2
FFA2
FFA1
FFA1
FFA1
FFA2
FFA2
FFA1
FFA1
FFA1
FFA1
FFA2
FFA3
FFA3
FFA3
FFA2
FFA3
FFA3
FFA4
FFA4
FFA4
FFA4
FFA4
FFA4
FFA3
FFA3
FFA4
FFA5
FFA6
FFA5
FFA4
FFA5
FFA6
FFA7
FFA7
FFA6
FFA7
FFA7
FFA8
FFA7
FFA7
FFA7
FFA7
FFA7
FFA7
FFA8
FFA8
FFA9
FFA8
FFA8
FFA8
FFA9
FFA9
FFA9
FFA8
FFA8
FFA9
FFA9
FFA9
FFAA
FFAA
FFAA
FFAA
FFAA
FFAB
FFAB
FFAB
FFAB
FFAA
FFAA
FFAB
FFAB
FFAC
FFAC
FFAC
FFAC
FFAC
FFAD
FFAE
FFAE
FFAD
FFAD
FFAE
FFAE
FFAE
FFAE
FFAD
FFAE
FFAE
FFAE
FFAE
FFAE
FFAF
FFAF
FFAF
FFAF
FFAF
FFAF
FFB0
FFB0
FFB0
FFB0
FFB0
FFB1
FFB1
FFB2
FFB2
FFB2
FFB2
FFB2
FFB2
FFB3
FFB3
FFB4
FFB5
FFB5
FFB4
FFB4
FFB4
FFB5
FFB5
FFB5
FFB5
FFB4
FFB4
FFB5
FFB6
FFB6
FFB7
FFB7
FFB6
FFB6
FFB6
FFB7
FFB7
FFB8
FFB8
FFB9
FFB8
FFB7
FFB7
FFB7
FFB8
FFB9
FFB9
FFB9
FFB9
FFB9
FFBA
FFBA
FFBA
FFB9
FFB9
FFB9
FFBA
FFBA
FFBB
FFBA
FFBA
FFBB
FFBB
FFBB
FFBA
FFBA
FFBA
FFBB
FFBC
FFBC
FFBC
FFBC
FFBC
FFBC
FFBC
FFBC
FFBC
FFBD
FFBD
FFBD
FFBD
FFBE
FFBE
FFBD
FFBC
FFBC
FFBD
FFBE
FFBE
FFBE
FFBE
FFBE
FFBE
FFBE
FFBF
FFC0
FFC0
FFC0
FFC0
FFC1
FFC2
FFC2
FFC1
FFC0
FFC0
FFC0
FFC0
FFC0
FFC0
FFC1
FFC1
FFC1
FFC0
FFC1
FFC2
FFC3
FFC3
FFC2
FFC2
FFC2
FFC3
FFC3
FFC3
FFC3
FFC3
FFC4
FFC4
FFC3
FFC3
FFC3
FFC4
FFC4
FFC4
FFC3
FFC3
FFC4
FFC5
FFC5
FFC5
FFC4
FFC4
FFC5
FFC6
FFC6
FFC6
FFC6
FFC7
FFC7
FFC7
FFC7
FFC7
FFC7
FFC7
FFC7
FFC7
FFC7
FFC7
FFC8
FFC8
FFC8
FFC9
FFC9
FFC8
FFC8
FFC8
FFC8
FFC9
FFC9
FFC9
FFC9
FFC9
FFC9
FFC9
FFC9
FFCA
FFCA
FFCB
FFCB
FFCB
FFCB
FFCA
FFCA
FFCA
FFCC
FFCD
FFCC
FFCC
FFCC
FFCC
FFCC
FFCB
FFCB
FFCB
FFCD
FFCD
FFCD
FFCD
FFCD
FFCD
FFCD
FFCD
FFCD
FFCE
FFCE
FFCE
FFCE
FFCF
FFCF
FFCF
FFCE
FFCE
FFCF
FFD0
FFD0
FFCF
FFCE
FFCF
FFD0
FFD0
FFCF
FFCF
FFD1
FFD1
FFD0
FFCF
FFCF
FFD0
FFD1
FFD0
FFCF
FFCF
FFD0
FFD1
FFD2
FFD1
FFD1
FFD2
FFD3
FFD3
FFD2
FFD2
FFD3
FFD4
FFD4
FFD3
FFD3
FFD2
FFD2
FFD2
FFD3
FFD4
FFD4
FFD4
FFD4
FFD4
FFD4
FFD4
FFD4
FFD5
FFD5
FFD5
FFD5
FFD5
FFD6
FFD7
FFD6
FFD6
FFD6
FFD7
FFD7
FFD5
FFD4
FFD4
FFD5
FFD5
FFD5
FFD5
FFD6
FFD7
FFD8
FFD7
FFD7
FFD7
FFD8
FFD8
FFD8
FFD8
FFD8
FFD9
FFD9
FFD9
FFD9
FFDA
FFDA
FFD9
FFD9
FFD9
FFD9
FFD9
FFDA
FFDB
FFDB
FFDA
FFD9
FFD9
FFDB
FFDC
FFDD
FFDC
FFDB
FFDB
FFDB
FFDB
FFDC
FFDD
FFDD
FFDD
FFDC
FFDC
FFDD
FFDD
FFDD
FFDD
FFDD
FFDE
FFDE
FFDE
FFDE
FFDE
FFDF
FFDF
FFDF
FFDF
FFDF
FFDF
FFDF
FFDF
FFE0
FFE2
FFE4
FFE3
FFE1
FFE0
FFDF
FFE0
FFE1
FFE1
FFE1
FFE1
FFE1
FFE0
FFE0
FFE0
FFE1
FFE2
FFE2
FFE2
FFE1
FFE2
FFE2
FFE3
FFE3
FFE2
FFE2
FFE2
FFE2
FFE3
FFE3
FFE2
FFE3
FFE3
FFE3
FFE3
FFE3
FFE4
FFE5
FFE4
FFE3
FFE4
FFE5
FFE5
FFE5
FFE5
FFE5
FFE6
FFE5
FFE4
FFE4
FFE5
FFE6
FFE6
FFE5
FFE5
FFE5
FFE6
FFE7
FFE6
FFE6
FFE6
FFE7
FFE7
FFE7
FFE7
FFE7
FFE7
FFE7
FFE7
FFE7
FFE7
FFE7
FFE8
FFE8
FFE9
FFE9
FFE9
FFE9
FFE9
FFEA
FFEA
FFE9
FFE9
FFE9
FFE9
FFEA
FFEA
FFEB
FFEB
FFEB
FFEA
FFEA
FFEA
FFEB
FFEB
FFEB
FFEB
FFEB
FFEC
FFED
FFEC
FFEB
FFEB
FFEB
FFEB
FFEC
FFEC
FFED
FFED
FFED
FFED
FFED
FFED
FFED
FFED
FFED
FFED
FFEE
FFEF
FFEE
FFED
FFED
FFEE
FFEF
FFEF
FFEE
FFEE
FFEE
FFEE
FFEE
FFEF
FFEF
FFEF
FFF0
FFEF
FFEF
FFEF
FFF0
FFF1
FFF0
FFEF
FFEF
FFF0
FFF1
FFF0
FFF0
FFF0
FFF1
FFF2
FFF2
FFF1
FFF1
FFF1
FFF2
FFF1
FFF0
FFF0
FFF0
FFF0
FFF0
FFF0
FFF1
FFF1
FFF2
FFF1
FFF1
FFF1
FFF1
FFF1
FFF2
FFF2
FFF3
FFF3
FFF2
FFF2
FFF2
FFF3
FFF3
FFF3
FFF2
FFF3
FFF3
FFF3
FFF3
FFF3
FFF3
FFF3
FFF3
FFF4
FFF4
FFF4
FFF4
FFF4
FFF4
FFF5
FFF5
FFF4
FFF4
FFF5
FFF6
FFF6
FFF6
FFF6
FFF6
FFF7
FFF7
FFF6
FFF6
FFF7
FFF7
FFF7
FFF7
FFF7
FFF7
FFF8
FFF8
FFF8
FFF8
FFF8
FFF8
FFF8
FFF7
FFF8
FFF8
FFF8
FFF8
FFF8
FFF9
FFF9
FFF8
FFF8
FFF8
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0002
0002
0002
0001
0002
0002
0002
0002
0001
0002
0002
0002
0001
0001
0001
0002
0002
0002
0002
0003
0003
0002
0002
0003
0004
0005
0004
0003
0003
0003
0004
0004
0004
0004
0005
0005
0005
0004
0004
0004
0004
0005
0006
0007
0007
0006
0006
0006
0007
0008
0007
0007
0006
0007
0008
0008
0008
0008
0007
0007
0007
0007
0008
0008
0008
0008
0008
0008
0009
000A
0009
0009
0009
0009
0009
0008
0008
0009
000A
000A
0009
0009
0009
000A
000A
000A
000A
000A
000A
000A
000A
000A
000B
000B
000B
000B
000B
000B
000B
000A
000A
000B
000B
000B
000B
000A
000B
000B
000C
000C
000C
000C
000C
000C
000C
000C
000D
000D
000C
000C
000C
000D
000E
000E
000D
000C
000D
000E
000E
000E
000E
000E
000F
000E
000E
000E
000E
000E
000E
000E
000E
000F
000F
000F
000F
000E
000E
000F
000F
0010
0010
000F
000F
0010
0010
000F
000F
000F
0010
0010
0010
0010
0010
0011
0010
0010
0010
0012
0012
0012
0011
0011
0012
0012
0012
0011
0011
0012
0012
0011
0011
0011
0012
0013
0013
0013
0012
0012
0012
0013
0014
0014
0013
0012
0012
0013
0014
0014
0013
0013
0014
0014
0014
0014
0014
0015
0015
0015
0015
0015
0015
0015
0015
0015
0015
0015
0015
0014
0014
0014
0015
0015
0015
0015
0016
0016
0016
0015
0016
0016
0017
0016
0016
0016
0016
0016
0016
0016
0016
0017
0017
0017
0016
0016
0016
0016
0016
0016
0017
0018
0018
0018
0017
0016
0017
0017
0018
0018
0017
0017
0017
0018
0018
0019
0018
0018
0019
0019
0019
0019
0019
001A
0019
0019
0018
0018
0019
0019
001A
001A
001A
0019
0019
0019
001A
001A
001A
0019
0019
001A
001B
001A
001A
0019
001A
001B
001B
001B
001B
001B
001B
001B
001B
001B
001B
001B
001B
001B
001C
001D
001D
001D
001C
001C
001C
001C
001D
001D
001C
001C
001C
001D
001E
001E
001D
001D
001D
001E
001F
001F
001F
0020
0020
0020
001F
001F
001F
001F
0020
0020
0020
0020
0020
0020
0020
0020
0021
0020
0020
0020
0020
0020
0020
0020
0021
0021
0021
0020
0020
0020
0020
0020
0020
0021
0021
0021
0022
0022
0022
0022
0021
0021
0021
0022
0022
0022
0021
0020
0021
0022
0022
0022
0022
0023
0024
0023
0022
0022
0024
0024
0024
0023
0023
0023
0023
0023
0023
0023
0024
0024
0024
0024
0024
0024
0023
0023
0023
0024
0025
0025
0025
0025
0024
0024
0025
0025
0025
0025
0024
0024
0024
0025
0025
0025
0025
0025
0025
0025
0025
0026
0026
0026
0025
0026
0026
0026
0025
0025
0026
0026
0026
0026
0026
0027
0027
0026
0026
0026
0027
0027
0026
0026
0026
0026
0026
0026
0027
0028
0028
0027
0026
0026
0027
0028
0028
0027
0028
0029
002A
0029
0028
0028
0029
0029
0028
0028
0028
0028
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
002A
0029
0029
0029
002A
002A
002A
002A
002A
002A
002A
002A
0029
0029
002A
002A
002A
002A
002B
002C
002B
002A
002A
002B
002B
002B
002B
002B
002B
002B
002A
002A
002B
002B
002B
002B
002B
002B
002C
002C
002B
002B
002B
002C
002C
002C
002C
002B
002B
002B
002C
002C
002C
002B
002C
002C
002D
002D
002D
002D
002C
002B
002B
002B
002C
002D
002C
002C
002C
002D
002D
002C
002C
002C
002D
002E
002D
002D
002D
002D
002E
002D
002D
002D
002D
002D
002C
002B
002B
002C
002C
002C
002B
002C
002E
002E
002F
002E
002F
002F
002E
002E
002E
002F
002F
002E
002E
002E
002E
002F
002F
002F
002F
002F
002F
002F
002F
002F
002F
0030
002F
002F
0030
0030
0030
0030
002F
002F
0030
0030
0030
0030
002F
0030
0030
0030
0030
002F
002F
0030
0030
0031
0031
0031
0031
0030
0030
0031
0031
0032
0032
0031
0031
0032
0034
0035
0034
0033
0032
0031
0032
0032
0032
0032
0032
0032
0032
0032
0032
0032
0032
0032
0032
0033
0032
0032
0032
0033
0033
0033
0033
0033
0033
0034
0033
0032
0033
0034
0034
0033
0032
0033
0034
0034
0032
0032
0033
0034
0035
0034
0034
0034
0034
0034
0034
0034
0034
0034
0033
0033
0034
0035
0034
0033
0033
0034
0035
0035
0034
0034
0034
0034
0035
0035
0036
0036
0035
0035
0036
0036
0036
0035
0035
0035
0035
0035
0035
0036
0036
0036
0036
0036
0036
0037
0037
0036
0036
0036
0037
0036
0036
0036
0036
0037
0037
0037
0036
0036
0036
0036
0036
0037
0036
0036
0036
0037
0037
0038
0038
0037
0036
0036
0037
0038
0038
0038
0037
0037
0037
0037
0037
0038
0038
0037
0036
0036
0037
0038
0039
0038
0038
0038
0038
0038
0038
0038
0038
0039
0039
0039
0039
0039
0039
0038
0038
0039
0039
0039
0039
0039
0039
0038
0037
0037
0038
0039
0038
0038
0038
0038
0038
0037
0037
0038
0039
0038
0038
0038
0038
0039
0039
0039
0038
0039
0039
0039
0039
0039
0039
0038
0038
0039
0039
0038
0038
0038
0038
0039
0039
0039
0039
0039
0039
0039
0039
0039
0039
003A
003A
003B
003B
003B
003A
003A
003A
003B
003B
003A
003A
003A
003B
003B
003C
003C
003B
003B
003B
003C
003C
003C
003D
003C
003B
003B
003B
003B
003C
003B
003B
003C
003C
003C
003C
003C
003C
003C
003B
003B
003B
003B
003C
003C
003C
003D
003D
003D
003C
003C
003C
003C
003C
003D
003D
003C
003C
003C
003D
003D
003D
003C
003C
003D
003D
003D
003D
003D
003E
003E
003E
003D
003C
003C
003C
003C
003C
003C
003D
003D
003D
003D
003D
003C
003D
003D
003E
003D
003D
003C
003D
003F
003F
003D
003D
003D
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003F
003F
003E
003E
003E
003F
003F
003F
003E
003E
003E
003F
003F
003F
003E
003E
003E
003E
003E
003F
003F
003F
003F
003F
003F
003F
003F
003F
003F
0040
0040
0040
003E
003E
003F
0040
0040
003F
003F
0040
0040
0040
003F
0040
0040
0040
0040
0040
0041
0042
0041
0040
0040
0040
0040
003F
003F
003F
0040
0040
0040
0041
0041
0041
0040
0040
0040
0040
0041
0041
0041
0041
0041
0041
0040
0041
0041
0042
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0042
0042
0042
0042
0041
0041
0041
0042
0042
0042
0042
0041
0040
0041
0041
0042
0042
0041
0042
0042
0043
0042
0042
0041
0042
0042
0043
0043
0043
0043
0043
0044
0044
0043
0043
0043
0044
0044
0043
0043
0043
0043
0043
0043
0043
0044
0044
0043
0043
0043
0043
0043
0043
0043
0043
0042
0042
0042
0043
0044
0044
0044
0043
0042
0043
0043
0043
0043
0043
0044
0044
0044
0044
0044
0043
0043
0043
0043
0044
0044
0044
0044
0044
0044
0044
0044
0043
0043
0043
0043
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0045
0045
0045
0045
0044
0044
0044
0044
0044
0044
0044
0045
0045
0044
0043
0042
0044
0045
0045
0045
0044
0044
0045
0045
0045
0045
0044
0045
0045
0045
0045
0045
0045
0044
0044
0044
0045
0046
0046
0045
0044
0043
0044
0045
0046
0046
0045
0045
0045
0045
0045
0045
0045
0045
0045
0044
0044
0045
0045
0045
0045
0044
0044
0044
0044
0044
0045
0045
0045
0045
0045
0046
0046
0046
0045
0045
0046
0047
0047
0046
0045
0046
0046
0046
0046
0046
0047
0047
0046
0046
0046
0046
0046
0046
0046
0046
0046
0046
0047
0047
0047
0046
0046
0046
0047
0047
0046
0046
0046
0047
0047
0047
0047
0047
0046
0046
0046
0047
0047
0046
0046
0046
0047
0047
0046
0046
0046
0046
0047
0047
0046
0046
0046
0046
0047
0048
0049
0049
0049
0049
0049
0048
0048
0049
004A
004A
0049
0048
0048
0049
004A
004A
004A
0049
0049
0049
0049
0049
0049
0049
0049
0048
0049
0049
0049
0049
0049
0049
0049
0049
0049
0048
0048
0048
0048
0048
0049
0049
0049
0049
0049
0049
0049
0049
0049
0048
0048
0048
0049
0049
0049
0049
0048
0048
0048
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0048
0048
0048
0048
0048
0048
0048
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0048
0048
0048
0049
004A
004A
004A
004A
004A
004A
004A
004A
004A
004A
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
0049
004A
004A
004A
0049
0049
0049
004A
0049
0049
0049
0049
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
0049
0049
0049
0049
004A
004A
004A
004A
0049
0049
0049
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
0049
004A
004A
004A
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
004A
004A
004A
0049
0049
004A
004A
004B
004B
004A
0049
0048
0049
004A
004A
004A
0048
0048
0049
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
004A
004A
004A
004B
004B
004B
004B
004B
004B
004A
004A
0049
004A
004A
004A
004A
0049
0049
004A
004A
004B
004B
004B
004B
004A
004A
004A
004A
004A
004A
004B
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
004A
0049
0049
0049
0049
0049
0049
0049
004A
004B
004B
004A
004A
004A
004B
004B
004A
004A
004A
004B
004B
004B
004B
004B
004B
004B
004A
004A
004A
004A
004A
004A
004A
004A
004A
004A
004B
004B
004A
004A
0049
0049
004A
004A
004B
004A
004B
004A
004A
0049
004A
004B
004B
004B
004A
004A
004A
004B
004A
004A
004A
004B
004B
004B
004A
004A
004A
004B
004C
004E
004E
004D
004B
004A
004A
004A
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004B
004B
004C
004B
004A
004A
004A
004B
004B
004B
004B
004B
004A
004A
004A
004B
004B
004B
004B
004B
004B
004B
004B
004B
004B
004C
004C
004B
004B
004B
004A
004B
004C
004C
004C
004C
004B
004B
004B
004B
004B
004A
004A
004B
004B
004C
004C
004B
004B
004B
004C
004C
004B
004A
004A
004B
004B
004A
0049
0049
004A
004B
004B
004B
004A
004A
004B
004B
004B
004B
004A
004A
004B
004B
004B
004B
004A
004A
004B
004B
004B
004A
004A
004A
004B
004B
004C
004C
004B
004B
004B
004B
004B
004C
004C
004B
004B
004C
004D
004C
004B
004B
004B
004C
004C
004C
004B
004B
004B
004B
004B
004B
004B
004A
004A
004A
004B
004B
004C
004C
004C
004C
004C
004C
004C
004C
004C
004C
004B
004C
004C
004B
004B
004B
004C
004B
004B
004B
004C
004C
004C
004B
004A
004A
004A
004A
004A
004A
004A
0049
0049
0049
004A
004B
004B
004A
004A
0049
0048
0049
004A
004B
004B
004A
004A
004A
004A
0049
0049
004A
004A
004A
0049
0049
004A
004A
004A
0049
004A
004A
004B
004B
004B
004B
004A
004A
004A
004A
004A
004A
004A
004A
004A
004A
004A
004B
004B
004C
004B
004B
004B
004C
004C
004B
004B
004A
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004A
004B
004B
004B
004A
004A
004A
004A
004A
004A
004A
004B
004B
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004B
004B
004A
004A
004A
004A
004A
004A
004A
004A
004B
004B
004B
004B
004C
004C
004B
004A
004A
004B
004B
004B
004A
004A
004A
004A
004A
004A
004B
004B
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004B
004C
004C
004B
004B
004B
004B
004B
004B
004B
004A
004A
004B
004B
004B
004B
004A
004A
004B
004B
004A
004A
004A
004B
004B
004B
004B
004B
004B
004A
004A
004A
004B
004B
004A
004A
004A
004A
004A
004A
004B
004B
004B
004A
004A
004B
004B
004B
004A
004A
004B
004B
004B
004A
004A
004B
004C
004B
004B
004B
004C
004C
004C
004B
004B
004C
004C
004C
004B
004B
004B
004B
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004C
004C
004C
004B
004A
004B
004C
004D
004C
004B
004B
004B
004C
004B
004B
004B
004B
004B
004A
004A
004A
004B
004C
004C
004C
004C
004C
004B
004B
004B
004C
004C
004C
004C
004B
004B
004B
004B
004B
004B
004C
004C
004C
004B
004B
004B
004B
004B
004B
004A
004A
004B
004B
004B
004B
004A
004B
004C
004D
004D
004C
004B
004A
004B
004D
004D
004B
004A
004A
004B
004B
004B
004B
004C
004B
004B
004A
004B
004B
004B
004A
004A
004A
004B
004C
004B
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004B
004B
004B
004A
004A
004B
004B
004A
004A
004A
004B
004C
004B
004B
004A
004A
004B
004C
004C
004B
004A
004A
004B
004B
004B
004B
004B
004B
004A
004A
004A
004B
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004A
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
004A
004A
0049
004A
004A
004A
004A
0049
0049
004A
004B
004A
004A
004A
004A
004A
004A
004A
004A
0049
0049
004A
004A
004A
004A
0049
0049
004A
004B
004B
004B
004A
004A
004A
004A
004B
004B
004A
004A
0049
004A
004A
004B
004B
004B
004A
004B
004B
004A
004A
004A
004A
004B
004A
0049
0049
004A
0049
0049
0049
0049
004A
004A
004A
004A
004A
0049
0049
004A
004A
004A
004A
004A
004A
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
0049
004A
004A
004A
004A
004A
004A
004A
004A
0049
0049
004A
004A
004A
0049
0049
0049
0048
0049
0049
004A
004A
0049
0049
004A
004B
004B
004B
004B
004C
004C
004C
004C
004B
004B
004B
004B
004B
004B
004B
004B
004B
004A
004B
004B
004B
004A
0049
004A
004A
004B
004B
004B
004B
004B
004B
004B
004B
004A
004A
004A
004A
004A
004A
004A
004A
0049
0049
0049
004A
004A
004A
004A
004A
004A
004A
0049
0049
004A
004B
004B
004B
004A
004A
004A
004A
004B
004B
004A
0049
0048
0048
0049
004A
0049
0049
004A
004A
004B
004A
004A
004A
004A
004A
0049
0049
004A
004B
004A
0049
0048
0049
0049
0049
0048
0048
0048
0048
0049
0049
0049
004A
004A
0049
0049
0048
0048
0049
0049
004A
004A
0049
0049
0049
004A
004A
0049
0048
0048
0048
0048
0049
0049
0049
0048
0048
0048
0049
0049
0049
0048
0048
0049
0049
0048
0048
0049
0049
004A
0049
0049
0049
0048
0048
0048
0048
0049
0049
0048
0048
0048
0048
0048
0048
0048
0048
0048
0048
0048
0048
0048
0048
0048
0049
004A
0049
0048
0048
0048
0049
0048
0047
0047
0048
0048
0048
0047
0047
0048
0047
0047
0047
0047
0048
0047
0047
0047
0048
0048
0048
0047
0047
0047
0048
0048
0048
0048
0047
0047
0047
0048
0048
0047
0047
0047
0047
0047
0046
0046
0046
0047
0047
0047
0046
0046
0047
0047
0047
0046
0046
0046
0047
0047
0047
0047
0047
0047
0046
0046
0045
0046
0046
0046
0046
0046
0046
0046
0046
0046
0047
0047
0047
0046
0046
0046
0046
0047
0047
0046
0046
0045
0046
0046
0047
0047
0046
0045
0045
0045
0045
0045
0043
0043
0044
0046
0046
0046
0045
0046
0046
0047
0046
0045
0045
0046
0047
0047
0047
0046
0045
0045
0046
0047
0047
0046
0045
0045
0045
0045
0045
0046
0046
0046
0046
0045
0046
0046
0045
0045
0045
0045
0046
0046
0046
0045
0045
0045
0046
0046
0046
0046
0046
0045
0044
0045
0046
0046
0046
0045
0045
0045
0046
0046
0045
0046
0047
0048
0048
0046
0045
0045
0045
0045
0045
0045
0046
0046
0046
0045
0045
0045
0045
0045
0045
0045
0044
0044
0044
0045
0045
0045
0045
0045
0045
0045
0045
0044
0044
0044
0044
0044
0045
0046
0046
0045
0044
0044
0044
0044
0044
0044
0045
0046
0046
0045
0044
0044
0045
0045
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0045
0045
0044
0044
0044
0044
0044
0044
0044
0044
0044
0044
0045
0045
0044
0044
0044
0044
0044
0045
0045
0045
0044
0044
0044
0044
0044
0043
0044
0044
0044
0044
0043
0043
0044
0044
0043
0044
0045
0045
0044
0043
0043
0044
0045
0045
0044
0044
0044
0044
0043
0043
0044
0044
0045
0044
0044
0044
0043
0043
0042
0042
0043
0044
0044
0044
0043
0043
0043
0043
0043
0043
0044
0044
0044
0044
0043
0043
0044
0044
0044
0044
0044
0044
0044
0043
0043
0043
0043
0043
0043
0043
0043
0043
0043
0042
0042
0042
0042
0041
0041
0042
0042
0043
0043
0043
0042
0042
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0042
0042
0043
0043
0042
0041
0040
0041
0041
0042
0042
0042
0042
0042
0042
0041
0040
0040
0041
0042
0042
0042
0041
0041
0040
0040
0041
0042
0042
0042
0042
0042
0042
0041
0041
0041
0042
0042
0042
0042
0042
0042
0041
0041
0041
0041
0041
0041
0041
0041
0042
0042
0042
0041
0041
0040
0040
0040
0041
0041
0041
0041
0042
0042
0042
0042
0042
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0041
0040
0040
0040
0041
0041
0040
0040
0040
0040
0041
0040
0040
0041
0041
0041
0041
0040
0041
0041
0041
0041
0040
0041
0041
0041
0040
0040
0040
0041
0041
0041
0040
003F
003F
0041
0042
0043
0042
0040
003F
0040
0040
0041
0041
0041
0041
0040
0040
0040
0040
0041
0041
0041
0041
0040
0040
003F
003F
003F
0040
0040
0041
0041
0041
0040
003F
0040
0040
0041
0040
0040
0040
0040
003F
003F
003F
0040
0040
0040
0040
0040
0040
003F
003F
003F
0040
0040
0040
003F
003F
0040
0041
0040
003F
003F
003F
0040
0040
003F
003F
003F
0040
0040
0040
0040
0040
0040
003F
0040
0040
0041
0040
0040
0040
0041
0042
0041
003F
003E
003F
0040
0041
0040
003F
003F
0040
0040
003F
003F
003F
0040
0040
0040
003F
003F
0040
0040
003F
003F
003F
0040
0040
0040
003F
003E
003F
0040
0040
0040
0040
0040
0040
0040
003F
003F
0040
0040
003F
003F
003E
003E
003E
003F
003F
0040
003F
003F
003E
003E
003E
003E
003F
003F
003F
003F
003F
003F
003F
003F
003F
003F
003F
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003F
003F
003F
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003E
003D
003D
003E
003F
003F
003F
003E
003E
003E
003E
003D
003D
003E
003E
003E
003D
003D
003E
003E
003E
003D
003C
003C
003D
003E
003F
003E
003E
003E
003E
003E
003E
003D
003D
003D
003E
003E
003D
003D
003D
003D
003D
003D
003E
003E
003D
003D
003D
003D
003E
003D
003D
003D
003D
003D
003D
003C
003C
003C
003C
003C
003C
003C
003C
003C
003D
003D
003D
003C
003B
003B
003D
003D
003D
003C
003B
003C
003C
003C
003C
003C
003C
003C
003C
003D
003C
003C
003C
003C
003C
003C
003B
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003D
003D
003C
003B
003A
003B
003C
003C
003C
003B
003B
003C
003C
003C
003C
003C
003C
003C
003B
003B
003B
003B
003C
003C
003B
003B
003B
003B
003C
003C
003C
003B
003A
003B
003B
003B
003A
003B
003B
003B
003B
003B
003B
003C
003C
003B
003B
003B
003A
003A
003A
003B
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003C
003B
003B
003B
003C
003B
003B
003B
003C
003C
003C
003B
003B
003C
003D
003D
003B
003B
003B
003C
003C
003C
003C
003C
003C
003B
003A
003A
003A
003A
003B
003B
003B
003B
003B
003B
003C
003C
003C
003B
003B
003B
003B
003C
003B
003B
003A
003B
003B
003C
003C
003B
003B
003B
003B
003B
003B
003B
003B
003A
003A
003B
003B
003A
003A
003A
003A
003A
003A
003A
003B
003B
003B
003A
0039
003A
003B
003B
003B
003A
003A
003A
003B
003A
003A
0039
0039
0039
0039
0039
0039
0039
0039
003A
003A
003A
0039
003A
003A
003A
0039
0039
0039
003A
003A
0039
0038
0038
0039
0039
0038
0038
0039
0039
0039
0039
0038
0039
003A
003A
0039
0038
0037
0037
0038
0038
0039
0039
0038
0038
0038
0038
0038
0038
0038
0038
0038
0038
0039
0039
0039
0039
0039
0039
0038
0038
0038
0037
0037
0038
0038
0038
0038
0038
0038
0039
0038
0038
0038
0039
0039
0038
0037
0038
0038
0038
0038
0037
0038
0038
0037
0037
0037
0038
0038
0038
0037
0037
0038
0038
0038
0037
0037
0037
0036
0036
0036
0037
0037
0037
0037
0036
0036
0037
0038
0038
0038
0037
0037
0037
0036
0036
0036
0037
0037
0037
0036
0036
0037
0037
0036
0036
0036
0037
0036
0036
0035
0036
0036
0036
0036
0035
0035
0036
0036
0036
0036
0035
0035
0035
0036
0036
0036
0036
0036
0036
0035
0034
0035
0036
0037
0036
0035
0034
0034
0034
0034
0033
0034
0035
0035
0035
0035
0035
0035
0035
0035
0036
0035
0034
0034
0034
0036
0036
0036
0035
0035
0035
0035
0035
0036
0036
0036
0035
0034
0035
0036
0036
0036
0035
0035
0035
0034
0034
0034
0035
0035
0036
0036
0035
0035
0034
0034
0035
0035
0036
0036
0035
0035
0034
0034
0035
0035
0035
0034
0035
0035
0035
0034
0034
0035
0037
0038
0037
0035
0034
0034
0035
0035
0035
0034
0035
0035
0035
0035
0034
0034
0034
0034
0033
0033
0033
0034
0035
0034
0033
0033
0034
0034
0034
0033
0034
0035
0035
0034
0033
0033
0033
0034
0033
0033
0033
0034
0035
0035
0034
0033
0033
0033
0033
0033
0034
0034
0034
0034
0033
0034
0035
0035
0034
0034
0033
0033
0033
0033
0034
0034
0034
0033
0033
0033
0033
0034
0033
0033
0034
0034
0033
0032
0032
0032
0032
0033
0032
0033
0033
0033
0033
0033
0033
0033
0033
0033
0032
0032
0032
0032
0033
0034
0034
0034
0033
0032
0032
0032
0032
0032
0033
0033
0033
0033
0033
0033
0033
0032
0032
0032
0033
0033
0032
0032
0032
0032
0032
0032
0031
0032
0032
0032
0032
0031
0031
0031
0032
0032
0031
0031
0031
0031
0031
0031
0033
0033
0033
0032
0031
0031
0030
0031
0031
0032
0032
0032
0032
0032
0032
0032
0031
0031
0030
0030
0030
0030
0030
0030
0031
0031
0030
0030
002F
0030
0030
0030
0030
0030
002F
002F
0030
0031
0030
002F
002F
0030
0031
0030
002E
002E
002F
002F
002F
002F
002F
0030
0030
002F
002F
002F
002F
002F
002F
002F
0030
0031
0031
0030
002F
002F
002F
0030
0030
0030
0030
0030
0030
0030
0030
002F
002F
0030
0030
002F
002F
0030
0031
0031
0030
002F
002F
002F
002F
002F
002E
002F
002F
0030
0030
0030
0030
002F
002F
0030
0030
0030
0030
0030
002F
002F
002E
002F
0030
0030
0031
0030
002F
002F
002E
002E
002F
002F
002F
002F
002E
002E
002E
002E
002E
002E
002F
002F
0030
002F
002F
002F
002E
002E
002F
002F
002F
002F
002E
002E
002E
002E
002E
002E
002E
002E
002E
002E
002F
002F
002E
002E
002E
002F
002F
002F
002F
002F
002F
002E
002E
002E
002E
002E
002D
002C
002C
002D
002D
002D
002D
002E
002E
002E
002E
002D
002D
002E
002E
002E
002E
002E
002E
002E
002E
002D
002D
002D
002D
002D
002D
002D
002D
002E
002E
002E
002D
002D
002E
002E
002E
002E
002E
002D
002D
002D
002E
002E
002E
002D
002D
002E
002E
002E
002E
002E
002E
002E
002E
002D
002D
002D
002C
002D
002E
002E
002E
002E
002D
002D
002D
002D
002D
002D
002D
002D
002D
002D
002D
002D
002D
002D
002E
002E
002E
002E
002D
002D
002D
002E
002E
002E
002D
002C
002C
002C
002D
002D
002D
002D
002D
002D
002D
002E
002E
002D
002C
002D
002D
002D
002C
002C
002C
002D
002D
002D
002D
002C
002C
002C
002D
002D
002D
002D
002D
002D
002D
002D
002C
002C
002C
002D
002D
002C
002C
002C
002C
002C
002C
002C
002C
002D
002D
002C
002C
002C
002C
002C
002C
002B
002B
002B
002C
002C
002C
002C
002D
002D
002C
002B
002B
002C
002D
002C
002B
002A
002B
002C
002C
002C
002C
002C
002C
002B
002B
002B
002B
002B
002B
002B
002B
002B
002B
002C
002C
002B
002B
002B
002B
002B
002C
002C
002C
002C
002C
002B
002B
002B
002B
002B
002B
002B
002B
002B
002B
002B
002A
002A
002B
002C
002C
002C
002B
002B
002B
002B
002B
002B
002A
002A
002A
002B
002B
002A
002A
002A
002A
002A
002A
0029
0029
002A
002B
002B
002B
002B
002B
002B
002B
002A
002A
002A
002B
002A
002A
0029
0029
0029
0029
0029
002A
002B
002B
002B
002A
002A
002A
002A
002A
0029
0029
002A
002A
002A
0029
0029
002A
002A
002A
0029
0028
0029
002A
002A
0029
002A
002B
002A
0029
0028
0029
002A
002A
002A
002A
002A
002B
002B
002A
002A
002A
002A
0029
002A
002A
002A
0029
0028
0029
0029
002A
0029
0029
0029
002A
002A
002A
0029
0028
0029
0029
002A
002A
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0029
0028
0028
0029
0029
0029
0028
0028
0028
0029
002A
0029
0028
0028
0028
0029
0029
002A
002A
002A
002A
002A
002A
002A
002A
002A
002A
002A
002A
002A
002A
0029
0029
0029
0029
0029
002A
002A
0029
0029
0029
0029
002A
0029
0029
0028
0029
002A
002A
0029
0029
0029
0029
0029
0029
002A
002A
002A
0029
0028
0028
0029
002A
002A
0029
0029
0029
0028
0028
0028
0029
0029
0028
0027
0028
0028
0029
0029
0028
0028
0028
0028
0028
0028
0028
0029
0029
0028
0028
0028
0028
0028
0028
0028
0028
0028
0027
0028
0028
0029
0028
0028
0027
0028
0028
0028
0028
0028
0028
0028
0028
0028
0027
0028
0028
0028
0028
0027
0027
0027
0028
0028
0027
0026
0026
0027
0027
0026
0026
0027
0027
0027
0026
0026
0025
0026
0027
0027
0027
0028
0028
0027
0026
0025
0025
0026
0026
0027
0027
0027
0026
0026
0026
0027
0027
0027
0027
0027
0027
0026
0026
0026
0026
0026
0026
0025
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0026
0027
0026
0025
0025
0025
0026
0027
0026
0025
0025
0025
0025
0025
0025
0025
0026
0026
0025
0024
0024
0025
0025
0025
0025
0025
0025
0025
0025
0026
0026
0025
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0024
0023
0023
0022
0023
0024
0024
0024
0024
0023
0023
0023
0023
0023
0024
0024
0024
0024
0024
0024
0024
0023
0023
0023
0023
0024
0024
0024
0023
0022
0021
0021
0022
0022
0021
0021
0021
0022
0022
0023
0023
0023
0024
0024
0023
0022
0023
0023
0024
0023
0022
0022
0023
0023
0023
0023
0023
0023
0023
0023
0023
0023
0022
0021
0021
0022
0023
0022
0022
0022
0022
0023
0023
0023
0023
0023
0022
0022
0022
0023
0023
0022
0021
0022
0023
0024
0023
0021
0021
0022
0022
0023
0022
0022
0022
0022
0023
0024
0025
0024
0023
0022
0022
0022
0022
0022
0022
0022
0022
0022
0022
0022
0022
0022
0022
0022
0023
0023
0022
0021
0021
0021
0022
0022
0022
0022
0021
0021
0022
0022
0022
0022
0022
0022
0022
0021
0021
0021
0022
0022
0022
0022
0022
0021
0021
0021
0021
0022
0022
0022
0022
0022
0021
0021
0021
0021
0022
0022
0021
0021
0021
0021
0021
0021
0020
0021
0021
0022
0021
0020
0020
0020
0021
0021
0021
0021
0021
0021
0021
0021
0021
0022
0021
0021
0021
0021
0021
0021
0020
0020
0020
0020
0020
0020
0020
0021
0021
0020
0020
0020
0020
0020
0020
0020
0021
0021
0021
0020
0020
0020
0020
0020
0020
0020
0021
0021
0021
0021
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0020
0021
0021
0021
0021
0021
0021
0020
001F
001F
0020
0021
0021
0021
0020
0020
0020
0020
0020
001F
001F
001F
0020
0020
0020
001F
001E
001E
001E
001F
001F
001F
001F
001F
001F
001F
001E
001E
001E
001E
001E
001E
001E
001E
001E
001E
001E
001E
001F
001F
001F
001F
001E
001E
001D
001D
001E
001E
001E
001F
001E
001E
001D
001D
001E
001E
001E
001D
001D
001E
001F
001E
001D
001D
001D
001E
001E
001D
001D
001D
001E
001E
001E
001E
001E
001E
001E
001E
001E
001F
001F
001E
001D
001D
001D
001E
001E
001E
001E
001E
001D
001D
001D
001D
001D
001D
001E
001F
001E
001E
001D
001D
001D
001E
001D
001D
001D
001D
001E
001D
001D
001C
001D
001D
001D
001D
001C
001C
001C
001D
001D
001D
001D
001D
001E
001E
001E
001D
001D
001D
001D
001C
001C
001C
001D
001D
001D
001D
001D
001D
001D
001D
001C
001D
001E
001E
001E
001D
001D
001D
001E
001E
001D
001D
001D
001D
001D
001D
001D
001C
001C
001C
001D
001D
001D
001D
001C
001C
001B
001B
001C
001D
001D
001C
001C
001C
001D
001D
001C
001B
001C
001C
001D
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001D
001D
001D
001C
001C
001C
001D
001D
001D
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001C
001B
001C
001C
001C
001C
001C
001C
001C
001B
001B
001C
001D
001D
001C
001B
001B
001D
001D
001D
001C
001B
001B
001B
001B
001B
001B
001C
001C
001B
001A
001B
001C
001C
001C
001C
001C
001C
001C
001C
001C
001B
001B
001B
001B
001B
001B
001C
001D
001C
001B
001B
001B
001B
001B
001B
001B
001C
001B
001B
001A
001B
001A
001A
0019
001A
001B
001B
001B
001A
001B
001D
001D
001C
001B
001B
001B
001B
001B
001A
001B
001C
001C
001B
001A
001B
001B
001C
001B
001A
001A
001B
001C
001C
001C
001B
001B
001A
0019
0019
0019
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001A
001B
001B
001B
001A
0019
001A
001B
001B
001A
001A
001A
001A
001A
0019
0019
001A
001A
0019
0019
0019
001A
001A
001A
0019
0019
0019
001A
001A
001B
001B
001A
0019
0019
0019
001A
001A
0019
0018
0019
0019
001A
0019
0019
0019
001A
001A
0019
0019
0019
001A
0019
0019
0018
0019
001A
001A
001A
0019
0019
0019
001A
0019
0019
0019
0019
0019
0019
0019
001A
001A
001A
0019
0019
0018
0018
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0018
0018
0018
0019
0019
0019
0019
0019
0019
0019
0019
0018
0018
0019
0019
0019
0019
0019
0019
0018
0017
0017
0018
0018
0018
0018
0018
0018
0018
0018
0018
0019
0019
0019
0018
0018
0018
0018
0018
0017
0018
0018
0018
0018
0018
0017
0017
0017
0018
0018
0018
0017
0017
0018
0018
0018
0018
0018
0018
0018
0019
001A
001A
0019
0019
0019
001A
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0019
0018
0018
0018
0018
0019
0019
0019
0019
0019
0019
0018
0018
0018
0018
0019
0019
0019
0019
0019
0018
0018
0018
0018
0018
0018
0018
0018
0017
0017
0017
0018
0018
0018
0018
0018
0018
0019
0018
0018
0018
0017
0018
0018
0018
0018
0018
0018
0018
0019
0018
0017
0017
0018
0019
0019
0018
0018
0018
0018
0017
0017
0018
0018
0018
0017
0017
0018
0018
0017
0016
0016
0017
0018
0018
0018
0018
0017
0017
0017
0017
0017
0017
0017
0017
0017
0017
0017
0017
0017
0017
0017
0016
0016
0016
0016
0016
0016
0016
0016
0017
0017
0017
0016
0016
0015
0015
0016
0017
0017
0016
0016
0016
0016
0016
0016
0016
0017
0017
0017
0016
0016
0016
0015
0015
0015
0016
0016
0015
0015
0015
0015
0015
0015
0015
0016
0016
0015
0015
0016
0016
0016
0015
0015
0015
0016
0016
0016
0015
0015
0015
0015
0015
0015
0015
0015
0015
0015
0015
0015
0014
0014
0014
0015
0015
0015
0015
0015
0015
0015
0014
0014
0014
0015
0015
0015
0014
0014
0014
0014
0014
0014
0015
0015
0015
0015
0014
0013
0013
0014
0015
0016
0015
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0014
0013
0013
0013
0014
0014
0014
0013
0013
0014
0014
0013
0011
0011
0011
0012
0012
0011
0011
0012
0013
0013
0013
0013
0014
0014
0013
0012
0013
0014
0014
0013
0012
0012
0013
0013
0014
0013
0012
0012
0012
0013
0013
0013
0013
0013
0013
0013
0013
0012
0012
0013
0014
0013
0013
0012
0013
0013
0014
0013
0013
0013
0013
0012
0013
0013
0013
0014
0014
0013
0013
0012
0011
0012
0013
0013
0012
0011
0013
0016
0017
0016
0014
0013
0012
0012
0012
0012
0012
0013
0013
0013
0012
0012
0012
0013
0013
0013
0012
0012
0013
0014
0014
0013
0012
0012
0013
0014
0013
0013
0013
0013
0013
0012
0013
0013
0014
0013
0013
0013
0013
0013
0012
0012
0012
0013
0013
0012
0012
0013
0012
0012
0012
0012
0012
0013
0013
0013
0013
0013
0013
0012
0012
0012
0013
0013
0013
0012
0012
0012
0012
0012
0012
0011
0011
0011
0011
0012
0011
0011
0011
0012
0012
0012
0012
0011
0011
0011
0011
0012
0012
0011
0011
0012
0012
0012
0012
0012
0012
0012
0012
0012
0012
0012
0012
0013
0013
0013
0012
0011
0011
0011
0012
0012
0011
0011
0012
0013
0013
0012
0011
0011
0012
0012
0011
0011
0011
0012
0012
0011
0010
0010
0011
0012
0011
0011
0010
0011
0011
0012
0012
0012
0012
0012
0012
0011
0011
0011
0011
0012
0012
0012
0012
0012
0012
0012
0012
0012
0011
0011
0011
0011
0010
000F
000F
000F
0010
0010
0010
000F
000F
000F
000F
0010
0010
0010
0010
0010
0010
0010
000F
000F
000F
0010
0010
0010
000F
000F
000F
000F
000F
000F
000F
000F
000F
0010
0010
0010
0010
0010
0010
0010
000F
000F
000F
000F
000F
000F
000F
0010
000F
000F
000F
0010
0011
0011
0010
000F
0010
0010
0010
000F
0010
0010
0010
000F
000F
000F
0010
0010
0010
0010
0010
0010
000F
000E
000E
000F
0010
000F
000F
000F
000F
000F
000F
0010
0010
0010
0010
0010
0010
0010
0010
000F
000F
000F
000F
000F
000F
000E
000E
000E
000F
000F
0010
0010
000F
000F
000E
000E
000E
000E
000F
000F
000F
000E
000E
000E
000E
000E
000E
000E
000E
000F
000F
000F
000F
000F
000F
000F
000F
000F
000F
000F
000E
000F
0010
0010
000F
000F
000E
000F
000F
000F
000E
000D
000D
000E
000E
000F
000F
000E
000E
000F
000F
000F
000F
000F
000F
000F
000F
000E
000E
000D
000D
000E
000F
000F
000F
000E
000E
000E
000E
000D
000E
000E
000F
000F
000E
000E
000E
000E
000E
000F
000F
000F
000F
000E
000D
000E
000F
0010
0010
000F
000F
000F
000F
000F
000F
000E
000E
000F
000F
000F
000F
000E
000E
000F
000F
000F
000F
000F
000F
000F
000F
000E
000E
000E
000F
0010
0010
000F
000F
000F
000F
000F
000E
000E
000E
000F
000F
000F
000E
000E
000F
000F
000E
000E
000E
000E
000E
000E
000E
000E
000E
000E
000E
000F
000F
000F
000F
000E
000E
000E
000E
000E
000E
000E
000E
000D
000D
000D
000D
000E
000E
000E
000D
000E
000E
000E
000E
000E
000F
000E
000E
000D
000E
000E
000F
000E
000E
000E
000E
000E
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000E
000E
000E
000D
000C
000C
000D
000E
000E
000E
000D
000D
000D
000D
000D
000D
000D
000D
000D
000E
000E
000D
000D
000D
000E
000E
000E
000E
000E
000E
000E
000E
000E
000E
000E
000E
000D
000D
000D
000D
000D
000E
000E
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000C
000C
000C
000C
000D
000D
000D
000D
000D
000D
000D
000E
000D
000C
000C
000D
000D
000D
000D
000C
000B
000C
000C
000C
000C
000C
000C
000C
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000D
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000B
000C
000D
000D
000D
000C
000C
000C
000C
000C
000C
000B
000B
000C
000C
000C
000D
000D
000C
000C
000C
000C
000D
000D
000C
000B
000B
000B
000C
000C
000C
000C
000C
000B
000C
000C
000C
000C
000C
000B
000C
000D
000E
000D
000C
000B
000B
000C
000C
000C
000B
000B
000C
000D
000D
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000B
000B
000C
000D
000D
000D
000D
000D
000D
000D
000C
000C
000D
000E
000E
000D
000C
000C
000D
000E
000D
000D
000C
000C
000B
000B
000B
000C
000D
000D
000C
000B
000C
000C
000D
000C
000C
000C
000C
000D
000D
000D
000C
000C
000C
000C
000C
000C
000C
000C
000C
000B
000B
000B
000C
000C
000B
000B
000B
000C
000C
000C
000C
000C
000C
000C
000C
000C
000B
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000C
000B
000B
000B
000B
000C
000B
000B
000B
000C
000C
000B
000B
000B
000B
000B
000B
000B
000B
000B
000B
000A
000B
000C
000B
000A
000A
000A
000A
000A
000A
000A
000A
000A
000B
000B
000B
000B
000B
000A
000A
000B
000B
000B
000B
000B
000B
000A
000A
000B
000B
000B
000B
000B
000A
000A
000A
000A
000A
000A
000A
000A
0009
0009
0009
000A
000A
0009
0009
000A
000B
000B
000B
000A
000A
000A
000A
000A
000A
000A
000A
000A
000A
000A
000A
000A
000A
000A
000B
000B
000A
0009
0009
000A
000B
000B
000A
000A
000A
000A
000A
000A
000A
000A
0009
0009
0008
0009
0009
0009
0009
0009
0009
0008
0007
0008
0008
0009
0009
0009
0009
0009
0008
0009
0009
0009
0008
0008
0008
0009
0009
0009
0008
0009
0009
0009
0009
0008
0009
0009
0009
0008
0009
0009
0009
0009
0009
0009
0009
0008
0008
0008
0008
0008
0008
0008
0009
0009
0009
0008
0008
0009
0009
0009
0008
0008
0009
0008
0007
0006
0006
0007
0007
0006
0006
0006
0007
0008
0009
0008
0008
0008
0008
0008
0008
0008
0008
0008
0009
0009
0009
0008
0008
0008
0008
0008
0008
0008
0008
0008
0008
0007
0007
0008
0008
0008
0008
0008
0008
0008
0007
0007
0008
0008
0008
0007
0008
0009
0009
0009
0008
0008
0009
000A
0009
0008
0008
0008
0008
0008
0009
0009
0009
0008
0007
0009
000B
000B
000A
0009
0008
0007
0007
0008
0008
0009
0009
0008
0008
0008
0008
0008
0007
0007
0008
0008
0007
0007
0008
0009
0009
0008
0007
0008
0009
0008
0007
0007
0008
0009
0008
0007
0008
0008
0009
0008
0007
0008
0008
0008
0008
0007
0007
0007
0008
0008
0008
0008
0007
0007
0007
0007
0007
0006
0006
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0008
0008
0008
0008
0008
0008
0007
0007
0007
0007
0008
0008
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0007
0008
0008
0008
0007
0007
0006
0007
0007
0007
0007
0008
0009
0009
0009
0008
0007
0007
0007
0007
0006
0006
0006
0007
0008
0008
0007
0006
0006
0007
0008
0007
0006
0006
0006
0006
0007
0008
0008
0008
0007
0006
0006
0007
0006
0006
0006
0008
0008
0007
0005
0005
0006
0007
0006
0005
0006
0007
0007
0006
0005
0005
0005
0006
0006
0006
0005
0005
0005
0005
0006
0006
0005
0005
0005
0005
0005
0005
0005
0005
0005
0006
0006
0006
0006
0005
0005
0004
0005
0005
0005
0005
0005
0005
0004
0004
0005
0006
0006
0006
0005
0005
0005
0006
0006
0006
0006
0005
0005
0006
0006
0006
0005
0004
0005
0005
0005
0005
0005
0006
0007
0007
0006
0005
0005
0005
0005
0005
0004
0004
0004
0005
0005
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0005
0005
0004
0003
0003
0004
0004
0004
0004
0004
0004
0005
0005
0004
0004
0004
0005
0005
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0004
0005
0005
0005
0004
0004
0004
0004
0004
0004
0004
0005
0005
0005
0005
0005
0005
0005
0005
0006
0006
0005
0004
0004
0005
0005
0004
0004
0004
0005
0004
0004
0005
0006
0006
0005
0004
0004
0005
0005
0004
0004
0004
0005
0005
0004
0004
0004
0005
0005
0005
0004
0004
0004
0004
0004
0005
0005
0005
0005
0005
0005
0005
0005
0004
0004
0005
0005
0005
0005
0004
0004
0005
0005
0005
0004
0004
0005
0005
0006
0005
0005
0005
0005
0005
0005
0005
0004
0004
0004
0005
0005
0005
0005
0005
0005
0005
0006
0005
0005
0004
0005
0005
0006
0006
0005
0005
0006
0006
0006
0005
0004
0004
0005
0005
0004
0004
0004
0005
0005
0004
0004
0004
0005
0005
0005
0005
0005
0005
0004
0004
0004
0005
0004
0004
0005
0005
0005
0005
0005
0005
0005
0004
0004
0004
0005
0005
0005
0004
0003
0004
0005
0006
0006
0005
0003
0003
0004
0005
0005
0004
0004
0004
0005
0005
0004
0003
0003
0004
0004
0004
0005
0005
0005
0005
0004
0004
0003
0004
0004
0004
0004
0004
0004
0004
0005
0005
0004
0004
0005
0005
0005
0005
0005
0004
0004
0004
0004
0004
0004
0004
0004
0003
0003
0004
0004
0004
0004
0004
0004
0004
0003
0003
0003
0004
0005
0004
0004
0004
0004
0005
0004
0004
0004
0004
0004
0004
0003
0003
0003
0004
0004
0005
0005
0005
0005
0004
0003
0003
0004
0004
0004
0004
0004
0005
0005
0004
0003
0003
0003
0003
0003
0003
0004
0005
0004
0004
0003
0003
0004
0004
0003
0003
0003
0004
0004
0004
0004
0003
0004
0004
0004
0004
0004
0004
0004
0004
0004
0003
0003
0004
0005
0005
0004
0004
0004
0004
0004
0004
0004
0005
0005
0004
0004
0004
0004
0004
0003
0003
0004
0004
0003
0002
0002
0003
0003
0003
0002
0003
0004
0004
0004
0003
0003
0003
0003
0003
0004
0004
0004
0003
0003
0003
0004
0004
0004
0004
0004
0004
0003
0003
0003
0004
0004
0003
0003
0004
0003
0002
0002
0002
0003
0003
0003
0002
0003
0003
0004
0003
0003
0003
0004
0003
0003
0004
0004
0004
0003
0003
0003
0003
0003
0003
0003
0004
0004
0005
0005
0005
0005
0005
0005
0005
0005
0006
0006
0005
0005
0004
0004
0005
0005
0006
0006
0005
0004
0004
0005
0005
0005
0005
0005
0004
0004
0004
0004
0004
0004
0004
0004
0004
0005
0005
0005
0005
0005
0005
0005
0004
0004
0004
0004
0003
0003
0003
0004
0004
0004
0003
0003
0003
0003
0002
0003
0003
0003
0003
0003
0003
0004
0004
0003
0003
0004
0004
0004
0004
0003
0004
0004
0004
0004
0003
0004
0004
0004
0005
0005
0004
0004
0003
0003
0003
0003
0003
0003
0003
0003
0004
0004
0004
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0003
0002
0002
0003
0004
0003
0003
0003
0004
0004
0003
0002
0003
0004
0004
0004
0003
0003
0003
0003
0002
0002
0002
0003
0002
0002
0003
0003
0002
0002
0002
0003
0003
0002
0002
0003
0004
0004
0003
0002
0002
0002
0002
0003
0003
0003
0002
0002
0002
0002
0002
0001
0001
0002
0003
0003
0002
0002
0002
0002
0002
0002
0002
0002
0002
0002
0003
0004
0004
0003
0002
0002
0003
0003
0003
0002
0002
0002
0002
0002
0002
0003
0002
0001
0001
0002
0002
0002
0002
0002
0002
0002
0002
0001
0002
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0000
0001
0001
0001
0000
0000
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0002
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0000
0001
0002
0004
0004
0002
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0002
0002
0002
0001
0000
FFFF
0000
0001
0002
0001
0001
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0002
0002
0001
0000
FFFF
0000
0001
0001
0001
0001
0001
0002
0002
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0000
0000
0001
0001
0001
0001
0002
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
0000
0001
0001
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFC
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFF9
FFF8
FFF8
FFF8
FFF8
FFF9
FFF9
FFFB
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFE
FFFE
FFFD
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFD
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFD
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFA
FFFB
FFFA
FFFA
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFFA
FFFB
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFA
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFF9
FFF9
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFF9
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFF9
FFFA
FFFB
FFFB
FFFA
FFF9
FFFA
FFFB
FFFB
FFFB
FFFA
FFF9
FFF8
FFF8
FFF8
FFF9
FFF9
FFF9
FFF9
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFE
FFFE
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFF9
FFFA
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFF8
FFF8
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFB
FFFB
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFF9
FFFA
FFFA
FFFA
FFFA
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFF9
FFF9
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFF9
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFF9
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFB
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFF8
FFF9
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFB
FFFB
FFFD
FFFD
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFF8
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFF9
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFF9
FFFA
FFFA
FFFB
FFFA
FFFA
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFD
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFF9
FFF8
FFF9
FFF9
FFF8
FFF8
FFF8
FFF9
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFB
FFFC
FFFD
FFFD
FFFD
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFA
FFF9
FFF9
FFF9
FFF9
FFF9
FFF8
FFF9
FFF9
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFF9
FFFA
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFF9
FFF9
FFF9
FFFA
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFC
FFFC
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFA
FFF9
FFF9
FFF9
FFF9
FFF8
FFF9
FFFB
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFA
FFFB
FFFC
FFFE
FFFF
FFFF
FFFD
FFFB
FFFA
FFFB
FFFB
FFFB
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFB
FFFA
FFFA
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFF9
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFA
FFFB
FFFB
FFFC
FFFB
FFFB
FFFA
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFA
FFFB
FFFB
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFD
FFFF
0000
0001
FFFF
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFD
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFB
FFFB
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFC
FFFB
FFFA
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFB
FFFB
FFFB
FFFB
FFFC
FFFB
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFC
FFFB
FFFA
FFFB
FFFB
FFFB
FFFA
FFFB
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFF
0000
0000
FFFE
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFA
FFFA
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFB
FFFB
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFB
FFFB
FFFC
FFFD
FFFF
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFF
0001
0002
0000
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFC
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
0000
0001
0001
FFFF
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFD
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
0000
0000
FFFF
FFFE
FFFE
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFC
FFFC
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
0001
0002
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFC
FFFC
FFFD
FFFE
FFFD
FFFC
FFFC
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0001
0001
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFC
FFFC
FFFC
FFFD
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
0000
0001
0002
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFF
FFFF
FFFF
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFE
FFFE
FFFE
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFC
FFFC
FFFD
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0001
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFC
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0002
0002
0001
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0001
0002
0002
0001
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFE
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0001
0002
0002
0001
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0002
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0002
0002
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0002
0002
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0002
0002
0002
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0001
0003
0002
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0001
0002
0002
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0001
0002
0002
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0002
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0002
0003
0001
FFFF
FFFE
FFFF
0000
0001
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0002
0002
0001
0001
0000
0001
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
FFFF
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0003
0002
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFD
FFFC
FFFD
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0000
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0001
0003
0003
0002
0000
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0002
0002
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0001
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
0000
0001
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0002
0002
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0001
0002
0002
0000
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0002
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0002
0003
0003
0001
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0002
0002
0001
0000
0001
0001
0001
0001
0000
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0002
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0002
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0001
0000
0000
0000
0001
0003
0003
0001
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0001
0003
0002
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0001
0000
0000
0000
0001
0002
0002
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0002
0001
0001
0000
0001
0001
0001
0001
0001
0001
0002
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0001
0002
0002
0002
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0001
0002
0002
0001
0000
0000
0001
0001
0000
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
FFFF
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0002
0003
0003
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0002
0002
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0002
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0002
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
0000
0002
0002
0001
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0002
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0000
0000
FFFF
0000
0001
0002
0002
0001
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0001
0003
0002
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0002
0001
0001
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFD
FFFC
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0001
0003
0004
0002
0000
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0002
0003
0002
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0002
0002
0001
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0002
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0001
0002
0003
0002
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0002
0002
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0002
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0002
0002
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0000
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0001
0003
0002
0001
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0001
0000
0000
0001
0002
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0002
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFC
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0002
0002
0001
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0001
0002
0002
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0001
0001
0002
0002
0002
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0002
0002
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0001
0002
0003
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0002
0002
0002
0001
0000
0000
0000
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0002
0001
0001
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0002
0002
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0002
0003
0003
0001
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0002
0002
0002
0001
0000
0000
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0001
0002
0002
0000
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0002
0002
0002
0002
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0002
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0002
0002
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0001
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0001
0002
0002
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0001
0002
0002
0002
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
FFFF
0000
0001
0001
0001
0000
0000
0001
0001
0002
0002
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
FFFF
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0001
0003
0003
0001
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0002
0002
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0002
0003
0002
0001
0001
0001
0002
0002
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0002
0001
0000
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0001
0002
0002
0000
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0001
0002
0002
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0001
0002
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFC
FFFD
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0002
0003
0003
0002
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0002
0001
0001
0000
0000
0001
0001
0001
0002
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0002
0002
0002
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0002
0003
0003
0002
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0002
0002
0001
0001
0001
0001
0000
0001
0001
0002
0002
0002
0002
0002
0001
0001
0001
0001
0001
0001
0002
0002
0002
0002
0002
0002
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0001
0002
0003
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0002
0001
0000
0000
0000
0001
0002
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0000
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0002
0002
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0002
0001
0000
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0002
0001
0001
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0001
0002
0003
0002
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0002
0002
0001
0001
0000
0000
0001
0001
0001
0001
0001
0002
0002
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0002
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0001
0003
0003
0001
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
FFFF
FFFE
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0003
0003
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0000
0000
0001
0001
0001
0001
0002
0001
0001
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0002
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFE
FFFE
FFFE
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0002
0002
0001
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0002
0001
0000
0000
0001
0002
0001
0000
0000
0001
0002
0001
0001
0001
0001
0001
0000
0000
0001
0002
0002
0001
0000
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0003
0003
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0001
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0001
0003
0002
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0002
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0002
0003
0001
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0002
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0002
0002
0002
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0001
0001
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0002
0002
0002
0002
0002
0002
0001
0001
0002
0003
0003
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0002
0003
0002
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0002
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0002
0003
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFD
FFFD
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0002
0002
0002
0002
0002
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0002
0003
0003
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0001
0002
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0001
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0001
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0001
0002
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0002
0003
0002
0001
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0003
0003
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0001
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0002
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0002
0001
0000
0000
0001
0002
0001
0000
0000
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0002
0002
0001
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0001
0001
0000
0001
0001
0001
0000
0000
0000
0001
0002
0001
0001
0000
0000
0000
0000
0001
0001
0002
0002
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0002
0002
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0001
0000
FFFF
FFFF
0001
0003
0003
0002
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0002
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0002
0002
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0001
0002
0002
0001
0001
0001
0001
0002
0002
0002
0001
0001
0001
0002
0002
0002
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0002
0002
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
0000
0001
0001
0001
0001
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0002
0002
0002
0001
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFD
FFFD
FFFD
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
0000
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0002
0002
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0002
0002
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFE
FFFF
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0001
0001
0002
0002
0002
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0001
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFE
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFC
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
0000
0001
0001
0000
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0002
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0002
0002
0002
0002
0001
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFD
FFFD
FFFF
0001
0002
0001
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0001
0000
0001
0001
0002
0001
0001
0000
0000
0001
0002
0002
0001
0000
0001
0001
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0001
0001
0001
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
0000
0001
0000
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0002
0002
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0001
0002
0001
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFC
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0002
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
0000
0001
0001
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0001
0002
0001
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFE
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0000
0001
0001
0002
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
0000
0000
0001
0001
0000
FFFF
0000
0001
0002
0002
0001
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0002
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0001
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0001
0002
0001
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0001
0003
0003
0001
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0001
0002
0002
0001
0000
0001
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0002
0002
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0002
0004
0004
0001
FFFF
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0002
0001
0001
0001
0001
0001
0002
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0002
0003
0003
0001
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0002
0001
0001
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0001
0002
0002
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0001
0003
0003
0002
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0002
0001
0000
0000
0000
0001
0000
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFD
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0001
0001
0001
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0000
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0001
0003
0003
0002
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0002
0001
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0002
0002
0001
0002
0002
0002
0001
0000
0000
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0002
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0001
0001
0001
0000
0001
0001
0002
0002
0001
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
FFFF
0000
0001
0001
0001
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0001
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0002
0003
0002
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0002
0002
0001
0001
0000
0001
0001
0001
0001
0000
0001
0001
0000
0000
0001
0001
0002
0002
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0002
0002
0002
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0002
0003
0001
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0002
0001
0001
0001
0002
0002
0001
0001
0002
0002
0001
0000
0000
0001
0002
0002
0002
0002
0002
0002
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0002
0002
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0002
0002
0002
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFD
FFFD
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0001
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
0000
0002
0003
0001
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0000
0001
0001
0002
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0001
0002
0003
0002
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0001
FFFF
FFFE
FFFE
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0002
0002
0001
0000
0001
0002
0001
0001
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0002
0003
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0002
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0003
0002
0001
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0002
0001
0001
0001
0001
0002
0001
0001
0001
0002
0002
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0001
0001
0000
0000
0000
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0001
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0000
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
0000
0002
0002
0002
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
FFFF
FFFE
FFFF
0000
0001
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0001
0003
0003
0001
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0002
0002
0002
0002
0001
0001
0001
0002
0002
0002
0001
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0000
0001
0002
0002
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0002
0002
0001
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0002
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0002
0002
0002
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0000
0000
0000
0001
0001
0001
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0001
0001
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0001
0002
0002
0001
0000
0001
0002
0002
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0002
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0002
0001
0001
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
FFFF
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0001
0001
0000
0000
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0002
0002
0002
0002
0002
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0002
0004
0003
0001
0000
0000
0000
FFFF
FFFE
FFFF
0000
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0001
0001
0001
0001
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0002
0001
0000
0000
0001
0001
0001
0002
0002
0002
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0002
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
FFFF
FFFF
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFD
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0001
0001
0001
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0002
0003
0003
0001
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFF
FFFE
FFFE
FFFD
FFFD
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFE
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0001
0001
0001
0000
0000
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0002
0001
0001
0000
0001
0001
0001
0000
0000
0001
0001
0001
0000
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0000
0001
0001
0001
0001
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0001
0001
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0001
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0001
0001
0000
0000
0000
0001
0001
0000
FFFF
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
FFFF
FFFF
0000
0000
0000
0001
0001
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFE
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFE
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0001
0000
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
FFFF
0000
0000
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0001
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFD
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0000
0000
0001
0000
0000
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFF
FFFF
FFFF
0000
0000
0000
0000
0000
0000
FFFF
FFFF
0000
0000
0000
0000
0000
0000
0000
0000
0000
FFFF
0000
FFFF
FFFF
FFFF
FFFE
FFFE
FFFE
FFFD
FFFD
FFFD
FFFE
FFFE
FFFE
FFFE
FFFE
FFFF
FFFF
0000
FFFF
FFFF
FFFE
FFFE
FFFF
0000
0000
0000
0000
0000
0000
0000
FFFE
FFFE
FFFF
0001
0001
FFFF
FFFE
FFFD
FFFE
FFFD
FFFD
FFFD
FFFF
0000
FFFF
FFFE
FFFD
FFFE
0000
0000
0000
0000
0000
0001
0000
FFFF
FFFF
0000
0000
FFFF
FFFF
FFFF
0000
0000
0000
0001
0001
0001
0001
0001
0000
FFFF
FFFE
FFFE
FFFF
0000
0000
FFFF
0000
0001
0001
0000
FFFE
FFFE
FFFF
0000
0000
0000
0001
0003
0004
0003
0002
0003
0003
0002
0000
0000
0001
0002
0002
0001
0001
0002
0002
0001
0000
FFFF
FFFF
FFFF
FFFF
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0002
0001
0000
0000
0001
0001
0001
0001
0001
0002
0003
0001
FFFE
FFFE
0001
0002
0002
FFFF
FFFE
FFFE
FFFE
FFFD
FFFC
FFFE
0001
0002
0000
FFFE
FFFE
0000
0000
FFFF
FFFF
0000
0001
0001
FFFF
FFFE
FFFF
0001
0001
0001
0001
0001
0001
FFFF
FFFF
FFFF
FFFF
FFFE
FFFC
FFFB
FFFC
FFFC
FFFC
FFFC
FFFC
FFFC
FFFD
FFFC
FFFD
FFFD
FFFE
FFFE
FFFE
FFFF
0001
0001
0001
0000
0000
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0001
0000
0000
0000
0000
0000
0000
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
FFFF
0000
0001
0002
0002
0002
0001
0001
0001
0002
0002
0003
0004
0004
0004
0003
0002
0002
0002
0002
0002
0001
0001
0001
0001
0001
0000
FFFF
0000
0001
0000
FFFE
FFFE
FFFF
0000
0000
FFFF
FFFE
FFFF
FFFF
FFFF
FFFF
0000
0001
0001
0000
FFFF
FFFE
FFFE
FFFE
0000
0002
0002
0000
FFFE
FFFF
0001
0001
FFFF
FFFD
FFFC
FFFD
FFFD
FFFC
FFFB
FFFC
FFFC
FFFD
FFFC
FFFC
FFFD
FFFE
FFFE
0000
0000
0000
0000
FFFF
FFFE
FFFD
FFFD
FFFE
FFFF
0000
FFFE
FFFD
FFFD
FFFF
0000
0000
FFFE
FFFC
FFFB
FFFC
FFFE
0000
0000
FFFF
FFFD
FFFE
0000
0002
0003
0003
0004
0003
0001
0001
0004
0008
0008
0005
0002
0004
0007
0007
0004
0001
0000
0001
0002
0001
0001
0001
0000
0001
0002
0002
0001
0000
0001
0003
0004
0004
0002
0002
0004
0006
0006
0006
0006
0007
0006
0004
0001
0000
0000
0001
0001
0000
FFFE
FFFD
FFFF
FFFF
FFFE
FFFD
FFFD
FFFD
FFFC
FFFC
FFFC
FFFE
FFFD
FFFA
FFF7
FFF8
FFFC
FFFD
FFFA
FFF8
FFFB
0000
0002
0000
FFFC
FFFA
FFFB
FFFE
0002
0005
0004
FFFE
FFF7
FFF3
FFF5
FFF9
FFFD
FFFE
FFFA
FFF2
FFEC
FFED
FFF6
FFFF
0001
FFFE
FFFD
FFFE
FFFC
FFF8
FFF7
FFFD
0006
0006
FFFD
FFF4
FFF4
FFFB
0002
0004
0004
0003
0001
FFFF
0000
0005
0007
0005
0001
0001
0004
0002
FFFC
FFF9
FFFF
000A
0011
000D
0003
FFF9
FFF7
FFFE
000B
0012
0010
0006
FFFF
0000
0007
000C
000B
0007
0004
0005
0006
0004
FFFF
FFFA
FFFC
0003
0009
0007
FFFE
FFF9
FFFD
0006
0008
0002
FFFC
FFFC
0003
0007
0002
FFF8
FFF4
FFFA
0003
0006
0001
FFFD
0000
0009
000D
0006
FFFB
FFF9
0002
000F
0015
0012
0009
FFFF
FFF9
FFFC
0007
0012
0011
0008
FFFF
FFFF
0001
FFFF
FFFC
FFFE
0005
0008
0006
0003
0003
0005
0005
0008
000F
0013
000A
FFFB
FFF4
FFFC
0009
000C
0004
0000
0003
0008
0007
0007
0010
001C
001F
0016
0009
0000
FFFE
0001
0005
0006
0001
FFF6
FFED
FFED
FFF4
FFFC
0000
0003
0004
0003
0002
0004
000A
000A
0002
FFFA
FFFB
0000
0003
FFFF
FFFB
FFFC
FFFE
0000
0001
0003
0005
0005
0004
0005
0008
0007
0001
FFFB
FFF8
FFF8
FFF7
FFF9
FFFC
FFFA
FFF0
FFE7
FFE9
FFF6
0001
0001
FFFC
FFFC
0000
0003
0002
0004
000B
0010
000F
0009
0006
0006
0007
0009
000E
0010
000D
0009
000B
000D
0006
FFFB
FFF8
0002
000E
000B
FFFD
FFF5
FFFB
0006
000C
000C
000A
0005
FFFE
FFFF
000D
001B
0019
0008
FFF9
FFF9
0003
000C
0012
0016
0013
0006
FFF9
FFFC
000A
0011
0005
FFF7
FFF8
0005
000B
0005
FFFC
FFF6
FFF0
FFE9
FFE9
FFF5
0001
FFFF
FFF1
FFE8
FFEF
FFFE
0008
0009
0005
FFFE
FFF6
FFF1
FFF3
FFF5
FFF3
FFF2
FFF2
FFF1
FFEB
FFE6
FFEB
FFF5
FFF8
FFF3
FFF1
FFF9
0001
FFFA
FFEC
FFE8
FFF0
FFF4
FFF0
FFF0
FFFA
FFFF
FFF3
FFE4
FFE7
FFF7
FFFE
FFF6
FFF0
FFF6
FFFB
FFF2
FFE6
FFEE
0008
0016
000D
0003
0009
0013
000D
FFFC
FFF7
0001
000A
000A
0009
000E
0011
0009
0000
FFFF
0008
000E
000C
0007
0004
0001
FFFE
FFFE
0002
FFFF
FFF8
FFFB
0007
000A
0000
FFFE
000C
0017
000D
0002
0011
002B
0028
0006
FFF9
001A
0036
0016
FFE1
FFED
0029
0031
FFED
FFCC
0015
0058
000A
FF83
FFAF
008E
0098
FE45
FA20
F690
F563
F614
F6CC
F6A0
F62A
F635
F69A
F6B7
F677
F656
F68B
F6C0
F6AA
F680
F693
F6CC
F6D4
F6A8
F69A
F6C9
F6F1
F6DB
F6B3
F6C0
F6F3
F6FD
F6D2
F6BA
F6E1
F710
F700
F6D0
F6D8
F71D
F742
F716
F6EA
F712
F75D
F753
F6FE
F6F6
F77B
F7E1
F768
F69B
F732
FA31
FE6A
016F
0201
0121
009D
0103
017F
0158
00E2
00D3
012C
0158
011D
00E1
00FD
0133
0125
00EF
00F1
012B
0143
0115
00F0
0113
0149
013E
0107
0101
0139
0153
0124
00F9
011A
0153
0141
00FB
00F2
0138
0158
010A
00B7
00E5
0157
0150
00C1
0091
014A
01E7
009D
FD05
F8EC
F69B
F69B
F785
F7D4
F76F
F72D
F772
F7C8
F7B6
F772
F772
F7B8
F7DA
F7B2
F788
F7A0
F7D2
F7D7
F7B4
F7AD
F7D2
F7E9
F7D2
F7B6
F7C5
F7E2
F7D8
F7B6
F7BA
F7EA
F7FE
F7D8
F7BC
F7E9
F82B
F822
F7E2
F7DE
F836
F870
F830
F7DF
F821
F8BD
F8BC
F7EA
F7AF
F9AF
FDB2
017B
0307
0280
01AF
01C8
025C
0279
020E
01CA
01FE
023E
0221
01DC
01DA
0213
0223
01F1
01CC
01F1
0228
0223
01F3
01E3
0205
021B
0202
01EA
01FF
0223
021D
01F9
01F4
0215
021F
01F7
01DB
01FC
0227
0208
01BB
01B7
0214
023F
01D3
0156
01A2
0276
0232
FF92
FB69
F819
F733
F802
F8AD
F861
F7DB
F7F8
F881
F8AE
F858
F815
F846
F891
F888
F84C
F850
F89A
F8C3
F89A
F86E
F883
F8AC
F8A1
F87D
F890
F8D2
F8E4
F8AB
F881
F8AE
F8EF
F8DC
F892
F88B
F8DF
F914
F8DF
F8A6
F8DE
F946
F93E
F8CD
F8B5
F941
F9A3
F90A
F83A
F91E
FC8A
00DF
038F
03B7
02BB
025C
02D9
033B
02FA
0291
029B
02ED
02FC
02BA
029A
02CC
02FC
02DB
029C
029A
02D0
02E8
02C5
02AA
02C4
02E3
02CC
029F
02A9
02E7
0304
02D7
02A3
02AA
02CE
02C5
0297
0293
02C3
02D2
0294
0262
0291
02DB
02B6
023D
0242
030C
0370
01CC
FE0A
FA1B
F821
F85D
F940
F967
F8E9
F8AE
F904
F960
F949
F900
F8FB
F933
F946
F91D
F909
F93A
F974
F96D
F93A
F92B
F950
F96A
F956
F93D
F94A
F963
F959
F939
F93D
F96F
F997
F991
F983
F998
F9B7
F9AA
F982
F983
F9B2
F9C2
F991
F978
F9CB
FA2B
F9E4
F91D
F938
FB80
FF7D
0315
0486
0409
033A
0334
03A8
03C8
0374
0337
035C
0392
0381
034F
0353
0387
0395
0363
0339
0353
0389
0390
0365
0342
0343
0348
0339
0336
0358
037A
036E
0346
033E
0362
0376
0357
032E
0330
0348
0341
0328
033C
0376
0371
030D
02D5
0355
0404
035F
0083
FC74
F964
F896
F94F
F9EE
F9BB
F94C
F959
F9C5
F9F6
F9C4
F996
F9B8
F9F2
F9F1
F9C3
F9B8
F9E3
FA09
FA01
F9EA
F9EF
FA01
F9FE
F9F1
FA00
FA25
FA2D
FA07
F9E5
F9F6
FA1B
FA1E
F9FF
F9F6
FA14
FA2E
FA26
FA1D
FA34
FA44
FA17
F9DA
F9F7
FA63
FA77
F9E1
F980
FAD0
FE33
0229
0499
04CE
03F4
038A
03E1
0439
0410
03BB
03BD
040B
042F
03FE
03C9
03D2
03F8
03F9
03DB
03D5
03EF
0400
03F2
03E0
03E5
03EB
03DC
03D0
03E9
0411
040B
03D0
03A5
03BB
03EE
03FC
03E8
03E6
03FD
03F7
03C7
03B3
03E5
0411
03D6
0377
03A7
046B
0487
0296
FECA
FB10
F94F
F99A
FA70
FA8D
FA0E
F9C5
F9FF
FA49
FA3E
FA0E
FA11
FA42
FA56
FA3F
FA37
FA60
FA89
FA7D
FA4C
FA2C
FA26
FA25
FA2A
FA51
FA90
FAAB
FA88
FA5B
FA65
FA96
FAA3
FA7E
FA67
FA89
FAB3
FAAB
FA91
FAAA
FAE8
FAED
FAAD
FA9C
FB01
FB5B
FAF6
FA2B
FA81
FD1A
0129
0477
0586
04E0
0429
0444
04BB
04CF
0481
0452
0470
048B
046C
0446
0458
0485
0488
0462
0450
046D
048B
0487
047C
0488
0490
046D
043A
0436
0464
047B
0455
042C
0446
0483
0489
044B
041D
0430
043F
040B
03CE
03F0
044F
0450
03D0
038C
0423
04D5
03F2
00C4
FCB3
FA04
F9A5
FA7D
FAF7
FAAD
FA51
FA6C
FAB7
FABE
FA97
FA9F
FADF
FAFF
FADC
FAB3
FABF
FADB
FACB
FA9F
FA97
FABD
FAD6
FAC3
FAB4
FAD2
FAF5
FAEA
FACB
FAE2
FB2D
FB53
FB27
FAED
FAF8
FB28
FB24
FAF2
FAFC
FB62
FBA7
FB5D
FAE2
FAE9
FB6A
FB84
FAD8
FA7C
FC12
FFBD
03A5
05B4
059F
04D2
049D
04FA
0527
04E4
04A0
04AF
04D2
04BC
048F
04A3
04F2
0524
050C
04E3
04DD
04E4
04CB
04A5
04AA
04DB
04F9
04E7
04CE
04D1
04CF
04A4
0478
048E
04D1
04DD
0493
0452
0477
04CF
04D8
0489
045E
0499
04CA
047E
0418
0466
0542
0532
02E4
FEE7
FB65
FA08
FA79
FB23
FB16
FAB4
FAB5
FB15
FB46
FB0F
FACC
FAD4
FB07
FB1A
FB07
FB02
FB14
FB17
FB01
FB00
FB2E
FB60
FB63
FB44
FB32
FB3A
FB3A
FB2D
FB39
FB63
FB6E
FB30
FAE4
FAEB
FB42
FB7C
FB58
FB20
FB34
FB79
FB85
FB53
FB58
FBB7
FBD2
FB1D
FA50
FB11
FE33
0273
057F
062D
0561
04C5
0500
0577
057D
052F
0510
053C
0561
054C
0526
0522
052F
052B
0522
0531
0545
052E
04EF
04CA
04DF
0508
0511
050C
0526
0557
0561
0532
0507
0510
0526
050A
04D4
04D3
0513
053C
0516
04E9
0509
0541
0512
0492
048A
0555
05E9
04A1
0121
FD14
FAAC
FA8C
FB71
FBD6
FB74
FB07
FB10
FB4F
FB57
FB2B
FB16
FB28
FB38
FB38
FB4A
FB73
FB7F
FB57
FB33
FB51
FB97
FBB2
FB8D
FB68
FB6F
FB79
FB52
FB18
FB1C
FB65
FB9F
FB97
FB7B
FB89
FBAC
FBA9
FB8A
FB99
FBDD
FBF9
FBBD
FB8F
FBDC
FC50
FC15
FB27
FAE4
FCD1
00B7
048C
065C
0615
053C
0514
0589
05D1
059F
0551
053A
0543
053D
0539
0559
057E
056C
0532
051E
0551
058A
0587
055E
054E
055C
055A
053D
053A
056C
059A
0588
0553
0549
0573
0581
0546
04FD
04EF
050A
050D
0502
0533
0593
059F
051A
04A2
0500
05DB
0598
0307
FEF4
FB9D
FA85
FB25
FBDA
FBC1
FB49
FB2D
FB6D
FB8B
FB60
FB42
FB6C
FBAD
FBBC
FBA6
FBA6
FBC1
FBC5
FB9F
FB7B
FB7A
FB83
FB78
FB70
FB89
FBA9
FB9A
FB6A
FB63
FBA9
FBF9
FC09
FBF0
FBFB
FC2C
FC32
FBF1
FBC2
FBEB
FC20
FBE6
FB62
FB4C
FBE5
FC6E
FC1B
FB7A
FC3A
FF42
035F
0646
06D6
05FA
0555
057D
05DA
05D5
059A
059F
05E1
05FF
05D2
059C
0599
05B9
05D0
05E0
05F9
0608
05EF
05C2
05B3
05C4
05BF
0591
0570
0588
05A9
058C
054F
0553
05AC
05E8
05AF
054A
0542
058B
0592
052D
0504
0591
05FF
04B9
0151
FD5F
FB0C
FAEE
FBB2
FBE0
FB6A
FB34
FB9B
FC0A
FBE8
FB72
FB4C
FB9E
FBF8
FBFA
FBC1
FB95
FB85
FB7D
FB88
FBBB
FBF1
FBF3
FBCE
FBCC
FC06
FC35
FC1D
FBE8
FBE8
FC0E
FC00
FBB5
FB9B
FBF2
FC55
FC41
FBE0
FBD5
FC37
FC49
FBAA
FB61
FD09
00CE
04CB
06D0
0694
05A9
057B
05EE
061A
05C3
0589
05D7
0646
0646
05E9
05B3
05D6
0602
05F7
05D8
05D8
05DF
05C4
059B
059B
05B5
05A2
055B
0538
056E
05B1
05A0
0556
0543
057C
059B
0569
0542
0587
05EA
05CF
0557
0558
0609
062A
042F
0045
FC8B
FAFB
FB78
FC48
FC36
FBA4
FB80
FBDD
FC0D
FBC2
FB74
FB9B
FBFE
FC14
FBCC
FB8A
FB8A
FBA1
FBA4
FBB3
FBEC
FC1B
FC08
FBDC
FBF3
FC48
FC72
FC3A
FBF9
FC16
FC6F
FC8F
FC65
FC4F
FC75
FC76
FC14
FBBE
FBF7
FC6B
FC3C
FB73
FB91
FE01
0227
05AB
06D2
0629
057C
05AB
061D
0610
05BC
05CA
0641
067F
063A
05DE
05D9
0604
0601
05DC
05E9
0628
0638
05FA
05CA
05F5
063B
0631
05E1
05B6
05CA
05C2
0573
053A
056F
05C9
05C1
0568
0555
05B2
05E9
0592
0544
05C7
0693
05E3
02C1
FE88
FBB0
FB46
FC16
FC65
FBE4
FB80
FBCC
FC47
FC44
FBE6
FBC6
FC0A
FC46
FC35
FC13
FC1C
FC2F
FC0D
FBD6
FBDC
FC1E
FC43
FC1F
FBF0
FBF4
FC08
FBEA
FBBA
FBCA
FC15
FC39
FC13
FC06
FC5F
FCBA
FC7D
FBD7
FBA9
FC46
FCCF
FC61
FBAA
FC87
FFCC
03EF
067E
06AB
05D5
059F
0623
0662
05F5
0589
05BF
0645
0663
0603
05AF
05BA
05DE
05D2
05BC
05DA
060A
05FE
05CC
05CE
060F
0630
05F8
05B4
05BB
05E3
05C7
057C
057E
05E3
0618
05BE
0550
057D
0612
062E
059E
0553
05FA
068A
051C
0152
FD2E
FB17
FB62
FC58
FC73
FBDE
FBA4
FC13
FC85
FC75
FC24
FC09
FC20
FC1A
FBF3
FBED
FC12
FC1A
FBEA
FBCB
FBFF
FC5C
FC84
FC64
FC3B
FC29
FC0D
FBE1
FBE0
FC2D
FC78
FC61
FC07
FBED
FC3C
FC7E
FC4E
FBFE
FC22
FC95
FC87
FBCA
FB9A
FD7F
015F
0534
06FB
06A6
05D7
05DD
0677
06AA
0637
05CB
05F1
065A
066E
061F
05DD
05E5
05FD
05ED
05DC
0604
0647
0651
0612
05CD
05B4
05AF
0599
0588
059E
05CA
05E0
05E5
0603
0624
0602
05A5
0582
05D9
0638
060B
0594
05B3
067D
0685
043A
0002
FC39
FADD
FB97
FC7A
FC53
FBAE
FB92
FC10
FC66
FC34
FBE6
FBEC
FC21
FC28
FC08
FC0C
FC37
FC46
FC29
FC19
FC3A
FC5D
FC54
FC42
FC59
FC7D
FC6E
FC3A
FC3C
FC80
FC99
FC42
FBDE
FBFA
FC73
FCA1
FC4D
FC10
FC5E
FCB4
FC48
FB81
FC07
FEEC
031F
0644
070B
0649
05B1
05F4
0677
0680
0624
05E6
05F0
0602
05F2
05DD
05DF
05E0
05CC
05C3
05E4
060E
060B
05DF
05C7
05DB
05E8
05C8
05A9
05C7
0610
0631
0615
05FA
0607
0606
05C3
057C
0599
05F8
05FB
0578
0531
05D4
06A3
05D0
0285
FE38
FB69
FB23
FC2C
FCB4
FC4F
FBD5
FBE5
FC26
FC10
FBCD
FBE2
FC4E
FC8D
FC62
FC26
FC2E
FC4B
FC2E
FBF8
FC03
FC49
FC65
FC36
FC13
FC41
FC78
FC55
FBFA
FBE9
FC39
FC76
FC5C
FC46
FC89
FCC9
FC82
FBF8
FBFE
FCB0
FD09
FC54
FB9D
FCDE
008E
04B6
06E6
06BA
05D6
05BA
0641
0675
0614
05BD
05DF
062B
0633
060F
060C
061D
05F8
05AD
05A0
05F0
063C
062C
05EB
05D9
05FE
0607
05D3
05A2
05A6
05BC
05B3
05B1
05EF
0638
0621
05AE
056F
05B5
0605
05BF
0531
0556
0658
06C5
04EC
00F1
FD01
FB35
FB8E
FC62
FC67
FBE2
FBBF
FC29
FC7A
FC47
FBEC
FBE7
FC29
FC43
FC1B
FC04
FC2E
FC5D
FC4D
FC1B
FC16
FC4A
FC7E
FC91
FC97
FC9B
FC7D
FC39
FC0E
FC2F
FC6B
FC6F
FC4F
FC6F
FCD3
FCF3
FC85
FC12
FC44
FCD0
FCB4
FBD2
FBB4
FDFF
0242
0601
073C
066A
058F
05CF
0681
0695
060A
05B0
05E2
0636
0648
063D
0654
0666
0631
05E2
05DC
0617
0623
05DA
059C
05C3
0615
061F
05E4
05CF
0601
061D
05E9
05B9
05EE
0649
0642
05DF
05B7
0605
0633
05C4
053C
0582
0650
05FA
0344
FF22
FBF7
FB2F
FBFA
FC98
FC54
FBD7
FBD6
FC24
FC2C
FBE1
FBB0
FBCC
FBEE
FBE2
FBD9
FC11
FC5E
FC67
FC2B
FC0D
FC45
FC94
FCA7
FC8A
FC83
FC9D
FC9E
FC69
FC33
FC29
FC2C
FC0E
FBF2
FC1C
FC72
FC90
FC63
FC61
FCCA
FD16
FC9C
FBDC
FC78
FF70
039C
068E
0704
0609
057F
0601
06AA
06A7
0642
0635
068A
06A8
0654
0603
061D
0664
0666
0626
0602
0612
060D
05D3
05A9
05C9
05FE
05F9
05CF
05D4
060A
0614
05D2
05A3
05D3
061C
060C
05B8
059A
05C2
05B7
0550
0536
05EA
068F
0569
01ED
FDC7
FB57
FB4F
FC46
FC9E
FC28
FBCF
FC0E
FC6E
FC64
FC0E
FBE3
FBFD
FC15
FC0C
FC10
FC36
FC53
FC45
FC33
FC4B
FC72
FC6F
FC49
FC46
FC79
FCA4
FC96
FC7A
FC8D
FCAD
FC8F
FC42
FC2C
FC71
FCAC
FC81
FC43
FC85
FD1C
FD1F
FC3B
FBA9
FD27
00E5
04EC
06FC
06B8
05B8
058B
0633
06B5
068F
0631
061F
0642
0635
05F2
05CC
05E4
0602
05FD
05FA
0619
0630
060E
05D3
05CA
05F5
0605
05D5
05A2
05AC
05CA
05B1
0579
0584
05E0
0618
05E0
058E
0599
05D8
05C0
055E
0572
062E
065A
0465
006E
FC99
FAF5
FB72
FC4D
FC42
FBAE
FB90
FC08
FC67
FC4C
FC13
FC22
FC4E
FC3D
FC0D
FC1D
FC66
FC81
FC49
FC1A
FC43
FC8D
FC8A
FC3F
FC19
FC4D
FC91
FC96
FC71
FC62
FC66
FC57
FC4C
FC7D
FCCF
FCD9
FC86
FC54
FCA1
FCF5
FC92
FBC4
FC17
FEBA
02DE
0639
073A
066F
0597
05A9
0631
065E
061E
05FA
062C
065C
0633
05DE
05C1
05EC
0616
060C
05EB
05E3
05F0
05F2
05E5
05DF
05E1
05D3
05B1
0597
059C
05B2
05C0
05CB
05DE
05E1
05BB
0593
05A6
05DD
05C6
0544
04EF
0566
0627
05A3
02E2
FEE9
FBF5
FB43
FBF7
FC67
FC06
FB93
FBBA
FC23
FC23
FBC4
FBAA
FC14
FC84
FC7D
FC28
FC03
FC27
FC45
FC31
FC1B
FC2C
FC4C
FC53
FC50
FC66
FC80
FC75
FC54
FC55
FC71
FC61
FC16
FBF9
FC5B
FCEA
FD05
FCA1
FC5C
FC8E
FCB4
FC3E
FBC1
FCC4
FFF7
0405
06AF
0703
061F
05B6
063B
06D3
06B3
0613
05AB
05C0
05F8
05FA
05D3
05B9
05B8
05BD
05C9
05DE
05E0
05B3
057A
0578
05B3
05E3
05D2
05A8
05A7
05C0
05AE
0577
0579
05D2
060A
05AE
051D
0538
0612
0652
0473
009D
FCD0
FB02
FB4D
FC28
FC44
FBBB
FB6E
FBB7
FC1C
FC27
FC00
FC0A
FC46
FC5D
FC32
FC0E
FC32
FC74
FC88
FC68
FC4E
FC55
FC58
FC45
FC3F
FC59
FC66
FC3F
FC16
FC3C
FC8B
FC81
FC07
FBBE
FC26
FCC2
FC98
FBC5
FBE3
FE5E
0289
0600
070E
064E
059D
05E7
0680
067D
05F8
05B2
05ED
062C
0608
05B6
05A3
05CF
05E6
05CB
05AE
05B1
05B3
059F
0597
05B9
05D9
05BF
058C
0594
05E0
0603
05B7
0554
0565
05DB
0609
05A1
0543
05A8
064E
05A0
02B0
FE9A
FBA1
FAF7
FBB8
FC35
FBDB
FB6B
FB97
FC16
FC3B
FBFD
FBE1
FC1B
FC46
FC15
FBD9
FC02
FC6B
FC85
FC2D
FBE0
FC03
FC56
FC63
FC2D
FC14
FC34
FC43
FC1F
FC11
FC4F
FC86
FC57
FBFF
FC1C
FCA2
FCAE
FBD2
FB2E
FC8C
0046
047F
06E1
06E1
05F0
05A5
0626
0690
065F
05F1
05CA
05DE
05D6
05A8
0596
05B3
05C2
05A4
0591
05BB
05F8
05F5
05BD
05AB
05DE
0602
05CC
0577
0571
05B6
05CF
058C
0556
058D
05E5
05D0
0574
059C
066A
0693
048E
008E
FCB5
FB06
FB6D
FC32
FC1A
FB84
FB6C
FBF2
FC5B
FC34
FBE3
FBEA
FC2C
FC36
FBFD
FBE3
FC14
FC43
FC2D
FBFD
FC04
FC35
FC46
FC2F
FC34
FC6A
FC83
FC4D
FC14
FC37
FC84
FC77
FC10
FBF7
FC7C
FCE4
FC50
FB40
FB89
FE5D
02AA
05FA
06E2
0625
057A
059A
05F5
05E9
059D
0596
05DD
0605
05E0
05B6
05CB
05F6
05E7
05A3
057A
0599
05D0
05DC
05B9
058E
057A
057D
0597
05C6
05E6
05CA
0582
0560
058C
05C0
059A
0540
0559
061E
06A1
0570
022A
FE3C
FBB5
FB5B
FC1A
FC6B
FBEC
FB67
FB8B
FC17
FC5B
FC30
FC07
FC29
FC56
FC3C
FBFC
FBF2
FC21
FC35
FC0A
FBE7
FC10
FC5B
FC6B
FC3A
FC19
FC34
FC5A
FC59
FC4B
FC58
FC5E
FC2B
FBF4
FC1F
FC87
FC70
FB9B
FB2C
FCC7
009A
04BC
06E9
06B9
05B8
0572
05EA
0631
05E3
0589
05A1
05F0
05FC
05CB
05BD
05E3
05E4
059C
0560
057D
05C6
05D2
0598
0573
0595
05C4
05BF
05A3
05A9
05BF
05A3
055F
054E
0588
05AD
0577
054A
05BE
0686
0644
03E0
FFF6
FC89
FB25
FB80
FC1D
FC04
FB84
FB60
FBB5
FC04
FBFA
FBD7
FBEC
FC1A
FC14
FBE0
FBCF
FBFD
FC25
FC16
FBFD
FC19
FC49
FC43
FC0E
FC05
FC46
FC72
FC36
FBD5
FBCF
FC1E
FC38
FBF1
FBCF
FC37
FCA1
FC42
FB76
FBE4
FEAF
02DD
0610
06DF
0614
056E
05A7
061D
0615
05B6
0592
05BC
05D1
05A7
058E
05C1
0604
05FD
05C1
05AC
05D5
05ED
05C8
05A2
05BA
05E0
05BD
056A
0559
05A4
05D3
058C
052E
054A
05BA
05BE
052F
04F1
05B2
0681
056F
01DE
FD9C
FB29
FB2B
FC18
FC43
FBA1
FB41
FB9F
FC1C
FC14
FBBB
FBA9
FBF4
FC2C
FC14
FBE9
FBE4
FBE4
FBBF
FB9A
FBBF
FC1D
FC55
FC35
FBFB
FBEA
FBF3
FBE3
FBD2
FC02
FC61
FC79
FC1B
FBBE
FBEB
FC5E
FC41
FB74
FB3C
FD1D
0105
04F6
06E0
0698
05A9
0572
05DB
0606
05AF
0569
059E
05FD
0604
05C2
05A7
05CD
05DB
05A0
0569
0587
05C9
05C6
057D
0556
057D
05A8
058E
055C
0568
059D
05A2
056D
0566
05B7
05ED
05A2
0542
058E
064E
0607
037F
FF67
FBFB
FADA
FB87
FC49
FC28
FBA3
FB8F
FBEC
FC16
FBD4
FB97
FBBB
FC02
FC03
FBCC
FBBC
FBEB
FC07
FBE3
FBBB
FBCE
FBF6
FBE6
FBB5
FBC5
FC19
FC43
FC05
FBBE
FBDC
FC25
FC0C
FB99
FB7F
FC06
FC6E
FBF3
FB39
FC03
FF2A
034D
0611
0682
05C1
0567
05CD
062B
05F9
0597
0592
05D8
05EC
05B2
058D
05BB
05FE
05FE
05C8
05AE
05C7
05D0
05A0
056A
0573
05AB
05C4
05A1
0580
0592
05B8
05BF
05BB
05D3
05E7
05A5
052D
0529
05DE
0655
04FD
0175
FD59
FAE4
FAC1
FBA2
FBF8
FB92
FB52
FBA8
FC07
FBD9
FB61
FB51
FBC0
FC17
FBF2
FBA5
FBA7
FBE5
FBF4
FBBF
FB9D
FBBB
FBD8
FBBE
FBA5
FBD6
FC20
FC0E
FBA4
FB70
FBBD
FC1B
FC09
FBC2
FBE0
FC52
FC4B
FB97
FB7A
FD82
017E
0543
06D2
064B
056C
056D
05F3
0619
05C9
059D
05D1
05F6
05BC
057A
05A0
0602
0614
05BC
0572
0587
05BC
05B5
0587
0588
05BC
05C8
058B
055C
0581
05C0
05B8
0583
058F
05D4
05BC
0509
047C
04F4
05F6
05B6
0303
FEDD
FBAA
FAD4
FB90
FC20
FBD0
FB54
FB71
FBEE
FC0E
FBA8
FB4B
FB64
FBBA
FBD9
FBB3
FB98
FBB3
FBDE
FBF1
FBF7
FC01
FBF3
FBB9
FB87
FB9F
FBED
FC0D
FBD7
FB9D
FBB6
FBFD
FC0B
FBE2
FBF9
FC70
FCAB
FC1B
FB6E
FC48
FF72
0396
0654
06A2
05A7
0527
0592
0601
05CA
055E
056C
05D4
05EF
059D
056D
05AD
05EE
05C1
056C
057B
05D5
05DF
0572
0525
056D
05E7
05E8
057C
054C
058F
05BC
0576
052E
0566
05C0
057C
04CF
04D2
05DC
0675
04BE
00BF
FCB0
FABE
FAF3
FBAD
FBB9
FB5A
FB4E
FB9F
FBBF
FB81
FB53
FB8B
FBE4
FBE8
FB9B
FB6B
FB8D
FBBA
FBA9
FB84
FB9F
FBE6
FBFA
FBC2
FBA2
FBDF
FC35
FC30
FBDB
FBB2
FBDF
FBFB
FBBC
FB8B
FBE6
FC68
FC23
FB2A
FB20
FD8B
01CE
0576
06AF
05FA
053B
057B
0627
064B
05DF
058A
0596
05B4
05A5
0596
05BA
05EC
05E3
05A7
057F
058C
05A4
0598
0576
056D
057B
0572
054A
0532
0547
0562
0551
052F
0542
0581
0586
0523
04D3
0533
05DC
054F
027E
FE5D
FB42
FA92
FB70
FC0D
FBBF
FB57
FB8F
FC01
FBEF
FB79
FB5F
FBC5
FBF9
FB93
FB22
FB57
FBF1
FC29
FBD9
FB9D
FBD4
FC13
FBE3
FB7D
FB74
FBCC
FBFD
FBCD
FBA8
FBE1
FC1B
FBE3
FB85
FBB3
FC5A
FC87
FBC1
FB19
FC4B
FFBB
03BD
061F
0642
0568
0515
0584
05E7
05B8
0559
0558
05A6
05C6
0590
055E
0575
059D
0583
0547
0547
0584
059C
0567
053A
0558
0581
0561
0523
0528
0564
0567
051C
0505
0569
05C0
0560
04A6
04AA
0597
05EB
0403
002A
FC7C
FACD
FB0D
FBCE
FBF6
FB8C
FB2F
FB34
FB6D
FB9D
FBBF
FBDD
FBE4
FBBD
FB80
FB6E
FBA9
FC00
FC0A
FBAF
FB59
FB79
FBDE
FBF1
FB97
FB67
FBC7
FC3B
FC16
FB8B
FB7C
FC19
FC6F
FBC3
FB0D
FC31
FFAE
03B4
0604
0633
059A
0574
05BA
05D1
0592
055D
0568
0588
0584
056C
0566
0571
0571
0565
055E
0558
054A
053E
0546
0559
0565
0561
0542
0510
04F7
0525
056F
0562
04EA
04AA
0538
0605
0574
028E
FE65
FB4A
FA83
FB39
FBC1
FB84
FB28
FB43
FB96
FBA0
FB69
FB60
FBA1
FBD2
FBAC
FB69
FB6A
FBAC
FBD3
FBB2
FB89
FB9C
FBCC
FBC7
FB89
FB6F
FBBB
FC26
FC28
FBBE
FB84
FBE7
FC5F
FC0D
FB21
FB22
FD61
014B
04C1
0624
05C4
0525
0532
0598
05AA
056A
0553
0593
05CE
05B5
0566
0530
052C
0538
0537
053B
055B
0583
057B
053B
0505
0517
054F
054E
0506
04DC
051D
0572
0540
04A3
0486
055A
05F9
048A
00C5
FCAD
FA9B
FAE2
FBDB
FC04
FB71
FB13
FB42
FB85
FB82
FB76
FB9F
FBC4
FB95
FB48
FB4A
FB9D
FBD0
FBAD
FB7B
FB8F
FBD7
FBF7
FBC3
FB76
FB6A
FBAD
FBF0
FBEE
FBC3
FBCA
FC15
FC2F
FBAC
FB10
FBC6
FEAD
02C0
05B8
064D
056C
04E6
0550
05C9
058C
0503
0500
0580
05C0
0572
051D
053D
0584
0570
0521
0519
0562
0576
051C
04CE
050D
059D
05CD
0566
04F2
04F7
0540
0533
04BE
048D
051C
05D6
055B
02D6
FF01
FBC4
FA91
FB25
FBFD
FBF7
FB51
FAFB
FB4F
FBC1
FBB8
FB54
FB1F
FB46
FB77
FB71
FB5F
FB7F
FBAF
FBA3
FB64
FB45
FB68
FB8A
FB74
FB4F
FB64
FBA3
FBB0
FB77
FB62
FBBF
FC2A
FBED
FB22
FB13
FD0B
00C6
0468
0626
05EB
0521
0504
057A
05AB
054E
04F2
0518
0580
059F
0563
0537
055A
0593
059A
057D
0572
0579
0566
0541
0548
057E
058D
053E
04DB
04D8
0533
0565
0521
04C9
04FF
05BB
05F4
047C
013A
FD83
FB16
FAA1
FB4F
FBC7
FB82
FB15
FB30
FBB5
FBF7
FBBB
FB7A
FB9C
FBE1
FBD2
FB7D
FB57
FB83
FB9E
FB67
FB27
FB41
FB85
FB78
FB24
FB25
FBB3
FC26
FBD6
FB24
FB0F
FBC8
FC45
FBA8
FAA9
FB1E
FDFB
0217
053F
0641
05C4
0532
053C
0580
056C
0507
04D0
0508
0560
0568
0520
04EF
050A
0537
0533
0512
051C
0553
056E
0550
053B
0563
058A
054F
04D3
04A9
0504
055B
0526
04C2
0500
05CB
05C3
0394
FFAB
FC17
FA95
FB03
FBD2
FBDD
FB5B
FB1D
FB5C
FB98
FB71
FB2F
FB46
FBA6
FBD6
FB9E
FB4F
FB48
FB73
FB79
FB50
FB49
FB84
FBB0
FB84
FB3E
FB53
FBBF
FBF9
FBB2
FB55
FB75
FBE3
FBD3
FB12
FAB9
FC3D
FFC1
03A6
05F6
0621
0543
04CE
052A
05A9
059C
0524
04E7
0524
057B
057C
0539
0516
0532
054D
0534
050E
0515
0531
0524
0501
0515
055A
0562
04FE
04AC
04F1
0583
0592
04F2
0486
050F
05D5
051E
021D
FE13
FB29
FA61
FAF1
FB7B
FB70
FB33
FB3F
FB87
FBA2
FB64
FB0F
FAF9
FB23
FB48
FB3E
FB27
FB39
FB70
FB8F
FB7A
FB62
FB78
FB9E
FB93
FB66
FB6B
FBA9
FBBF
FB7E
FB55
FBAB
FC16
FBC5
FAE2
FAFC
FD7A
01B8
054B
066A
05A0
04D0
04FC
058B
058D
050D
04C7
050B
056C
0577
0549
053A
054B
053F
0516
0515
054D
0566
051E
04B3
04A3
04FB
053A
04FF
0495
0499
0518
0571
0528
04AA
04CD
058D
05A5
03C6
0025
FC89
FAAC
FAB5
FB5E
FB7C
FB11
FADB
FB31
FB99
FB84
FB0E
FAD5
FB25
FBA3
FBC7
FB8A
FB56
FB6A
FB8E
FB74
FB3C
FB42
FB8E
FBC2
FBA5
FB79
FB8E
FBBD
FBA8
FB66
FB78
FBF0
FC13
FB59
FAA2
FBB4
FF31
037B
061E
0643
053D
04C4
052D
0596
0569
050D
0515
0562
056B
051C
04EC
0526
057A
0576
0520
04E3
04F2
0511
04F6
04BC
04BE
050E
0551
0539
04F2
04E2
050B
0502
0493
0445
04BB
0590
0539
028E
FE63
FB13
FA3C
FB2B
FBE7
FB75
FAA4
FA9B
FB4B
FBB5
FB64
FAF9
FB18
FB7D
FB7A
FB08
FACF
FB2A
FBAC
FBC8
FB90
FB72
FB85
FB70
FB1A
FAF7
FB62
FBF9
FC0B
FB8D
FB32
FB78
FBEB
FBBF
FB10
FB28
FD41
0107
049D
0645
05ED
0505
04E1
0578
05D6
0578
04E1
04CD
0530
0560
0516
04C6
04DE
0526
0526
04EA
04EA
053C
055D
04FC
0486
04A0
052B
056E
0526
04E6
0526
0571
0518
0463
045E
0548
05C6
042C
0077
FC8D
FA6D
FA61
FB1C
FB5B
FB09
FAD5
FB24
FBA3
FBC9
FB7F
FB30
FB37
FB77
FB91
FB6F
FB5D
FB86
FBAE
FB89
FB34
FB16
FB46
FB6A
FB47
FB25
FB67
FBD7
FBDF
FB72
FB3A
FB96
FBE1
FB5D
FA9E
FB61
FE8E
02D4
05BC
061D
0514
047E
04F5
0599
0592
0513
04D4
0504
052D
04F6
049C
048B
04C3
04E9
04D3
04BF
04E8
0522
052A
0517
0535
0575
056D
04F8
0498
04CD
054B
053C
0478
03F4
049A
05D1
05BE
0338
FF2C
FBC6
FA69
FAAF
FB44
FB52
FB02
FAE3
FB2C
FB8F
FBAB
FB78
FB47
FB58
FB94
FBB0
FB8E
FB60
FB5C
FB75
FB78
FB5E
FB50
FB4D
FB27
FAEA
FAE9
FB3E
FB83
FB5D
FB17
FB3C
FBAB
FB97
FAC6
FA6F
FC2C
0005
0407
0619
05F6
0506
049C
04D2
050C
0505
04F9
051E
054B
053D
0503
04EB
0514
0545
053E
0517
0512
0535
053A
04F3
04A0
04AB
0511
0548
04F8
048C
04B0
0551
059E
053E
04E3
053C
059B
046A
0116
FD18
FA9E
FA62
FB34
FB95
FB42
FAF7
FB2B
FB88
FB8A
FB2B
FAD1
FACC
FB0F
FB52
FB63
FB4E
FB39
FB26
FAFA
FAC2
FAB9
FAF9
FB4A
FB67
FB58
FB5A
FB6C
FB3D
FACD
FAB6
FB62
FC28
FBF3
FAFE
FB26
FDDE
0229
0566
060B
050D
0465
04CC
0566
055C
04EB
04C6
04FF
051F
04F9
04E2
0515
055D
0568
052F
04EC
04D8
04F5
0518
0520
0518
0522
0537
052D
04FD
04DB
04F2
0512
04E6
0490
04A5
0542
0549
0357
FF92
FBF9
FA6A
FAC2
FB5F
FB34
FAB1
FAAF
FB26
FB67
FB2F
FAF1
FB0C
FB44
FB43
FB2A
FB48
FB81
FB73
FB16
FAD2
FAEA
FB23
FB23
FAEE
FAE5
FB3F
FBB0
FBB8
FB43
FADC
FB0C
FB98
FBB3
FB14
FABA
FC22
FF9E
039A
05FA
0615
051D
0490
04C1
0515
0524
0514
051E
052F
052F
052F
0541
0544
051A
04EA
04F5
0536
055B
0534
04F4
04E5
04FF
0505
04DE
04B4
04BA
04FA
053B
051F
049C
0448
04B3
0559
04B1
01C9
FDB4
FAC6
FA41
FB2B
FBAA
FB27
FA8C
FA9C
FAF8
FAFC
FAC4
FAC6
FAF9
FB07
FB05
FB46
FBA4
FB93
FB05
FAA7
FAF2
FB70
FB67
FAF6
FAE3
FB5C
FBB3
FB8B
FB68
FBA5
FBA8
FAFC
FAA8
FC5F
0037
0417
05DB
0585
04CB
04E3
056F
05A0
0572
0559
055A
0528
04D9
04CF
0514
054B
0540
0520
050E
04E9
04A3
047D
04A9
04E1
04C4
0486
04B0
052C
0536
048D
0417
04B5
05A1
04E9
01B5
FD88
FACB
FA61
FB17
FB61
FAF3
FA85
FA8E
FAD1
FAFA
FB0A
FB1D
FB20
FB0B
FB0A
FB3D
FB62
FB30
FAD8
FAE1
FB5A
FBB2
FB7D
FB14
FB11
FB66
FB85
FB4F
FB50
FBBF
FBE7
FB37
FAAD
FC26
FFFC
0419
060C
0599
04A1
04A6
0552
0582
0506
04A7
04D7
0523
0511
04D1
04C6
04DF
04DA
04CC
04EB
0513
04F7
04AD
0495
04B6
04BA
048A
0487
04DA
04FB
0480
0408
048E
059C
0530
020E
FD98
FA8E
FA20
FB0C
FB85
FB30
FADD
FB03
FB40
FB35
FB1E
FB3D
FB55
FB1E
FAD3
FADD
FB26
FB3E
FB17
FB11
FB4C
FB6B
FB2F
FAEA
FB07
FB5F
FB79
FB53
FB6B
FBCE
FBCA
FB0E
FAAF
FC49
FFF7
03D2
05BE
0585
04B0
0491
050D
054F
0519
04DC
04E5
04FB
04E4
04CB
04E9
0515
0504
04C0
049D
04B1
04C4
04C0
04D5
0507
050E
04CE
04A8
04E4
0516
04B2
0410
042E
0511
0506
026E
FE0B
FA9E
F9E8
FAE2
FB68
FAE4
FA71
FAD9
FB78
FB66
FACB
FA81
FAC5
FB0A
FAF7
FAD8
FAEF
FB04
FAF3
FB0F
FB7E
FBBC
FB58
FAC8
FAC9
FB3E
FB5B
FAF5
FAD4
FB64
FBD4
FB4E
FAC1
FC31
000A
0414
05DA
0553
046B
0475
0509
0549
052C
0528
0548
0541
0525
0546
058B
056B
04DB
048A
04DA
0533
04EC
0459
044E
04D8
0530
04F3
04AA
04D1
0501
04A8
0431
048F
057F
0530
0255
FE0D
FAF0
FA54
FB2D
FBA8
FB39
FAAE
FABC
FB25
FB4E
FB19
FADF
FACE
FACB
FABD
FAB5
FAB9
FAB9
FABB
FAE4
FB31
FB61
FB4B
FB25
FB35
FB5A
FB3F
FAFC
FB0D
FB86
FBB5
FB2A
FAC5
FC29
FFB5
03A0
05A5
0561
0478
0466
04F4
051C
04B5
047F
04D7
0536
0516
04C6
04D8
053F
056E
0544
052E
0551
0543
04D0
0475
049F
04F8
04F1
04A4
0499
04CE
04BB
045B
046F
0521
050A
0293
FE4A
FACE
F9FE
FB01
FBB9
FB63
FAF0
FB1F
FB7D
FB5D
FAFB
FAF5
FB38
FB22
FAA3
FA69
FAC7
FB31
FB21
FAE4
FB02
FB4E
FB4A
FB0F
FB20
FB73
FB6F
FAF3
FAB4
FB1D
FB6F
FAE2
FA56
FBC8
FFA6
03C2
0594
050D
0438
0475
0526
0528
0492
0458
04B9
04FD
04B3
0459
047C
04E2
0509
04FD
0518
0541
0513
04A6
0487
04DC
051B
04E2
049F
04D7
0534
04FB
045E
0467
0530
0519
0294
FE61
FB13
FA45
FB19
FBA8
FB51
FAE8
FB1F
FB8E
FB8D
FB2A
FAE4
FADA
FAD9
FAE4
FB22
FB6A
FB61
FB14
FAFA
FB3C
FB63
FB0F
FA9D
FAA5
FB03
FB12
FAC7
FAE3
FB9A
FBF2
FB27
FA50
FB88
FF50
038C
05AC
055A
046A
0467
050A
0541
04DC
0488
04A1
04CB
04B6
0493
04A8
04D9
04E9
04E4
04F5
0507
04E4
04A9
04AA
04DD
04DC
049B
0499
050E
0559
04DD
041C
0435
0517
0500
026F
FE3F
FB07
FA4C
FB19
FB88
FB10
FA96
FAC0
FB1D
FB13
FAD3
FAE4
FB3D
FB53
FB01
FAB8
FAC7
FAEE
FAEC
FAF2
FB35
FB75
FB5C
FB1F
FB2C
FB6C
FB5A
FAEF
FAD2
FB48
FB89
FAE5
FA55
FBCC
FFAC
03C7
05A0
051F
043D
0461
0508
0519
049D
046D
04CA
0515
04F2
04D3
0518
0562
053A
04E0
04D7
0506
04F0
0493
046A
0490
0492
0442
042B
04AF
052B
04CD
040C
0440
056B
057E
02B4
FE14
FA93
F9D8
FAC7
FB5F
FB1E
FAEF
FB4D
FB92
FB2E
FA94
FA82
FAE2
FB0F
FAE2
FAC7
FAF6
FB29
FB27
FB1F
FB3E
FB4D
FB18
FADD
FB02
FB64
FB7D
FB3A
FB18
FB47
FB34
FA8D
FA54
FC0C
FFC1
0388
0561
053E
04B3
04DA
054F
0542
04CE
04AD
0508
0548
050A
04B4
04C3
0512
0525
04ED
04C7
04CC
04A7
043B
03F3
0429
049E
04E8
0509
053B
054E
04EB
045F
047C
0538
0503
0260
FE0A
FA9C
F9CB
FAB4
FB55
FB09
FAAE
FADF
FB1A
FAD2
FA76
FABA
FB5E
FB7B
FAEB
FA84
FACC
FB37
FB24
FADF
FB0E
FB8C
FBAA
FB4E
FB05
FB0F
FB04
FAB1
FA9D
FB20
FB82
FAF7
FA57
FBAE
FF96
03F3
0619
05B8
04BB
04A4
051C
0526
04BD
049A
04EA
051E
04E6
04AB
04C0
04DC
04AC
0471
0485
04B1
0493
045B
0486
0500
052D
04DD
049E
04CE
04F0
047A
03F6
046A
0581
0548
0262
FDFC
FABD
F9F9
FAAB
FB26
FAFE
FADB
FB15
FB44
FB11
FAD0
FAED
FB3F
FB4F
FB14
FAEC
FB06
FB2B
FB34
FB3F
FB5F
FB64
FB28
FAE7
FAEF
FB1D
FB12
FAD9
FAEC
FB5F
FB83
FAE0
FA60
FBB5
FF55
037C
05CC
05AF
04AC
0465
04E9
0541
0504
04B3
04B8
04CE
0499
0450
0462
04BA
04DE
04B1
0499
04C5
04E0
04A7
0465
0476
04AF
04AE
0488
049A
04D0
04B5
0458
0476
0535
0532
02D0
FE87
FAE4
F9D8
FAB3
FB62
FB10
FA9C
FACE
FB36
FB16
FAA0
FA91
FAFA
FB30
FAEE
FABD
FAFB
FB3F
FB18
FAD8
FAFE
FB55
FB51
FB03
FB01
FB62
FB89
FB2A
FAD9
FB19
FB61
FAE7
FA4F
FB72
FEFE
032D
0590
05A3
04DB
048B
04A4
0493
0468
048D
04EB
04FB
04B2
0498
04EC
0536
050E
04BE
04B8
04D5
04B0
0466
046B
04B6
04C6
0479
0453
04A1
04D7
0463
03CD
042D
0552
055B
02CA
FE8F
FB35
FA3A
FAD3
FB5B
FB39
FAF8
FB07
FB23
FAFC
FACA
FAE2
FB22
FB30
FB07
FAF1
FB06
FB15
FB08
FB01
FB08
FAEE
FAB1
FAB4
FB30
FBB2
FB98
FB0D
FAF1
FB87
FBE0
FB2C
FA4E
FB45
FEC2
02EF
0545
0536
046B
0473
0518
0546
04CD
0474
04A3
04DD
04AA
0464
049C
051F
0539
04C1
0458
0476
04CB
04D9
04AB
048D
047A
044C
0434
0479
04DA
04C4
0457
046E
053B
054D
02FD
FEC1
FB24
FA0F
FACB
FB50
FAE2
FA6E
FABA
FB43
FB36
FAB8
FA89
FAD3
FB0A
FAF5
FB02
FB66
FBA6
FB5E
FAF2
FAE9
FB14
FAFF
FAD2
FB0F
FB8E
FB8F
FAF4
FAA2
FB28
FBA1
FAF1
F9EA
FAE6
FECB
0373
05E8
059F
0489
045B
04DE
050D
04C2
049C
04CB
04D7
049C
048E
04E1
0517
04CD
046F
0482
04CE
04C4
047E
048D
04EE
04FE
0489
0440
04A7
0523
04CF
040E
0430
054E
0581
0300
FE95
FAFA
F9DF
FA71
FAE7
FAAA
FA74
FAC6
FB29
FB08
FAA2
FAA0
FB0F
FB58
FB1F
FAB8
FA9F
FAD6
FB05
FB02
FB00
FB2F
FB60
FB3E
FACF
FA96
FAE8
FB56
FB22
FA64
FA70
FC9D
009C
0464
0608
058F
049D
0482
0507
0542
04F6
04AA
04BB
04E7
04DA
04B3
04B7
04CA
04A3
045B
0466
04DC
0532
04EA
0456
042F
0492
04D1
0474
0404
0462
055B
0567
0325
FF0F
FB4E
F9BD
FA3A
FB1D
FB24
FA8C
FA4C
FAAF
FB1B
FB06
FAB3
FAB2
FB0B
FB41
FB15
FADC
FAEB
FB16
FB0A
FAE0
FAFD
FB62
FB8B
FB31
FACB
FAF2
FB70
FB6A
FAB2
FA86
FC64
0032
03F9
05C0
0570
049A
048E
051B
054A
04D9
0476
04A7
050C
04F9
0480
0452
04AF
0507
04CE
0449
0420
046C
04A9
0490
0482
04D1
050E
04A3
03E2
03D2
04AC
050D
0355
FFA3
FBFB
FA43
FA7D
FB33
FB3B
FABC
FA7E
FABF
FB13
FB1B
FAF4
FAE2
FAE3
FACE
FAAB
FAB7
FB05
FB4D
FB44
FB01
FAE2
FB08
FB2D
FB13
FAFA
FB3C
FB9F
FB71
FAA0
FA5D
FC1E
FFE0
03BD
05A9
0568
0481
0462
04F8
0548
04ED
0474
0471
04BD
04D7
04A3
047B
0499
04CB
04D6
04D0
04E4
04F0
04A9
0428
03F1
0444
04AC
048D
040D
0404
04C5
053A
03C8
0032
FC3E
FA18
FA2C
FB03
FB22
FA95
FA51
FAAA
FAFA
FAC4
FA7C
FAC2
FB5B
FB76
FAE6
FA71
FAB3
FB3C
FB43
FAD3
FAB2
FB2C
FB9C
FB6A
FAF9
FB11
FB9B
FB9E
FAC0
FA3F
FBC9
FF77
036A
0595
05A4
04E2
049D
04EC
051C
04D5
047C
048A
04E3
050A
04CC
047D
0475
04A7
04C3
04B0
049F
04AE
04B1
0480
0448
044C
0470
045B
0417
0435
04E4
0533
03C0
005B
FC99
FA6F
FA4D
FAED
FAFE
FA82
FA52
FABC
FB28
FB0A
FAA6
FA95
FAE7
FB1E
FAFC
FAD5
FB02
FB54
FB5C
FB1A
FAF8
FB20
FB36
FAEF
FAA3
FADD
FB78
FBA3
FB00
FA87
FBBD
FEFE
02D3
0542
059F
04F2
0499
04EB
0543
051B
04AF
0483
04A8
04BE
0494
046B
048D
04D3
04DF
049F
046C
0488
04C5
04D4
04B5
04A5
04A6
0477
041F
041D
04B5
0517
03D9
008C
FC99
FA25
F9FA
FAE5
FB41
FAB6
FA36
FA78
FB15
FB43
FAF1
FABC
FAF0
FB26
FAF2
FA94
FA97
FB01
FB44
FB0F
FABA
FABD
FB03
FB18
FAF0
FAF8
FB52
FB76
FAFB
FA93
FBA9
FEC6
02A3
053B
05BA
0510
04A3
04D8
0511
04D8
047E
0487
04E1
050F
04E5
04BD
04DE
050A
04DC
046E
043D
0475
04B0
0488
0439
0445
04AC
04DA
0488
0446
04AA
052C
044D
0143
FD34
FA50
F9B6
FA86
FB22
FAF0
FA94
FAB5
FB14
FB14
FAA8
FA5D
FA86
FAD6
FAE5
FAC0
FABB
FAE2
FAFC
FAFC
FB19
FB5B
FB67
FB01
FA96
FAC5
FB6F
FBA1
FAD8
FA10
FB08
FE4D
025E
050A
0588
04ED
04AB
0509
0546
04EC
046D
046A
04CE
04F9
04AF
0463
048E
04FE
0522
04D6
048C
049B
04C6
04A7
045C
0462
04C5
04EB
0474
03F1
042F
04E1
0478
01D6
FDD8
FAC2
F9F7
FABA
FB51
FAFF
FA72
FA77
FAE3
FB05
FAB9
FA83
FAB3
FAF6
FAE6
FAAE
FABA
FB08
FB2A
FAF4
FAC7
FAF2
FB2B
FAFE
FA94
FA9A
FB3F
FBBB
FB4E
FA83
FAFF
FDB6
01A8
04AE
0586
04D7
042C
044B
04C3
04E5
04B2
049C
04C5
04D4
0495
0457
047E
04EC
051C
04DF
0496
04A3
04DA
04D0
0487
047C
04DA
0520
04CF
0440
043D
04B5
0457
01FA
FE2F
FB03
F9F5
FA93
FB42
FB25
FAB6
FAB5
FB11
FB2F
FAE5
FAB3
FAF0
FB4B
FB3F
FAD5
FA89
FA9D
FAD6
FAF6
FB15
FB56
FB77
FB20
FA83
FA54
FADB
FB68
FB22
FA61
FAB7
FD4E
015D
04AF
05C0
050F
0446
045A
04D8
04EC
048E
045A
048D
04BD
0495
045C
0489
04F9
0512
04A0
0431
0455
04DB
0516
04CE
0479
047A
048E
0455
0417
0473
0532
04FC
02A8
FEC9
FB69
FA1D
FA95
FB45
FB31
FAB2
FA92
FAE7
FB20
FAED
FAA6
FAB6
FAFE
FB14
FAE5
FACA
FAF3
FB1D
FB00
FACE
FAEE
FB4B
FB5B
FAEC
FA94
FAEE
FB9B
FB9B
FACD
FA9A
FC92
0070
040E
0585
0503
0436
043F
04C4
04F0
04B8
04B3
0508
052D
04C5
043A
0428
0487
04CA
04B4
048F
049B
04A7
047F
0463
04B2
052E
051E
0457
03B5
0421
0528
0513
02AF
FEBB
FB56
FA09
FA7C
FB31
FB2F
FABE
FA9B
FAE2
FB0D
FACE
FA8C
FAC6
FB4D
FB75
FB05
FA9C
FAD9
FB6F
FB80
FAD4
FA37
FA66
FB0C
FB48
FAEA
FAA4
FAE0
FB1A
FAD7
FAE4
FCB7
0068
0417
05BF
0556
047C
0467
04CB
04D7
0490
0488
04C7
04BD
044F
042A
04AC
0523
04BC
03E0
03C4
04B7
058B
052F
043A
0425
0533
05EA
0519
0399
0352
049B
0576
03B9
FF8F
FB70
F99E
FA21
FB3A
FB6F
FAD1
FA5E
FA9D
FB1C
FB2E
FACA
FA8E
FAE5
FB73
FB84
FAF6
FA66
FA74
FAFB
FB53
FB20
FAB4
FA90
FAD3
FB37
FB74
FB5F
FAE8
FA53
FA79
FC4A
FFB2
0340
054A
057B
04E8
04A8
04C2
04B2
0479
0493
04FB
04FC
0446
03A6
040D
0526
0591
04B8
03AD
03D3
0508
05D2
0550
0446
03ED
045B
04A9
0473
0454
04B1
04B7
0321
FFE5
FC87
FAA1
FA6B
FAE7
FB1C
FAE0
FA98
FA9C
FAF4
FB58
FB64
FAEF
FA5B
FA54
FB0F
FBDC
FBD0
FAE0
FA0A
FA3D
FB3C
FBED
FB9A
FAB7
FA44
FAAD
FB5A
FB6C
FAD0
FA94
FC09
FF5A
031B
055C
0578
049B
045A
04E8
0534
04AB
041E
048A
0579
0576
0423
02F3
035D
04E0
059D
04CD
03A8
03A3
048B
051A
04D1
0466
0469
0481
0453
045A
050B
0573
03DF
0011
FC12
FA1A
FA3C
FACE
FAB2
FA5D
FA8E
FAFC
FAEC
FA88
FAAF
FB84
FC05
FB6F
FA71
FA4F
FB31
FBFA
FBC8
FB00
FA98
FADB
FB42
FB53
FB2C
FB19
FB0D
FAD2
FA90
FAEA
FC7D
FF57
02B0
0532
05E1
0507
0417
0448
054F
05C7
04F6
03BE
0384
0470
054A
0511
0423
0396
03D8
0472
04D3
04DC
04A2
043C
03EB
0413
04AE
050F
04B3
0415
0415
0473
03AD
00D2
FD07
FA7C
FA00
FA62
FA4F
FA09
FA8F
FBB9
FC22
FB26
F9FE
FA34
FB9C
FC90
FC1B
FB03
FA8C
FAE2
FB48
FB5A
FB60
FB6F
FB1B
FA5C
FA0C
FAD9
FC0C
FC28
FAEC
FA06
FB57
FEDB
02BC
0533
05E6
057A
049A
03D1
03B4
047D
057E
059C
049B
0380
0369
0441
04FD
04EB
045A
03F3
03EC
0426
0494
050D
051E
047C
03B8
03CE
04CA
054D
03DA
008C
FD03
FABA
F9E8
FA02
FAA2
FB81
FBFC
FB86
FA81
FA0D
FAB2
FBAA
FBDB
FB36
FAA0
FAA8
FAFD
FB3D
FB85
FBE0
FBC8
FAE6
FA04
FA4F
FBA3
FC60
FB84
FA5D
FB45
FECB
02E9
0549
0594
050E
04AE
0469
042B
0459
0515
05A2
0536
0422
0387
03F1
04C6
0530
050B
049F
0417
03AB
03DD
04D2
05A7
0539
03CA
030D
0400
053A
0445
0094
FC55
FA02
F9E0
FA79
FACD
FB17
FB91
FBAF
FB00
FA30
FA4D
FB46
FBE8
FB6E
FA72
FA05
FA5D
FAE7
FB37
FB4C
FB27
FAC3
FA7D
FADD
FBB2
FBF5
FB26
FA75
FBC7
FF65
035D
058B
05B7
053E
0513
04F4
0479
040B
0447
04F6
0541
04D2
0439
0410
0452
04B1
0516
055D
051B
0436
037F
03ED
053A
05ED
0533
0410
03FD
049B
03D1
007E
FC3C
F9BE
F9CF
FAD4
FB1C
FABB
FABC
FB40
FB59
FA95
F9CD
FA03
FB07
FBC2
FB8C
FAC8
FA3C
FA56
FAFD
FBBA
FBEF
FB47
FA37
F9C1
FA55
FB2F
FB4B
FB08
FC0D
FF38
0331
05AC
05DA
04FB
048B
04A0
0479
040E
0427
050D
05E1
05B0
04AB
03D4
03C9
0455
0504
0581
057C
04C7
03D9
03AC
049B
05B2
05AA
049D
03D7
03D8
0349
00B1
FCBD
F9E2
F99F
FAEA
FBAF
FB44
FAB2
FAD9
FB44
FB15
FA67
FA1B
FAA1
FB80
FBFA
FBB5
FAD0
F9D4
F989
FA5E
FBB8
FC3B
FB48
F9E4
F9A7
FAC2
FBE9
FC5D
FD21
FF81
02DF
0517
051A
0431
042E
0512
0560
0479
0399
040F
055E
05E5
04FB
03AA
034D
0421
055B
0618
05F3
0505
03DC
0356
03F5
053B
0604
05B8
04B8
037F
01D4
FF5A
FC93
FA9E
FA02
FA30
FA76
FAD5
FB8C
FC2D
FBEE
FADC
FA0D
FA47
FB08
FB5D
FB27
FAFE
FB06
FAC7
FA3B
FA39
FB38
FC3E
FBE3
FA45
F91A
F994
FB01
FC2F
FD5F
FFC8
0354
0609
0647
04DD
0400
048B
053A
04C1
03B0
038C
049A
058B
0546
043C
03A5
0401
04CD
055F
0577
0518
045F
03C3
03F1
04FE
0606
0600
04CE
0315
013A
FF02
FC71
FA5F
F9C1
FA72
FB40
FB47
FACD
FA9C
FAE5
FB2A
FB11
FACC
FAB3
FADF
FB38
FB93
FBA4
FB1B
FA28
F9B4
FA79
FBE3
FC61
FB2A
F95F
F8EB
FA7D
FD0D
FF52
0112
02C1
045B
0542
0532
04B9
0482
0497
04A9
04BB
0508
056F
0572
04E1
042A
03CF
03DC
0418
047C
0507
0549
04BF
03C2
0383
049D
0610
063F
04BD
029B
00C6
FEF3
FC90
FA41
F974
FA72
FBB3
FBA7
FA8E
F9E9
FA61
FB0B
FAE2
FA39
FA27
FAFB
FBD6
FBDC
FB2F
FA86
FA51
FA91
FB2C
FBDC
FC03
FB27
F9C6
F931
FA54
FCC3
FF50
015F
032F
04F0
0618
0609
0508
041F
041A
04D1
0584
0599
050F
0461
0429
0493
0519
04F6
0423
039C
0442
0584
05CF
048F
0335
0398
058F
06DB
05B1
029C
FF90
FD87
FBEF
FA45
F938
F9A0
FAF7
FBB4
FB29
FA42
FA2C
FAD8
FB44
FAF0
FA6A
FA66
FAD3
FB24
FB18
FAE1
FAB5
FAA5
FAC6
FB20
FB5C
FAFE
FA1C
F9A3
FA86
FCC7
FF87
0207
041F
05B6
0652
05AB
0474
03E8
0483
057F
05C8
0532
0478
043F
0486
04ED
052D
0520
04BB
0449
0452
04F0
0567
04FB
040F
03EC
0510
0634
057E
02A8
FF50
FD10
FBE2
FACF
F9A9
F954
FA4A
FB9B
FBD5
FAB2
F966
F940
FA55
FB9B
FC05
FB65
FA69
F9FC
FA76
FB42
FB76
FAE7
FA6B
FAC8
FB88
FB77
FA58
F997
FABA
FD88
0047
01ED
0320
04CB
0664
068B
0521
03CF
0412
056F
0630
0594
0482
041B
0457
0485
0480
04B1
052A
0563
050E
048C
045B
0473
048B
04B5
0527
0572
049B
0244
FF55
FD0B
FBB4
FABA
F9D2
F975
FA11
FB29
FBB6
FB3B
FA3C
F99F
F9E8
FAEF
FC01
FC3F
FB51
F9F5
F982
FA70
FBAD
FBDB
FB08
FA86
FAFB
FB68
FAB6
F9AE
FA66
FD8F
0152
036E
03D1
0432
0569
064B
058F
03DD
0333
045B
0600
0667
056A
044A
0405
0471
04DD
04EC
04B0
0466
044A
0470
04A5
0497
045B
0481
0543
05BE
049C
01AA
FE4F
FC17
FB28
FA9C
FA0C
F9FC
FABC
FB93
FB94
FAD3
FA3C
FA45
FA7F
FA84
FAA2
FB23
FB8C
FB45
FAAF
FAC5
FB9A
FC06
FB41
FA2A
FA33
FB47
FBD2
FB22
FAC4
FCB8
00B7
044B
058D
050D
04A0
050A
057F
0532
0483
045F
04FB
05A7
05AE
04FF
0423
03CD
0451
0533
0571
0497
037B
036A
047F
055F
04F2
03F8
0402
04FF
04E1
022C
FE1D
FB55
FAC7
FAFB
FA71
F9A4
F9F2
FB40
FBE3
FAF4
F99C
F980
FAA2
FB9B
FB93
FB0B
FAC8
FACA
FAC5
FAE4
FB7A
FC2A
FC26
FB59
FA9F
FA9A
FAEB
FB14
FB9C
FD8F
00E0
0411
05AC
05AE
0531
0501
050B
04F9
04CC
04B0
04BF
050C
0590
05CD
0518
03A8
02E5
03E3
05B3
0620
0469
027C
02A7
04A4
05F6
0548
0402
03EB
043D
028A
FE58
FA49
F919
FA5F
FB5D
FA9C
F976
F9CE
FB61
FC3C
FB59
F9C3
F927
FA02
FB76
FC5B
FC29
FB30
FA49
FA45
FB2A
FC13
FC15
FB51
FAB6
FAB9
FAED
FB1F
FC25
FECE
0258
04DC
056D
0515
0544
05E8
05D4
04C4
03E9
0432
04FB
0528
04C3
04AA
04F3
04BF
03DD
0375
0469
05B0
0579
03C0
029E
0383
0542
05AB
0470
032B
02AE
01AA
FEB2
FAB7
F865
F903
FAFC
FBD4
FAE7
F9AE
F9AB
FAD9
FC02
FC1B
FB28
FA27
FA27
FB34
FC28
FBD8
FA93
F9FA
FB09
FCA0
FCD3
FB70
FA4F
FAC4
FBE1
FC1B
FBFC
FDB9
01EF
0613
0726
0551
039F
0426
05C7
0635
0513
0401
0415
04A6
04AF
0459
0461
04B7
049F
0403
03B6
0425
049B
044A
0395
0381
0437
04D2
0494
03A9
0276
00C3
FE32
FB47
F948
F8FA
F9E1
FAEF
FB79
FB60
FAC8
FA26
FA2E
FB12
FC01
FBF3
FB08
FA87
FB27
FC08
FBE8
FB04
FAD4
FBCD
FC93
FBEC
FAAD
FAA6
FC06
FD1E
FD06
FD55
0023
04CF
0813
07AD
04F2
0319
039F
0537
05EC
0551
0457
03D2
03CF
040C
0464
04AC
04AF
0476
0448
0438
0404
03A1
037E
03EA
0479
0483
040C
038C
02DC
0108
FDB8
FA4D
F8C2
F97C
FADD
FB4C
FAE2
FAB6
FB0E
FB32
FAD6
FAA1
FB17
FB9C
FB54
FA8D
FA73
FB5F
FC42
FC25
FB80
FB6B
FBEA
FBEC
FAFF
FA29
FAA4
FC60
FE54
0003
01E2
042A
0603
065E
054F
0400
0374
03D0
04A2
0566
05A0
0509
03F2
034A
03B6
04BF
0544
04CA
03F0
037B
037E
03B8
0439
0509
055C
040C
011B
FE1E
FC99
FC3C
FB7F
F9E4
F8CA
F992
FB9C
FCD6
FC1A
FA5D
F964
F9E6
FB33
FC40
FC77
FBCA
FAA1
F9D9
FA49
FBCE
FD13
FCCB
FB1B
F98C
F998
FB86
FE8A
018E
03C5
04D3
04F8
04F0
0545
05A6
054E
0439
0377
03F0
0524
05B2
0509
0408
03CC
0453
04BA
048C
0434
0426
0435
041E
042F
04CA
056A
04C8
0247
FEC7
FBD9
FA46
F9BB
F9A9
F9F9
FAB7
FB7B
FBAB
FB29
FA86
FA66
FAE6
FB9A
FBEC
FB89
FAA6
F9F3
FA26
FB42
FC67
FC8C
FB87
FA31
F994
FA20
FBBD
FE26
00EB
0344
0487
04DD
0526
05D8
0643
0573
03B8
02B5
0393
0584
0689
05A7
03DF
02FA
03A6
050D
05E9
05A4
0488
035A
02F4
03D7
0596
06B5
05A2
022C
FDF1
FB17
FA82
FB38
FB8E
FAD2
F9D1
F9C6
FAF2
FC3E
FC60
FB35
F9F8
F9ED
FB06
FBFC
FBCB
FAC8
FA24
FA85
FB6A
FBF0
FBC2
FB2F
FA9C
FA5C
FAF5
FCFC
0046
038B
0553
055C
04BE
0493
04CD
04A7
03F6
038F
042B
0553
05C8
04F9
03B9
0351
041F
0543
059F
04EE
03E0
0359
03B4
04A7
0592
05C0
049A
01FA
FE8A
FBA0
FA60
FAC2
FB88
FB7B
FAA6
FA32
FAE9
FC25
FC78
FB5F
F9F0
F9AC
FAD6
FC34
FC78
FB8D
FA6F
FA0F
FA93
FB80
FC32
FC1B
FB15
F9D3
F9D5
FC50
00C2
04E9
0687
0570
039A
0322
0449
058B
0580
0459
0379
03CA
04CF
055A
04E9
0416
03C7
0432
04CB
0502
04CB
047B
0456
046F
04C5
051B
04C4
02F6
FFAC
FC25
FA0E
F9FC
FAE9
FB53
FAD7
FA56
FAA7
FB73
FBBD
FB32
FA9C
FAD2
FBA4
FC0D
FB77
FA6D
F9F7
FA76
FB55
FBC4
FB7D
FAD0
FA38
FA21
FAF9
FD17
003E
0369
0551
057F
04C0
045A
04C8
0560
053E
0464
03B6
03E4
0498
04ED
048E
0413
0438
04F6
0594
0585
04EC
044A
03FE
0425
04B1
0545
0506
030B
FF6B
FBA2
F990
F9CB
FB21
FBD6
FB50
FA6A
FA40
FAF5
FBBC
FBE2
FB82
FB2A
FB20
FB2A
FAFD
FAA6
FA73
FA8B
FACC
FAFF
FB0F
FAFD
FACC
FAAA
FB2A
FCFD
0031
03B6
05F2
0614
04DB
03D8
03EE
04AB
0512
04CA
0456
043A
045B
0450
041B
042E
04BC
054F
0548
04A6
040A
0404
048E
052F
057C
0534
040E
01CD
FEBC
FBD8
FA39
FA2C
FAF6
FB90
FB8F
FB49
FB31
FB45
FB30
FAD6
FA92
FAC4
FB54
FBBB
FB97
FB12
FAB2
FAC9
FB31
FB84
FB7C
FB1A
FA9B
FA74
FB4B
FD91
00EA
0410
05A5
0553
0417
0351
038B
0441
04B2
04B2
0497
0498
0496
0473
045C
0488
04CB
04BB
043A
03B8
03B8
043D
04C7
04EE
04B9
0453
0387
01D9
FF2F
FC49
FA52
F9F3
FACE
FBEA
FC7B
FC54
FBB4
FAF7
FA7A
FA96
FB55
FC34
FC5E
FB7B
FA35
F9B6
FA7F
FBDD
FCA0
FC42
FB45
FA7D
FA51
FACB
FC0E
FE4A
0129
03AC
04E8
04DD
045E
041F
041E
03FB
03B8
03B7
0423
0491
0480
0403
03B1
03F5
0495
04FC
04D9
045C
03E9
03C0
03EE
0467
04F6
0510
0405
0193
FE5B
FBA2
FA65
FA91
FB36
FB7E
FB66
FB6F
FBC3
FBF3
FBA3
FB2E
FB45
FBF2
FC5F
FBD5
FAC3
FA52
FB04
FC0F
FC55
FBA5
FAC9
FA74
FAA5
FB2B
FC4C
FE70
0141
03A9
04E4
0530
053D
0528
0483
0359
029D
0331
04B2
05A6
0510
038C
02A9
0340
04A5
057D
051C
040D
0354
0379
043B
0503
055D
04F8
0385
00F3
FDD9
FB60
FA69
FABB
FB42
FB42
FB0F
FB61
FC27
FC71
FBB3
FAAA
FA86
FB70
FC48
FC19
FB3E
FAD3
FB35
FBB3
FBAD
FB6E
FB81
FBB2
FB5F
FAC3
FB41
FDE1
01CC
04DD
05BB
0505
044D
0444
045D
03FC
0370
0379
042D
04C8
0499
03DE
0379
03EA
04C1
0525
04BB
03F2
037A
0394
0401
0473
04CA
04BE
03B0
0136
FDF2
FB69
FAA5
FB1F
FB6A
FAEE
FA8B
FB3C
FC84
FCDE
FBC1
FA7A
FAA1
FC09
FCF6
FC48
FAD4
FA40
FAFC
FBF9
FC38
FBE0
FB92
FB51
FAC7
FA6C
FB84
FE9B
026C
04DA
0514
0445
0414
04CF
0556
04C4
038F
02F3
037D
0479
04D6
0457
03AC
038E
03EF
0439
041C
03E0
03EB
0432
0469
0492
04EB
0527
0433
014A
FD4B
FA60
F9F7
FB40
FC25
FBA7
FABF
FAD0
FBCB
FC6A
FC01
FB4F
FB45
FBAF
FBA8
FB15
FAE7
FBAF
FCA6
FCA2
FBA8
FAE5
FB0D
FB71
FB30
FAC8
FBCB
FEDE
029B
04E2
0503
043C
0418
04C2
052C
049B
0391
0323
03AD
0479
04A6
0429
03C2
03FE
048B
04AD
0436
03BB
03CB
0433
045E
0436
042B
043A
036D
00E1
FD46
FAA4
FA49
FB57
FBDA
FB20
FA5C
FAE3
FC52
FD17
FC75
FB52
FAEA
FB4F
FBB4
FBBD
FBC7
FBFD
FBDC
FB19
FA72
FAE9
FC3E
FCEE
FC18
FAF7
FBC5
FF24
0333
0574
054B
043F
03F8
0486
04D0
0443
0384
037A
041B
048A
0442
03B1
0391
03F6
0449
042B
03F6
0425
0482
0461
03A6
0324
038B
042A
035B
0065
FC9D
FA46
FA44
FB64
FBEF
FB8A
FB2C
FB8C
FC2B
FC24
FB74
FAF6
FB36
FBCA
FBF4
FBA0
FB59
FB70
FB9F
FB9B
FBA0
FC0F
FCA8
FCA3
FBC8
FB2A
FC52
FF8C
0345
0562
053A
040B
0377
03DE
045D
0433
03B6
03B4
0441
04A5
046C
040C
0425
0489
0478
03D3
0371
03EF
049E
044D
030E
026A
035F
04AF
03F1
0073
FC4F
FA42
FAC4
FBED
FBF7
FB25
FADB
FB81
FC1D
FBDE
FB3A
FB27
FBAC
FBF0
FB86
FB0E
FB37
FBB6
FBBA
FB38
FB20
FC03
FD10
FCED
FB8D
FA9F
FBE6
FF4B
02EB
04F0
0522
049A
045A
046E
045F
040E
03D8
0404
045E
047A
0442
040C
0423
0469
0484
045B
0431
0431
041F
03B1
0335
0373
0494
0560
041A
0068
FC1E
F9B5
F9F1
FB4D
FBE1
FB63
FAFB
FB64
FBF7
FBC0
FAF8
FAB7
FB63
FC12
FBD7
FB11
FAE1
FB87
FC0F
FBC2
FB3B
FB7A
FC31
FC06
FAA4
F9D1
FBA5
FFEA
0403
05A6
0517
0453
047F
04F0
04AC
03FE
03F0
04AC
0530
04B9
03D2
038E
0419
0496
0465
03EB
03DD
042C
042D
03B6
0388
044F
0576
0578
0365
FFE3
FC9A
FAC3
FA60
FAB3
FB17
FB57
FB6E
FB4D
FAF2
FA9A
FAA1
FB21
FBC5
FC0A
FBBC
FB30
FAF5
FB3B
FBAC
FBDA
FBC2
FBB9
FBDC
FBC9
FB3A
FAD3
FBDF
FEEA
02BF
0542
0577
0464
03D2
0457
050F
0511
049E
0486
04DB
04E7
045A
03DA
040D
0495
0498
040F
03D6
0452
04BC
044C
039D
03FF
0563
05CD
0380
FF48
FBD6
FAD8
FB70
FBB5
FB13
FA8A
FAE7
FB9A
FBA9
FB0F
FAA3
FAD7
FB38
FB3F
FB12
FB26
FB7A
FB9A
FB61
FB2B
FB3E
FB55
FB1F
FB07
FC01
FE70
017E
03D0
04C1
04C2
04A0
04B3
04C7
04A2
0456
041D
041F
045B
04B6
04FB
04FB
04C0
0493
04A2
04C0
04A0
045C
0472
04FB
052B
03EF
0130
FE28
FC3A
FBA4
FB8A
FB35
FAD2
FADE
FB43
FB78
FB4F
FB29
FB48
FB61
FB16
FAA2
FA90
FAE0
FAFE
FAAD
FA79
FADE
FB5B
FB09
FA1D
FA35
FC97
0076
0390
0488
041F
03F1
0481
0506
04DF
0473
0478
04DC
04FA
0498
0435
0445
0499
04CB
04DC
0503
051B
04CC
0450
0478
0580
0638
04F3
017D
FD9A
FB54
FB03
FB62
FB4F
FAED
FAF0
FB60
FB91
FB2C
FAA3
FA87
FAD5
FB23
FB3F
FB3C
FB1D
FACC
FA87
FAC0
FB68
FBA3
FACB
F9A9
FA10
FCE1
00D7
03AE
0467
0401
03F4
047F
04CB
045D
03BE
03B2
0446
04ED
0543
0551
0531
04E5
0496
049B
04F2
0512
049D
041D
047B
0590
05C8
03AE
FFC5
FC47
FAEF
FB63
FC00
FBD6
FB5D
FB58
FBBB
FBF0
FBC2
FB7C
FB44
FAEA
FA6C
FA37
FA91
FB09
FB0A
FABD
FAD0
FB4D
FB4A
FA4E
F989
FADF
FE9A
02B9
04E9
04DC
0424
040E
045E
0447
03D9
03C8
0431
0465
0402
03A3
03FC
04D1
0546
0517
04D5
04E3
04DC
0471
043C
04FF
0618
05A2
028D
FE35
FB2E
FAA1
FB63
FBAF
FB32
FAE3
FB52
FBE3
FBD4
FB56
FB30
FB9F
FC12
FC05
FB99
FB30
FAE2
FAA0
FAA2
FB11
FB6D
FAEB
F9BA
F97B
FBB8
FFEF
03B9
0524
0486
03BC
03E6
0484
04A4
0441
0408
0434
0458
042A
03F1
03EF
03F4
03D1
03E0
047D
0534
0525
045E
0427
0549
0681
0583
01B7
FD3F
FACE
FAE7
FBD5
FC09
FB9C
FB70
FBA8
FBAD
FB5C
FB4A
FBC1
FC2A
FBF0
FB6A
FB55
FBA5
FB95
FAF2
FA8E
FB06
FB9F
FB26
F9E5
F9DA
FC75
00A9
03D5
048F
03D5
0375
03ED
0463
0442
0400
0435
0496
046F
03C3
0356
03A1
043B
048E
049D
04BC
04D0
0483
041C
046F
0588
05F2
0415
0046
FCCB
FB88
FC17
FCA1
FC34
FB86
FB81
FBDE
FBC5
FB2E
FAEC
FB65
FBF8
FBF6
FB8D
FB5B
FB6C
FB4B
FAFB
FB14
FB9F
FBA6
FA88
F970
FA75
FE16
0243
046B
0423
032E
031D
03B5
03E7
038F
0374
03F3
046F
045D
0416
043A
04A7
04B1
043D
03FB
044C
049A
0449
03DC
0465
05A9
05CA
0348
FF0F
FBC1
FAF5
FBCE
FC6E
FC34
FBE7
FC25
FC75
FC34
FB9E
FB62
FB8A
FB7B
FB0C
FADA
FB40
FBAB
FB69
FAD9
FAED
FBA3
FBC9
FACE
FA19
FBAC
FF8B
0355
04D9
0454
03A3
03CC
0427
03E5
0367
037E
0416
0457
0406
03D9
0448
04C2
0494
0415
042B
04D0
0503
045B
03DE
0491
0597
04C7
0150
FD14
FAC2
FAFC
FC0C
FC32
FB81
FB20
FB7C
FBEE
FBEB
FBBA
FBCC
FBE9
FBA0
FB1E
FB0D
FB89
FBDF
FB97
FB2E
FB47
FB8B
FB19
FA2E
FA80
FD54
0190
0488
04D3
03AC
0340
0424
051D
0516
0464
03ED
03DE
03D1
03C5
041F
04BF
04E3
0440
039D
03D0
047D
04A0
042B
0438
0528
057A
036B
FF6E
FC0B
FB1C
FBD9
FC32
FB70
FAB0
FAF3
FBB6
FBE7
FB76
FB2D
FB5E
FB85
FB5A
FB61
FBFF
FC97
FC41
FB2E
FA96
FB0D
FBA6
FB55
FAAE
FB7E
FE83
023B
0478
04AC
0426
042B
0497
048E
03F5
0399
03FC
04A5
04D6
0487
0431
03FF
03B2
034E
0352
03F3
0490
047C
040E
0445
0529
052C
02D2
FEB8
FB4C
FA4D
FB23
FBF8
FBE8
FB85
FB7E
FB9F
FB6B
FB11
FB24
FBA5
FBF7
FBDC
FBCD
FC1E
FC5F
FC13
FB9F
FBC3
FC42
FBF4
FA92
F9C4
FB90
FFCA
03DB
0569
04A1
0389
037A
040F
045B
0448
0459
049C
049A
0431
03D7
03E1
03F8
03AE
0342
034C
03C5
03FB
03B6
03B7
049F
058D
04A5
0141
FD16
FAAC
FAD5
FC13
FC8C
FBFD
FB71
FB89
FBCD
FB98
FB1A
FAFA
FB55
FBB5
FBD2
FBEB
FC30
FC55
FC13
FBC2
FBDD
FC18
FBA7
FAB2
FACA
FD42
0149
0467
0509
040C
036B
03DB
046B
043D
03C4
03E8
0499
04F0
0481
03E1
03B6
03EB
0410
041A
0446
046C
0427
03AD
03D7
04CD
0532
035D
FF82
FBE6
FA9C
FB6B
FC5F
FC2F
FB69
FB31
FB98
FBBF
FB44
FAD3
FB21
FBE1
FC36
FBE0
FB63
FB32
FB2F
FB23
FB3C
FB95
FBB1
FB17
FA75
FB6E
FEBC
02DA
0548
051C
03D1
0354
03EC
047F
0465
0428
0467
04CD
04AB
0421
03F1
0455
04A9
0477
0431
0463
04BF
049E
043C
0483
0564
053A
028D
FE2F
FAC9
FA14
FB32
FC10
FBD8
FB59
FB61
FBA6
FB81
FB10
FAF2
FB40
FB6C
FB2C
FAEC
FB1E
FB7B
FB79
FB33
FB3A
FB8A
FB60
FA86
FA41
FC39
0054
0451
05E8
0517
03D9
03C3
047F
04C7
0449
03E9
0454
0511
053E
04C1
044A
0449
047F
0490
048B
049B
0491
044D
0443
04EA
0584
0458
00B1
FC43
F9C6
FA25
FBA6
FC21
FB60
FAC9
FB1F
FB9C
FB4C
FA83
FA43
FAC7
FB5C
FB84
FB7D
FB8B
FB6E
FB00
FAC7
FB40
FBD8
FB7B
FA65
FA8C
FD78
0216
0584
0612
04D2
03EF
0436
04C7
04CB
048F
04C0
0540
0566
050B
04B0
04A7
04AB
0477
0450
0483
04C5
048B
0407
041E
0506
0566
0384
FF6D
FB58
F990
FA34
FB71
FBB7
FB22
FABE
FAE7
FB0F
FACA
FA72
FA88
FAE7
FB07
FAD7
FAC6
FB09
FB49
FB45
FB41
FB7B
FB86
FAE6
FA48
FB58
FEDA
0348
0607
0610
04CA
042E
049F
0516
04F0
04AB
04E9
0565
0570
0500
04AF
04BE
04CE
049C
0482
04C9
0508
04B9
043F
0482
055C
051A
024F
FDD0
FA40
F964
FA78
FB72
FB57
FAD6
FAC7
FAFD
FAD7
FA5E
FA30
FA8E
FB08
FB37
FB42
FB63
FB62
FAFD
FA92
FABF
FB57
FB69
FAAD
FA78
FC79
0088
0468
0608
0589
04B0
04AF
0527
0549
0514
0511
0550
0551
04E9
0491
04A2
04CB
049C
0452
0478
04F7
051E
04B7
0475
04E0
0530
03E2
0097
FCD2
FA8B
FA3E
FAC9
FAF5
FAA0
FA5D
FA72
FAA0
FAAE
FAB7
FADD
FAFF
FAF2
FADC
FB08
FB62
FB74
FB06
FA85
FA7D
FADA
FB02
FAE2
FB70
FDC1
0184
04E5
063A
05AA
04C7
04AE
050D
050C
049F
0474
04DB
0561
0581
054A
050E
04D8
0492
047E
04EA
0583
058D
0508
04CD
052A
04E7
028D
FE89
FB1C
F9FD
FA94
FB19
FAE4
FAC8
FB56
FBD1
FB5E
FA5F
F9E4
FA2D
FA91
FAA7
FABA
FB01
FB16
FAA6
FA26
FA41
FAD3
FB36
FB94
FD16
0037
03AB
059A
05AC
0521
050D
053E
0504
046D
0433
04B4
0578
05D8
05B9
056A
052D
050E
0503
04F0
04C8
04BB
0503
0539
045E
01E9
FEAC
FC24
FB06
FAC4
FA8F
FA58
FA85
FB01
FB3E
FB07
FAC3
FABA
FAAD
FA6E
FA4F
FA8C
FACC
FAB1
FA89
FAC8
FB1C
FAD3
FA46
FB0A
FE0E
0201
0483
04D0
045D
04A2
0553
0568
04EC
04C3
051F
0547
04E6
049A
04EE
0571
0570
050D
04F4
0523
0507
04BB
050B
05BF
0507
01B3
FD37
FA60
FA33
FB1A
FB45
FAC0
FAA9
FB25
FB3C
FA8A
F9F3
FA3F
FAFD
FB4C
FB13
FAC2
FA7C
FA39
FA4A
FAD9
FB3A
FAB0
F9F3
FAEF
FE7D
02DD
056C
0587
04E4
0504
0575
052A
0463
043D
04FD
05CA
05FC
05B4
0543
04BD
0456
047E
052D
0593
0529
04AC
0519
05B6
046D
0096
FC5B
FA50
FA8C
FB14
FAB5
FA24
FA5C
FB16
FB5C
FAFB
FA80
FA27
F9BE
F97A
F9F4
FAFA
FB78
FB03
FA90
FAE0
FB35
FAAA
FA38
FBE9
FFFF
0412
05BD
053E
04AD
0511
0584
0533
04B3
04CC
0520
0507
04DF
0567
0648
066E
05B2
050D
050D
0519
04B6
048E
0536
0578
035B
FF03
FB2C
F9FD
FAA0
FAE7
FA5B
FA33
FAE8
FB6B
FAF4
FA44
FA6C
FB1D
FB25
FA4F
F99D
F9B5
FA14
FA44
FA9C
FB34
FB43
FA88
FA8D
FD0C
015D
04C6
059B
04F5
04D7
0587
05B6
04EB
044B
04C5
05A5
05C2
052D
04CB
04ED
053D
0594
05F4
05FA
0543
0465
047C
055A
050E
021C
FDBF
FAD9
FA95
FB4B
FB19
FA42
FA22
FAD7
FB3F
FAD7
FA4C
FA3B
FA67
FA7A
FAA6
FB0F
FB2D
FA98
FA06
FA72
FB5E
FB51
FA69
FAEF
FE58
02D8
054D
0502
041C
046B
0554
0561
04A6
0470
0515
058B
0542
0504
0574
05DE
0579
04CC
04C1
0515
04E6
0466
0498
0537
0452
00CE
FC73
FA3A
FAC7
FBE5
FBAE
FAC1
FAA5
FB49
FB6D
FACB
FA61
FABB
FB2A
FAF2
FA5F
FA29
FA5F
FAA0
FAE1
FB48
FB6E
FADD
FA70
FC02
FFF4
0409
05B7
0501
0409
0432
04D4
04DB
046D
046A
04EB
0533
04ED
049A
04A4
04CF
04E8
0527
0579
0545
0485
044D
0528
05A2
039C
FF32
FB21
F9D8
FAD7
FBBD
FB6B
FADB
FB0B
FB7A
FB49
FAC4
FAC3
FB32
FB57
FB20
FB20
FB6D
FB6F
FAFA
FAB7
FAFE
FB0E
FA5E
FA2B
FC69
00EE
04EE
0611
050F
044A
04AB
0521
04CD
0448
046D
04F3
04FC
047D
0439
0479
04B4
0498
0487
04B9
04C6
0491
04C6
058E
0579
02E7
FE71
FAC5
F9D0
FAC9
FB88
FB34
FAB7
FAE2
FB3E
FB15
FAA9
FAA6
FB0B
FB59
FB77
FB9C
FBAC
FB62
FAFE
FB04
FB49
FB09
FA56
FAB7
FD89
01DF
051A
05C1
04F0
0484
04D3
04F4
049D
047C
04F3
0579
0579
051E
04DA
04A7
044A
03FF
0438
04BC
04DB
049E
04CC
0553
04A8
019F
FD5D
FA66
F9DD
FA9A
FB00
FAE0
FB00
FB80
FBA2
FB15
FA77
FA5A
FA83
FA98
FACD
FB54
FBB6
FB79
FAFE
FAF7
FB3B
FB19
FACE
FBCB
FEE6
02D3
0551
05AD
0541
0556
0597
0524
0442
03F8
0486
052D
055F
0551
054E
052B
04C4
047A
04AC
0503
04F5
04B7
04DF
04F4
037B
0001
FC3F
FA5B
FA72
FAE1
FA92
FA1C
FA63
FB20
FB63
FB00
FAAC
FAC3
FAE0
FABB
FAB8
FB0E
FB3F
FAEC
FA92
FABB
FB06
FADA
FAD8
FC80
0022
03ED
05C6
0595
0507
053B
05A3
0568
04DC
04CB
052F
0560
052D
04F8
04E5
04B3
046B
047A
04F4
0548
0517
04DE
050F
04D2
02BF
FEF7
FB91
FA4A
FA97
FAC7
FA54
FA17
FA8A
FAFE
FAC6
FA45
FA49
FACC
FB1B
FB03
FB05
FB55
FB77
FB31
FAFE
FB1E
FB03
FA89
FAF0
FD91
01BD
04FF
05CA
0510
04C2
0556
05BA
0552
04E7
053C
05D4
05D0
0540
04CD
049D
0466
043D
047A
04E3
04D7
0467
0473
0520
04E2
021E
FD9E
FA34
F99B
FAA3
FB1F
FA9A
FA3C
FAA4
FB1C
FAEC
FA63
FA2E
FA65
FAAF
FAF8
FB60
FBAF
FB88
FB29
FB2F
FB79
FB38
FA8F
FB29
FE3B
028F
058B
060A
0542
04DD
0517
0530
04EF
04DC
0523
0541
04FF
04DF
0526
0545
04CD
0446
044D
048B
0464
042A
04A9
0568
0495
0140
FCFF
FA6C
FA3E
FADB
FACD
FA6C
FAA3
FB37
FB49
FADC
FAB2
FAFD
FB2C
FAFE
FAE0
FB15
FB36
FAFC
FAF2
FB88
FBFD
FB55
FA62
FB6E
FF3D
0387
0580
050A
0453
04B9
0578
0569
04D2
04B3
051D
053B
04CE
0484
04BC
04EA
04AD
0482
04CA
04F4
0481
041E
0494
050B
03A0
FFF5
FC20
FA73
FAE7
FB96
FB55
FACA
FACF
FB13
FAE9
FA88
FA8C
FADC
FAFC
FB00
FB50
FBB5
FB90
FAFC
FADB
FB6E
FBBD
FB1D
FAD0
FCCD
00E8
047B
0573
049B
0412
0481
04F0
04CD
04AC
0508
056F
0556
0504
04FD
0508
0497
03EF
03E9
047D
04B0
0448
0453
0528
0518
0268
FE05
FAD9
FA64
FB49
FB81
FAF4
FAE3
FB8B
FBC0
FAF2
FA24
FA4C
FAE1
FAF5
FAC5
FB1C
FBC9
FBEE
FB7D
FB49
FB81
FB52
FA98
FAEB
FDD6
0255
0578
05BC
04A4
045A
04FD
0539
04AA
0444
04A5
0544
0578
0553
0531
0501
049A
0445
0459
047A
0426
03DB
048E
05B0
0507
016A
FCC1
FA1E
FA44
FB4A
FB66
FADB
FAD6
FB67
FB9B
FB17
FA8D
FA80
FA9E
FA9F
FADB
FB68
FB9C
FB23
FACC
FB49
FBDA
FB59
FA6A
FB4D
FEFA
037A
05EC
05C3
04F0
04FC
0560
050E
044E
0418
0477
04BB
04C8
0515
058C
0579
04C4
044F
04AB
052F
0503
0497
04E4
055C
03F8
0007
FBAC
F99E
FA15
FB08
FB01
FA75
FA66
FADB
FB37
FB51
FB7D
FBB0
FB86
FB0D
FAD3
FAFB
FB00
FAB9
FAB7
FB21
FB24
FA5D
FA2B
FC5F
00B4
04AC
063E
05DA
054E
0558
054B
04C6
0478
04D4
052D
04CE
042E
0423
048A
04A7
047B
04B2
0553
0589
050D
04D0
0570
05A2
036B
FEF6
FAF4
F99B
FA43
FACD
FA71
FA1E
FA81
FB0A
FB12
FADA
FAF8
FB52
FB61
FB29
FB2B
FB72
FB72
FB07
FACC
FAFF
FAFC
FA7A
FAA3
FCE7
00E4
046F
05DC
0590
0516
0534
057E
0578
054E
0550
0557
052A
04EB
04C8
04A6
0477
047E
04CF
04F2
0494
043F
04A7
0553
04B8
020C
FE7F
FC04
FB36
FB12
FAB6
FA68
FA8E
FABA
FA65
F9F6
FA25
FAC3
FAF8
FAA5
FA98
FB36
FBB5
FB58
FABA
FAF3
FBBF
FBBE
FADA
FB12
FDF7
0240
0509
0534
0457
044F
0511
0569
050F
04E5
0560
05DD
05BD
055B
0549
0550
04F2
0475
0488
0510
052D
04A3
045B
050A
05C9
04CC
018B
FDA0
FB2C
FAC5
FB54
FB92
FB36
FAB6
FA88
FAB9
FAFD
FAFF
FAB6
FA69
FA64
FAA5
FAEA
FAF3
FABA
FA6C
FA49
FA78
FAE5
FB37
FB38
FB66
FCCF
FFDF
0360
0558
0530
0457
0474
056E
05E5
053F
0465
045C
04E9
0526
04F8
0506
0576
05A2
054C
052A
05A5
05EA
051D
03F5
03FA
0512
0506
0226
FDBB
FAC0
FA71
FB2C
FAFD
FA09
F9C9
FAA3
FB80
FB8F
FB42
FB44
FB5B
FAF7
FA48
FA0C
FA59
FA7F
FA35
FA38
FB0E
FBE2
FB75
FA27
FA09
FC9D
00EC
0471
05A8
054B
04FE
0566
05D5
059C
04F4
0488
0487
0497
0482
047B
04BE
0519
0532
050F
050D
0544
0554
050F
04FA
0584
05D9
044F
0072
FC1D
F9E0
FA4D
FB85
FB94
FA93
F9FB
FA63
FAE6
FACA
FA91
FAFA
FBB0
FBD0
FB5E
FB34
FB90
FB9B
FACD
F9F6
FA1D
FACD
FAB9
FA0C
FAD5
FE5F
02FA
0590
0525
03BA
0394
04B2
0590
0586
055D
05AB
05D6
052F
0437
03EC
0455
0495
0459
0451
04F0
0595
0575
04F1
0511
05BC
0548
0276
FE57
FB6E
FB05
FBEF
FC39
FB5F
FA6C
FA3E
FA7F
FA7A
FA47
FA98
FB7F
FC1F
FBC8
FAF2
FA99
FAEF
FB3F
FB14
FAD4
FAF6
FB22
FAD0
FA91
FBDD
FF30
02EE
04E6
04C2
0434
04A9
05A5
05DD
0531
04B0
04E0
050C
048D
03F9
0445
0535
059A
050A
0471
048E
04CF
0464
03CE
043F
0578
056E
02AF
FE6F
FB5B
FAA3
FB04
FADF
FA38
FA1E
FAD0
FB76
FB7E
FB4F
FB66
FB7E
FB29
FAB3
FACB
FB63
FBAA
FB4E
FB19
FBBD
FC82
FC04
FA5D
F9A8
FBD0
003B
0434
05BA
054A
04C8
0522
05A3
0563
049D
0434
0467
04A5
048D
0471
04A9
04E8
04B2
042F
040B
0461
0487
042C
0416
0506
0604
04EA
00FE
FC53
F9D5
FA2E
FB6A
FB95
FACF
FA76
FAF6
FB76
FB5F
FB31
FB76
FBC4
FB7E
FAF9
FB0F
FBBF
FC13
FB96
FB0B
FB36
FB8E
FB0E
FA24
FAC0
FDF4
024A
052C
059A
04DC
048E
04F1
0547
052B
04E3
04B0
0476
0435
043A
0495
04C2
0455
03C3
03DE
04A6
0520
04B1
040C
0454
055C
0569
0305
FEDF
FB55
FA1F
FAC5
FB7D
FB43
FAA3
FA96
FB2E
FBA7
FB87
FB28
FB1E
FB6D
FBB4
FBCD
FBDE
FBDB
FB8C
FB21
FB32
FBCE
FC11
FB4D
FA72
FB7E
FF1F
0375
05D1
058E
0472
0446
04E8
0526
04B7
046F
04C0
050A
04AB
0404
03E5
044E
0486
044C
0428
046B
0497
0446
040D
04AB
057E
04C1
01A8
FDA1
FAFE
FAA4
FB7A
FBFD
FBC4
FB43
FACD
FA65
FA3E
FAB2
FB9B
FC3D
FC18
FB85
FB38
FB62
FB93
FB7D
FB5E
FB7D
FB8A
FB0E
FA6A
FAEA
FD6F
0130
0427
04F4
041A
0356
03C2
04E7
05A1
0586
051E
04F3
04EC
04B6
045B
042D
043C
0453
0464
049F
04FC
0519
04D1
04A1
04EA
04E8
033F
FFD8
FC8E
FB58
FC0E
FCB2
FBEC
FA8C
FA2C
FB03
FBC6
FB8F
FAE5
FAB8
FB06
FB32
FB23
FB47
FBA2
FB9F
FB0A
FA92
FAD4
FB5B
FB4B
FAEC
FBB4
FE67
01D1
03FF
046F
0455
04C7
056E
0557
0485
03F7
0446
04EA
0518
04CD
04A5
04DA
0507
04E6
04C0
04E6
051B
04F1
048B
0485
04F3
04D6
030D
FFBA
FC6E
FAAE
FA97
FB16
FB45
FB2A
FB33
FB67
FB70
FB38
FB0C
FB1E
FB2D
FAF0
FA96
FA87
FACB
FB06
FB1A
FB4D
FB9C
FB6E
FA79
F9C8
FB20
FEED
034D
05BB
0599
0482
042F
04AC
0501
04D5
04BC
0509
0540
04F2
0487
04A8
0531
0569
0525
0501
053B
052E
0472
03E2
049B
05FE
05C2
028C
FDE4
FAC6
FA72
FB6B
FBAC
FAFF
FA9B
FB0D
FB89
FB43
FA96
FA65
FACE
FB2A
FB14
FADD
FAE0
FAEF
FAC3
FA9B
FAD9
FB36
FB0A
FA7C
FAD9
FD36
00EB
03F7
0502
04A2
045F
04DD
0569
0543
04B3
048A
04FB
0569
0557
0504
04EF
051B
0526
04F2
04C4
04C3
04BA
049F
04E1
05A3
05E3
042B
0064
FC78
FA88
FAC4
FB7E
FB5B
FAB6
FAA0
FB27
FB62
FAF8
FAA2
FAF3
FB5B
FB07
FA3D
FA0C
FAC2
FB7C
FB87
FB58
FB98
FBC7
FAE9
F989
F9E2
FD52
0240
0585
05C4
0495
0435
04FB
05A5
0572
04F9
04EB
0501
04AC
0433
0457
0517
0596
054D
04BB
0486
048C
0453
0424
04CE
0622
065F
03EE
FF74
FB8A
FA2B
FADC
FBA7
FB63
FA99
FA49
FA93
FADF
FADF
FAE2
FB24
FB6D
FB77
FB6D
FB96
FBC6
FB9C
FB2E
FB03
FB2D
FAFF
FA21
F9A1
FB33
FF18
0351
0578
0535
044F
0469
054C
05C0
055F
04E7
04EE
0514
04D2
0461
044F
0484
045D
03CB
0390
0422
04E1
0506
04E3
0562
063C
05A3
025E
FDB6
FA7F
FA22
FB4E
FBDB
FB38
FA74
FA5D
FA8E
FA79
FA6F
FB05
FBEB
FC2F
FBA6
FB3E
FBAC
FC5C
FC4D
FB88
FAFF
FB0D
FAF9
FA5F
FA5B
FC80
009B
0476
0606
0577
0486
0460
04CA
0523
0567
05CC
0608
059F
04C8
044F
0481
04B4
0443
0389
0360
03EA
0477
04A2
04E7
059C
05DA
0424
004D
FC26
F9E4
F9F9
FAF3
FB4A
FADC
FA7D
FAA1
FAE6
FAD4
FA80
FA49
FA4F
FA78
FAD3
FB84
FC4F
FC9B
FC30
FBA1
FB8C
FBAA
FB39
FA7A
FB03
FDFF
0261
0593
0628
0546
0502
05CF
0653
0594
0456
03FA
04AC
057C
05C2
05B4
0593
0520
044A
03BD
0411
04BD
04B1
03F0
03B5
047A
04CA
02DC
FF07
FBA6
FA73
FAC2
FACA
FA01
F964
F9C2
FAAA
FB3F
FB67
FB7D
FB7A
FB18
FAA7
FAD5
FB97
FBF2
FB4A
FA64
FA7A
FB78
FC08
FB83
FB2C
FCC5
0041
0395
0509
04FA
04F5
05A2
0639
05F2
052E
04D7
050D
0517
0493
040C
041D
0485
0498
045B
0476
0511
0567
04EB
0451
04A3
0577
04DD
01B1
FD65
FAAA
FA7C
FB40
FB14
FA16
F9C4
FAA5
FB95
FB89
FB04
FB2D
FC06
FC65
FBB0
FABA
FA87
FAF1
FB14
FAC4
FAAA
FB08
FB3D
FAF1
FB1D
FD15
00A2
03D5
0516
04CA
0488
050E
05A1
056B
04A2
0417
040A
040C
03DA
03BE
0401
0475
04D2
0531
05BD
0626
05F1
0554
0523
0590
056D
0357
FF97
FC34
FAE5
FB56
FBDA
FB7F
FADB
FADA
FB6E
FBD9
FBD0
FBBB
FBE4
FC02
FBC8
FB78
FB7C
FBAC
FB75
FAC4
FA35
FA3B
FA6F
FA35
F9EF
FAE7
FDD2
01AD
0487
0568
0515
04E7
0533
053D
047D
037A
0330
03CC
0482
0494
043B
042E
0492
04CD
047A
0412
044F
0525
05CA
05CF
05AC
05EA
0605
04C3
01B6
FE0D
FB7E
FAA9
FAD2
FB0A
FB20
FB66
FBE8
FC44
FC36
FBED
FBC0
FBB7
FB99
FB51
FB12
FB0E
FB32
FB3E
FB0E
FAC2
FA9C
FAA1
FA89
FA2E
FA1D
FB55
FE3E
01EB
04A7
0579
04ED
0450
044D
0483
046A
041B
0406
0438
044E
041C
03F6
0434
04B1
04F9
04E5
04C7
04EE
0530
0531
04F1
04E5
0544
0570
044F
0170
FDCC
FB25
FA7C
FB38
FBEC
FBE4
FB9B
FBB4
FC01
FBDE
FB45
FAF1
FB57
FBF4
FBFA
FB71
FB25
FB6F
FBB4
FB59
FAC5
FAD5
FB7E
FBB8
FAFA
FA55
FB86
FEEC
02DD
0533
0550
045B
03C2
03DD
0417
03FE
03D0
0404
0498
0510
050D
04AF
0451
040D
03C6
038B
03AC
0441
04DA
04F3
04B0
04C7
0571
05B5
0434
00BE
FCE2
FA99
FA7A
FB73
FC1F
FC1A
FBEF
FC0C
FC2F
FBE2
FB37
FAC4
FAEE
FB75
FBD7
FBF0
FC02
FC2F
FC34
FBD1
FB43
FB09
FB21
FAE9
FA1C
F9B5
FB42
FF0E
0356
05C0
059C
045C
03C9
0430
0498
045C
03F7
0422
04B4
04E8
0482
041F
0448
04AE
04A2
0421
03DA
0433
04B2
04B5
0477
04D6
05F1
0675
04CA
00F0
FCCA
FA68
FA34
FAED
FB47
FB21
FB20
FB8B
FBF0
FBDB
FB7F
FB57
FB79
FB7E
FB34
FAF3
FB23
FB96
FBB0
FB3D
FACD
FAF7
FB70
FB4B
FA51
F9C2
FB4A
FF14
034A
05B6
05D8
0513
04E3
054F
055B
049D
03D4
03D5
0477
04EB
04DC
04C0
04FE
054B
051F
0495
0458
04B5
052B
0524
04D0
04EB
0586
058B
03BB
0026
FC66
FA3A
FA00
FA9B
FAD8
FA9B
FA9B
FB2A
FBBC
FBAE
FB24
FAC9
FADE
FAF3
FAAF
FA73
FAC9
FB71
FB94
FAFE
FA8C
FAFA
FBA9
FB57
FA10
F9B6
FC1D
00C6
0518
06E4
0655
0540
04F2
0534
0534
04D7
04B3
0517
0590
0580
04F7
04A7
04FA
0584
058D
0503
048F
04AD
0507
04FA
0499
04AE
056A
0592
038A
FF54
FB03
F8D5
F91A
FA46
FAE5
FAE4
FAEF
FB26
FB05
FA65
F9EC
FA34
FAED
FB3D
FADC
FA67
FA78
FADD
FAF6
FAAD
FA9D
FB30
FBE1
FBCC
FB03
FAE6
FCD8
00A0
0468
066F
068F
05F9
05A6
0586
052C
04CC
04FE
05B8
061F
05A5
04E0
04D2
058B
060D
05A9
04EB
04D3
0565
059B
04DC
03F0
0406
04F8
0514
02E5
FEEB
FB48
F9B9
FA19
FADA
FACC
FA24
F9D2
FA38
FACC
FAEB
FAA2
FA79
FA9A
FAA6
FA59
FA10
FA47
FACC
FAEF
FA88
FA53
FAF2
FBD7
FBE2
FB0C
FAEF
FD25
0144
0506
0683
05F1
0503
04E5
055A
059A
057B
056A
0597
05B1
056F
0516
0520
0592
05EF
05DA
0584
0554
054F
0519
0496
0445
04A9
055D
050B
02AA
FEC0
FB2D
F984
F9B9
FA83
FADE
FADF
FB07
FB47
FB19
FA6D
F9F2
FA33
FAC6
FAC9
FA21
F9B0
FA2B
FB17
FB63
FAD1
FA4E
FAA5
FB5C
FB5D
FAA3
FAA9
FCDA
00C9
0465
05FD
05C8
0542
0560
05B6
056C
048B
03FD
0465
0562
0617
0630
060C
05FF
05D9
055B
04D3
04DA
056F
05CD
0569
04C8
04DE
0593
0570
0324
FF3D
FBD9
FA8C
FAE9
FB4C
FAD0
FA0F
FA07
FAC7
FB7B
FB7F
FAFF
FA7F
FA2F
F9F2
F9D1
FA04
FA82
FAD8
FAAF
FA54
FA63
FAF2
FB46
FABF
F9EC
FA59
FCF9
00EB
0413
0514
0488
041B
04B3
05B5
0617
05BE
0566
0581
05A2
0548
04BD
04C6
0588
063C
062E
05A1
0565
05AB
05CD
055B
04EA
0548
0618
05B9
0309
FEE9
FB9F
FAA2
FB4E
FBDA
FB57
FA5F
F9F2
FA2B
FA59
FA19
F9E3
FA49
FB20
FBA1
FB5B
FAAA
FA30
FA17
FA19
FA0F
FA28
FA72
FA89
FA1B
F9B3
FA91
FD65
014C
045A
0560
04EF
048E
0506
05C7
05E3
054F
04E1
052C
05CE
0604
059C
0518
04EA
04F9
0504
0522
0591
061D
0634
05B6
055B
05CC
0673
05AE
0288
FE15
FAA8
F9A6
FA54
FAEE
FAA2
FA1E
FA52
FB1F
FB93
FB32
FA86
FA4F
FA8C
FAA6
FA65
FA3C
FA92
FB10
FB14
FAA1
FA6B
FACA
FB10
FA76
F982
FA02
FD27
01EB
05C7
070B
064F
0571
0574
05C8
0582
04B6
044B
04B3
0561
058A
0534
050A
056C
05ED
05F2
057A
04FC
04AD
045B
0407
043C
0547
064A
0599
0266
FDE9
FA73
F954
F9DA
FA67
FA43
F9FE
FA4C
FAFC
FB4A
FAF0
FA7A
FA86
FAF9
FB33
FAE8
FA73
FA58
FAA0
FAF9
FB45
FBB1
FC30
FC39
FB71
FA91
FB28
FE08
0218
051F
05E7
054A
0501
05A8
0656
061C
0549
04EA
0558
05D1
05A0
0506
04C9
0507
0525
04C8
046A
04A5
0535
0532
0457
038C
03C6
0494
0441
01B3
FDDE
FAFC
FA5A
FB2D
FBB0
FB1A
FA2C
F9EB
FA54
FA97
FA51
F9FF
FA2D
FAB1
FB01
FB0A
FB38
FBA8
FBD3
FB51
FA98
FA8F
FB55
FBF4
FB9D
FAF2
FB9D
FE7E
027F
0575
061C
051C
0428
0447
0514
0599
0584
0557
0588
05DA
05BF
052B
04A9
049D
04C4
04B0
047D
049F
050F
052A
04B6
0472
051B
05F7
0524
01AF
FD0E
F9E9
F979
FA8D
FB3A
FAFD
FABD
FB20
FB9A
FB5A
FA8B
FA23
FA9E
FB61
FB98
FB3F
FB03
FB39
FB6C
FB28
FAB8
FACA
FB5E
FB8F
FAC4
F9DE
FAAD
FE00
0280
05C4
0692
05CB
0520
053C
057A
0528
0485
044E
04A9
04FD
04D9
0490
04B0
0526
054A
04D8
0462
0491
0528
0549
04B2
0444
04DD
05E1
056F
0263
FDE3
FA6C
F973
FA31
FAE3
FABE
FA52
FA5A
FAC1
FB07
FB1D
FB60
FBD7
FC06
FB9A
FAF4
FAA8
FAB6
FAA4
FA5A
FA65
FB34
FC3E
FC65
FB53
FA40
FAFD
FE26
0258
055A
0616
055B
04C7
0514
05AF
05CD
0577
054E
0570
054A
0486
03BF
03CA
049C
0555
0573
0566
05B6
05F6
0552
03FB
034A
040C
0517
0451
0111
FD08
FA85
FA3D
FB00
FB66
FB31
FAFA
FB0D
FB01
FA80
F9E3
F9DE
FAA3
FB94
FBE5
FB6D
FAC1
FA7C
FAA0
FABC
FAA1
FAA2
FB01
FB69
FB60
FB30
FC03
FEA6
025B
0554
0660
05F7
055E
0533
0520
04D3
049E
04EF
0587
05B7
0553
04EB
04FB
0539
0517
04A9
0492
0514
059C
0597
054C
0579
0615
05F7
040C
00A5
FD49
FB36
FA64
F9FF
F98A
F949
F9A4
FA76
FB22
FB3C
FAF5
FAD0
FB07
FB4D
FB35
FAC8
FA89
FACD
FB36
FB2A
FAB1
FA79
FAC4
FAD9
FA09
F922
FA16
FDC8
0299
05D5
0677
05E5
05E2
0686
06C2
062E
0586
0565
056A
04F3
0430
03E3
0446
04CB
04FF
050F
053D
055B
0534
0513
0566
060B
067C
0684
0642
057F
0390
0048
FCAC
FA35
F961
F974
F9A3
F9D7
FA2D
FA62
FA4A
FA59
FB0E
FC0A
FC64
FBE5
FB52
FB3C
FB2E
FA7E
F990
F971
FA43
FAE1
FA85
F9DC
F9F4
FAA5
FB08
FB46
FCCB
0055
047C
06F0
06ED
05D3
0548
0584
05AF
0545
0489
03ED
03A7
03CF
0453
04DA
0512
0529
0599
0659
06AA
060E
0520
04E6
0567
059F
0503
0456
0457
0441
027E
FEE1
FB46
F9A6
FA04
FAD0
FAFA
FADA
FB1E
FB9E
FBC8
FB9B
FB8E
FBB2
FB95
FB10
FA94
FA83
FA9D
FA7C
FA45
FA67
FACD
FAE5
FA97
FA91
FB44
FC16
FC3E
FC2B
FD47
0030
03AB
05D0
05F8
0519
0470
045F
049D
04E4
050F
04F5
04A2
047D
04CB
0531
0525
04C9
04D1
0571
05E7
057B
049C
044C
04AA
04D1
0465
043E
04EA
053C
035D
FF50
FB70
F9F9
FAB4
FB9F
FB75
FAC7
FAA1
FB0F
FB65
FB5A
FB28
FAF4
FABB
FAB7
FB25
FBA7
FB79
FA8A
F9DB
FA58
FB93
FC46
FBF0
FB45
FAED
FAAC
FA54
FACE
FD3E
0134
049D
05CD
0521
0446
0448
04D9
0547
056A
056B
0550
0519
04FB
050A
04F3
047D
041A
0465
052C
0587
0515
048F
04BE
0545
052E
047E
0451
0506
052A
0309
FF03
FB72
FA22
FAA5
FB50
FB48
FAF6
FAD5
FABE
FA7F
FA69
FAC7
FB45
FB64
FB4E
FB89
FC01
FBFF
FB3B
FA6A
FA5B
FAE6
FB40
FB2D
FB24
FB47
FB0C
FA6B
FAB0
FD37
0171
0508
0631
0569
0488
0493
050C
0528
04E8
04B7
04B3
04BD
04DC
050C
04F6
0461
03C6
03DE
049C
051A
04DB
0488
04F2
05BF
05ED
0574
055E
05D9
0540
0219
FD75
FA3C
F9FA
FB52
FBFC
FB77
FB00
FB56
FBD0
FBB1
FB57
FB62
FB8E
FB3C
FAAD
FAC1
FB91
FC33
FC04
FB79
FB3D
FB1C
FA88
F9D4
F9E5
FAA5
FAEF
FA7D
FAEA
FDC2
021D
0543
05B8
04A8
0410
0468
04C2
049E
047D
04AE
04AA
041E
03B4
0425
0503
0551
04F4
04B0
04DA
04E9
048C
0463
04FF
05C3
05AC
04FA
04EC
0598
0529
022D
FDE2
FB09
FAC9
FBA9
FBCF
FB2F
FAE5
FB45
FB8D
FB5D
FB5A
FBFA
FC9A
FC6A
FBA0
FB0E
FAE5
FAC1
FAA7
FB13
FBE9
FC2D
FB5B
FA5C
FA5F
FB11
FB1E
FA85
FB30
FE72
02CF
0568
054D
0444
0438
0503
0544
04A7
041F
043B
0455
03D6
034B
0384
044B
04BF
04A5
0487
04AF
04BF
0490
0497
0516
056D
04FF
0464
04A5
054D
045B
00D3
FC7E
FA1C
FA55
FB62
FB9F
FB46
FB5E
FBE5
FC08
FBAA
FB94
FC09
FC42
FBC0
FB3C
FB87
FC35
FC40
FBA9
FB6A
FBCE
FBF7
FB55
FABA
FB1F
FBEF
FBD2
FB19
FBF9
FF9B
0411
0654
05BB
045F
0423
04AC
04A5
03F0
0396
03FF
0469
043D
03F7
0436
04A7
049E
0428
03D3
03B7
0383
035E
03D2
04BE
0522
0480
03D4
0433
04D2
0396
FFEA
FBF4
FA39
FAC0
FB8C
FB65
FAFD
FB48
FBF0
FC0A
FBA7
FBA3
FC22
FC48
FBAF
FB22
FB66
FC12
FC4D
FC2C
FC5C
FCC0
FC7A
FB6C
FABF
FB43
FC10
FBD2
FB1C
FC25
FFC8
03F7
05FA
058D
04B2
04DF
057D
0565
04A7
042A
042A
0413
03B7
03A9
0426
047D
0423
0398
03A6
0420
0448
0415
0430
04B5
04DA
0447
03F2
04AD
0556
03BD
FF90
FB53
F99B
FA3F
FB13
FAE0
FA6E
FAC0
FB82
FBD7
FBCC
FC11
FC98
FC8E
FBD2
FB5B
FBC9
FC5C
FC25
FB75
FB4A
FBB0
FBBB
FB27
FADF
FB72
FBF8
FB78
FAE8
FC72
007B
049E
0650
05BD
0501
0534
057A
04E2
03EB
039D
03EF
040B
03BC
03B8
044B
04C5
0496
0435
044E
04A6
049E
0466
04AD
0552
0556
0472
03D2
0462
04FF
037B
FF8C
FB8E
F9D9
FA3C
FADC
FADB
FAEF
FBAD
FC70
FC66
FBD8
FB9C
FBC7
FBB8
FB57
FB55
FBEC
FC50
FBDC
FB1F
FAF7
FB3D
FB23
FAB4
FAD4
FBA8
FC06
FB3E
FAB7
FC96
00D0
04BE
0615
0557
049B
04BF
04E3
0457
03BB
03D9
0469
049E
047A
049F
0504
04D6
03DE
031F
0381
048D
0528
051E
0514
0537
0501
0465
043F
04EF
051D
030E
FF0C
FB8E
FA79
FB2B
FBBD
FB7E
FB40
FB93
FBED
FBB5
FB3E
FB2D
FB68
FB59
FB08
FB24
FBDE
FC87
FC95
FC56
FC2C
FBBE
FAB9
F9DC
FA38
FB7B
FC07
FB46
FAF6
FD37
018B
050B
05B9
04A4
041D
04BC
053E
04CD
0423
042A
049D
04A7
044A
0449
04D0
0519
049E
03DA
0385
039A
03BD
040C
04C6
057A
0568
04B9
047D
0500
04D8
026D
FE45
FAD5
F9D6
FA94
FB40
FB31
FB0C
FB46
FB7F
FB6C
FB6C
FBD9
FC46
FC15
FB7D
FB4A
FBB1
FC08
FBDC
FB94
FBA5
FBC1
FB7C
FB34
FB84
FC07
FBAC
FA8F
FA9D
FD86
024B
05F5
06BE
05BB
04FF
0516
0511
0480
041C
0473
04E9
049C
03BD
034D
03B8
0465
04AA
0496
0482
0478
046F
04A2
0512
0526
0470
03A0
03E1
04FD
04ED
020C
FD64
F9E5
F94A
FA76
FB42
FB07
FABB
FB0E
FB87
FB83
FB39
FB43
FB9D
FBC1
FB80
FB40
FB49
FB69
FB73
FB8C
FBB6
FB93
FB02
FAA1
FB05
FBBD
FBD1
FB6D
FC29
FF22
032C
05C5
05D6
04BE
0460
04F6
0568
0526
04CC
04F0
0542
0531
04DA
04CC
0517
0538
04ED
0493
047A
0478
0467
048A
050D
0578
0548
04D5
04E0
051D
0403
00A9
FC6F
F9E6
FA11
FB6D
FBEE
FB44
FA91
FA85
FAA9
FA74
FA2D
FA59
FAD0
FAFA
FABB
FA97
FADE
FB3D
FB53
FB36
FB20
FB07
FAE0
FAED
FB4B
FB6C
FAC2
FA01
FAFA
FE92
0340
0641
066B
0529
048B
050C
05AD
05B7
0582
0592
05C3
05AA
0553
0527
0539
0537
04FF
04DA
0507
0557
058B
059E
058A
0523
048B
0478
0555
062B
0523
0193
FD20
FA46
F9D4
FA67
FA6F
F9EB
F9CB
FA53
FACD
FABA
FA73
FA77
FAAB
FAAF
FA96
FABD
FB1B
FB37
FAEE
FAB5
FADE
FB09
FAC3
FA4A
FA33
FA7B
FA9E
FAB7
FBD7
FEBA
027D
0535
05EB
0572
052B
0579
05D1
05D6
05BB
05AB
057C
051D
04EA
0535
05B0
05BE
0548
04D6
04D1
0501
0509
04F5
0517
057F
05FC
066E
06A5
05F8
03A1
FFCF
FC0A
FA11
FA30
FB1E
FB80
FB28
FABF
FAAC
FAC5
FAE0
FB12
FB5B
FB6E
FB18
FA96
FA51
FA5F
FA8C
FABD
FAF7
FB13
FAD5
FA69
FA5C
FAC1
FAE2
FA42
F9CC
FB3F
FF1B
039F
065F
06A7
05D0
055B
055D
0519
0471
040E
0442
0493
0482
0446
0463
04DC
053C
0551
056B
05BA
05E7
059C
0521
0502
0545
0566
052E
0513
0583
0603
0569
0304
FF66
FBFB
F9F8
F9A4
FA72
FB7A
FC0B
FC0C
FBDF
FBDE
FBF9
FBEC
FBAB
FB6B
FB49
FB1B
FAB7
FA40
F9FE
F9FF
FA2B
FA8C
FB39
FBE4
FBEA
FB1E
FA3A
FA22
FAD2
FB86
FC07
FD38
FFE2
0343
0574
0572
0435
0374
03B6
042F
042B
03FA
043D
04E0
0541
052F
0528
058E
060C
060B
057E
04D5
0464
0429
0423
0476
050A
055D
050E
0474
044C
04BC
04DB
038F
00C3
FDA1
FB8E
FB0D
FB90
FC20
FC28
FBB7
FB37
FAF4
FAE0
FAC4
FA85
FA44
FA35
FA68
FABE
FB11
FB4D
FB73
FB94
FBC4
FBF9
FBF8
FB95
FB13
FAF9
FB5F
FBA5
FB34
FA9B
FB61
FE61
026E
0532
057E
0460
03C2
0449
0513
053B
04FA
050E
0586
05BA
0558
04DE
04D7
0511
04F9
0485
043C
0465
0499
0460
03F0
03E2
0459
04D1
04E8
04EC
0542
056E
043F
012B
FD4A
FA89
F9F3
FAD2
FB9F
FB94
FB1F
FAFA
FB2E
FB38
FADC
FA86
FAA8
FB20
FB61
FB33
FAF5
FB11
FB75
FBBF
FBD0
FBDA
FBF1
FBDD
FB84
FB38
FB40
FB53
FAFA
FA9A
FB8E
FEBA
0325
0673
0715
05B6
0447
03F7
0466
04B0
04A4
04AC
04F2
0518
04E0
049C
04BC
0527
0555
04FF
046D
0410
0401
0412
042A
045E
04A8
04D9
04DF
04F3
0530
0514
03AA
008C
FCAB
F9CA
F911
FA0F
FB4B
FBAF
FB5D
FB1C
FB49
FB8C
FB83
FB46
FB2A
FB39
FB36
FB15
FB15
FB58
FB9E
FBA2
FB8E
FBB4
FBF6
FBD3
FB36
FABE
FAEC
FB5D
FB56
FB24
FC32
FF60
0384
0648
0687
0561
04B4
0504
0566
0519
0487
0471
04C8
04DC
0476
0429
046D
04E0
04D3
0447
03F2
043D
04C1
04E0
0496
046A
049E
04DF
04D0
049F
04B2
04C2
03C3
00FC
FD29
FA2A
F95F
FA63
FB8C
FBA3
FAF0
FA7A
FAA3
FAE4
FAD7
FADF
FB83
FC6B
FCA4
FBE3
FB10
FB27
FBEC
FC47
FBC6
FB29
FB37
FBA3
FB9A
FB14
FADC
FB53
FBD2
FBD4
FC23
FE18
01A8
04EB
0617
056B
04A9
04EF
05AC
05D4
0551
04E7
04F6
0510
04C0
043D
0404
0424
044B
0458
047A
04BB
04CA
0473
03FB
03D3
0409
044B
0471
04B7
0544
0594
04BC
0252
FEF9
FC02
FA6E
FA41
FAAD
FAE2
FABA
FA9A
FACC
FB21
FB43
FB33
FB3C
FB78
FB94
FB55
FB07
FB2B
FBAF
FBF8
FBB3
FB5B
FB8A
FC21
FC6D
FC18
FB7C
FAFD
FA83
FA17
FA92
FCEF
00CF
0449
05B6
0557
04C4
04EA
054A
0529
04C2
04CE
0545
055C
04C8
0443
0480
0522
053F
04BB
045A
0490
04CF
046E
03BE
03AC
0466
050C
04E9
047A
04B2
0570
0559
0357
FFE5
FCA6
FAD5
FA6C
FAA2
FAE8
FB35
FB95
FBD2
FBA8
FB2F
FAD4
FAE4
FB30
FB43
FAFB
FAC3
FB09
FB9A
FBCE
FB69
FAFC
FB29
FBC4
FC06
FB9D
FB18
FB0D
FB3C
FB27
FB44
FCD5
002F
03C2
057E
0510
0412
0402
049E
04BD
0424
03CF
045F
052A
0543
04CB
04A3
0508
0542
04CC
0430
0440
04ED
0561
0532
04D4
04C2
04C5
0478
0425
046A
050C
04C8
02A7
FF43
FC4E
FAFB
FB19
FBAE
FC15
FC3C
FC36
FBF7
FB90
FB44
FB42
FB68
FB68
FB30
FAFA
FB00
FB30
FB3E
FB04
FABA
FAC2
FB31
FBB0
FBD2
FB91
FB4E
FB44
FB3A
FAFE
FB26
FCBE
FFF9
037B
0573
0565
0483
0425
045C
0456
03E0
03BA
0461
052F
0538
049A
0453
04D8
0576
0564
04DC
04AE
04F7
04F9
044E
039E
03B0
0450
04AF
04AA
04F1
05B0
05C5
03DB
002B
FC8E
FAA9
FA7B
FADE
FB0A
FB20
FB63
FBA6
FBA2
FB7E
FB8E
FBC0
FBA2
FB0F
FA87
FA9D
FB3C
FBC4
FBD9
FBC0
FBE9
FC47
FC61
FBFC
FB6E
FB31
FB39
FAFD
FA60
FA41
FBD6
FF47
0325
0594
0600
0576
0542
0583
0568
0499
03CF
03D9
0481
04E5
04B5
0486
04D6
053B
04F9
0426
03A0
03DD
0452
0449
03E7
03D9
0446
04A4
04AD
04DC
0582
05C1
042C
0093
FCA2
FA59
FA26
FADB
FB46
FB48
FB5B
FB9C
FBBA
FB9C
FB88
FB9F
FB9A
FB46
FAF4
FB17
FB95
FBD6
FB9B
FB58
FB93
FC1C
FC46
FBDF
FB7C
FBAD
FC1C
FBEF
FB0E
FAA6
FC17
FF6B
030D
0536
056D
04A8
0411
03F9
0409
0413
0450
04D3
0532
04FE
0473
044C
04CE
055E
053E
0492
0435
0495
051D
04FD
043D
0399
037C
038F
0380
03A7
0460
04F9
03F6
00D0
FD03
FAD2
FB08
FC51
FCDD
FC3C
FB61
FB2B
FB6F
FB8E
FB56
FB14
FAFD
FAFA
FB00
FB2F
FB7D
FB90
FB39
FAD6
FAF6
FB93
FC13
FC1C
FC11
FC75
FCF9
FCC3
FBBC
FB28
FC7C
FFAC
0304
04CA
04D7
0454
043F
0483
0493
0458
043D
0475
04A6
047B
0431
044D
04D8
0540
050E
0489
0461
04C6
0528
04EB
0433
03AD
03B4
03F2
03F6
03E5
0427
0479
03BD
0120
FD54
FA44
F95E
FA4E
FB8D
FC03
FBD6
FBBC
FBF5
FC2F
FC2E
FC17
FC13
FBFE
FBAB
FB41
FB13
FB28
FB3F
FB3D
FB5B
FBB6
FBFE
FBEB
FBBE
FBED
FC49
FC00
FAD8
FA19
FB88
FF65
03C8
065B
0680
057E
04C9
04AB
049B
0455
0416
0404
03E3
0399
0386
0403
04C7
0522
04DA
046E
046D
04C3
04E5
0494
0420
03F6
041C
044C
0472
04BF
052E
0529
03D8
00F1
FD48
FA65
F95A
F9ED
FAE5
FB44
FB15
FB06
FB70
FBF2
FC10
FBD2
FB9D
FB9A
FB9B
FB86
FB8F
FBC9
FBE7
FBA4
FB46
FB4A
FBB1
FBEF
FBB2
FB56
FB55
FB7D
FB50
FB1C
FC11
FEDC
0286
053B
0614
05B7
0540
0511
04ED
04C5
04D7
0516
0510
04A1
044D
048C
0503
04EC
042B
037F
0393
042E
04A3
04B8
04BD
04DE
04CA
044F
03DB
0410
04D0
0519
03E2
010C
FD8B
FAC5
F9AC
FA2A
FB40
FBD8
FB99
FB09
FACA
FAE8
FAF6
FACB
FAB5
FAF5
FB58
FB92
FBB1
FBEC
FC24
FBFF
FB7F
FB25
FB48
FB96
FB96
FB60
FB73
FBCF
FBE7
FBAB
FC1F
FE4A
01C0
04C3
0600
05B6
0508
04A4
0472
045B
0498
0522
0575
053A
04D9
04DD
0519
04E2
042B
03C2
0448
0547
05B7
053E
0473
03FD
03E0
03E2
041E
04B3
052F
04C3
031D
00B8
FE54
FC65
FB1B
FA96
FAC3
FB27
FB3B
FB04
FAF8
FB47
FB83
FB49
FAD7
FAAE
FAE2
FB1A
FB30
FB5D
FBAD
FBC3
FB60
FAEB
FB04
FBA9
FC3C
FC58
FC38
FC12
FBB1
FB25
FB67
FD88
0130
0481
05E1
0585
04DF
04D8
0522
0533
0521
0533
053A
04E7
0483
049B
051B
053C
049C
03DC
03DA
0485
0509
04F2
04A9
049D
0496
0430
03A0
0377
03DC
046A
04CF
04F4
0486
02E5
0005
FCFF
FB3C
FAF8
FB24
FADB
FA69
FA87
FB20
FB70
FB29
FACC
FAD3
FB15
FB35
FB4E
FBA9
FC14
FC02
FB6E
FB06
FB38
FB9C
FBAB
FB91
FBD9
FC6D
FCA4
FC3B
FBB6
FB8E
FB83
FB4C
FB8F
FD65
00B4
03D2
053A
051A
04C2
04E7
052E
0535
053F
058D
05B9
053D
0466
0413
0477
04D1
0487
0403
03FA
0458
0474
041E
03D6
03F5
0433
0433
041A
0432
045D
045F
0487
0545
05F3
04EF
0186
FD42
FA8B
FA29
FAC9
FAEB
FA8D
FA87
FAFF
FB44
FB06
FAD4
FB1D
FB7C
FB6C
FB39
FB84
FC2E
FC73
FC0F
FBA3
FBBE
FC18
FC15
FBC2
FBA9
FBD8
FBC1
FB28
FA95
FA72
FA6E
FA50
FAF2
FD6C
015C
04C8
0616
05AB
051A
0522
053B
04EF
04B4
0502
056B
0535
0486
0428
0455
0471
0413
03AB
03C2
041C
041E
03D3
03DD
0461
04C8
04C0
04D0
055E
05D7
0588
04DD
04D3
0525
041A
00B1
FC70
F9FE
FA28
FB35
FB52
FAA4
FA63
FACF
FB16
FAE3
FAE3
FB81
FC11
FBD5
FB36
FB42
FC1A
FCBC
FC75
FBCC
FB91
FBAC
FB82
FB09
FAC0
FAC6
FABE
FA99
FAC2
FB4B
FB85
FB20
FB38
FD5C
015F
0507
0661
05BD
04DC
04B0
04CB
04AB
049E
04FF
0565
0530
0486
041E
0428
0422
03D0
03B6
042E
04B3
04AF
046C
049C
0529
0555
04F1
04BD
0527
0577
04E7
0410
042B
04E2
0425
00CA
FC82
FA21
FA66
FB80
FBAC
FB2B
FB28
FBB1
FBC7
FB20
FAB0
FB1F
FBC2
FBAD
FB28
FB2E
FBDE
FC51
FBF8
FB57
FB1D
FB32
FB13
FACD
FAD7
FB31
FB51
FB1F
FB2D
FBA8
FBD5
FB4E
FB36
FD2B
0106
048C
05C4
04FA
0405
03F3
044B
0466
047C
04EA
0554
052D
04B6
04A9
050A
051B
0481
03DB
03DA
044A
0490
04AA
0505
0579
0556
049E
0451
04ED
0581
0505
0411
0418
04F0
0472
0138
FCE3
FA87
FB0F
FC66
FC6B
FB65
FAE4
FB31
FB39
FA87
FA05
FA7A
FB4E
FB80
FB2A
FB30
FBC2
FC0F
FBA6
FB2D
FB4F
FBAB
FB8C
FB1B
FB03
FB4D
FB5F
FB1A
FB0E
FB6A
FB7F
FAF4
FAEE
FCF8
00CF
0437
0571
0509
04A3
04D1
04F0
04B6
04B6
0545
05CA
059E
050B
04D1
04F5
04DA
045E
0421
046E
04B5
048B
046E
04E0
0553
04EA
0403
03ED
04F1
05AC
0505
03FD
0454
05A4
0541
01A4
FCBE
F9EC
FA24
FB5B
FB82
FAC6
FA7C
FAE6
FB21
FACD
FAA7
FB2F
FBC1
FB94
FAFF
FAF6
FB98
FC14
FBE3
FB74
FB54
FB63
FB34
FAE9
FAFD
FB6B
FBA1
FB62
FB17
FAFD
FAB3
FA36
FAA5
FD31
0151
04C8
05ED
0556
04D2
052C
059A
0558
04C6
04A9
04F8
051C
04EE
04CD
04D1
04AD
044E
041A
044B
0486
047B
0486
0514
05A9
0561
0472
042A
050A
05D2
054B
0439
044F
055B
04EC
016B
FC94
F9B7
F9E3
FB17
FB47
FAC1
FADE
FB97
FBB8
FAFA
FA76
FAE9
FB9B
FB90
FAFD
FAD2
FB36
FB67
FB0B
FABA
FAE6
FB1C
FAE5
FAA9
FAF3
FB70
FB7A
FB4B
FB9F
FC49
FC25
FB02
FAAC
FD0C
017B
0518
05EE
04ED
0435
0479
04E4
04E1
04CD
04FB
0518
04E2
04B9
04FF
055F
054A
04F4
0505
056E
055E
04AD
045D
0519
05F5
05A0
045D
03B9
044E
04F0
0490
03ED
045D
054F
0470
00C5
FC6D
FA57
FAED
FBFE
FBC6
FAD2
FA97
FB3F
FBAA
FB3D
FAA0
FA99
FAF1
FAFA
FAAB
FA8C
FAD4
FB27
FB34
FB18
FB09
FB09
FB1C
FB62
FBC5
FBCB
FB38
FA9C
FABD
FB5C
FB5C
FA7A
FA39
FC60
00A2
0494
0629
05A5
04D1
04C6
051E
0528
04F5
04F3
0525
0543
0548
0556
0551
0511
04D4
0500
0561
0544
047E
03EC
0450
0526
0545
049F
0454
04EA
056A
0504
0494
055D
0694
05AE
018F
FC81
F9DD
FA51
FB88
FB75
FA99
FA7F
FB3D
FB9E
FB29
FAB2
FAE1
FB3D
FB13
FA91
FA69
FAB9
FB03
FB1C
FB55
FBAB
FB98
FB03
FAAA
FB03
FB70
FB30
FAAD
FADF
FB96
FB84
FA5A
F9E9
FC3A
00D6
04EB
065C
05C7
051D
052E
0551
04F7
0477
044D
046C
0491
04BB
04F5
0507
04C8
048D
04C6
053C
0543
04CE
04A5
0535
05C8
0589
04D7
04BF
0556
0583
04B4
03F7
0487
05AC
0515
01A4
FD17
FA37
F9ED
FABE
FB05
FAB6
FABA
FB54
FBD3
FBAB
FB29
FAE4
FAF8
FB18
FB1B
FB1D
FB2D
FB32
FB24
FB14
FAFA
FABA
FA66
FA44
FA71
FAAC
FAC6
FB05
FBAF
FC43
FBDA
FA99
FA3A
FC6A
00AD
0486
05ED
0545
047B
04AD
0543
054A
04CE
0486
04B7
0503
0523
0531
054A
0557
054E
0553
0561
0536
04C4
048C
04FA
059B
0593
04E9
0495
050E
0577
04F2
0425
0462
0564
0505
01CC
FD26
FA13
F9DF
FB0D
FBA5
FB74
FB72
FBCE
FBBF
FAFF
FA53
FA6A
FAE5
FAFE
FAAC
FA86
FAC2
FAF0
FAD4
FACC
FB24
FB88
FB88
FB4D
FB38
FB33
FAF4
FAB8
FB00
FB96
FB89
FAA2
FA53
FC5D
0082
0460
05EF
0584
04ED
0519
0563
0506
0451
0424
04B9
057D
05D5
05B5
0556
04E4
048C
0483
04C1
04EC
04CB
0499
049F
04B8
0494
045D
0494
053C
05A1
054D
04DC
052B
05CD
050D
01EE
FDAB
FAA2
F9EA
FA8B
FB0A
FB07
FB0E
FB53
FB66
FB08
FAAB
FABF
FB08
FB0E
FADA
FAE7
FB5A
FBD5
FC02
FBF2
FBCE
FB8A
FB1D
FAD2
FAEA
FB1D
FAF1
FA87
FA82
FAF3
FB0E
FA75
FA52
FC45
0038
0408
05B4
056B
04E3
0512
055E
050F
0494
04C1
0574
05C2
054C
04AC
047C
049B
04A1
0497
04BD
04EE
04B8
042D
03EF
0458
04FC
054E
055A
0567
055F
0519
04F3
056A
05FB
0527
021A
FE01
FB14
FA5A
FAE2
FB49
FB47
FB60
FBA2
FB83
FADD
FA46
FA4B
FAC1
FB24
FB5A
FBA2
FBF5
FBF2
FB76
FAE5
FAB0
FAD5
FB20
FB7D
FBCA
FBA6
FAE4
FA16
FA16
FAE6
FB8C
FB69
FB52
FCBC
FFD3
0301
04A6
04BC
0475
0492
04C6
04A8
047E
04CA
0570
05D0
059C
052E
04F0
04D1
048D
0432
0409
042B
0475
04C9
0526
0573
0581
0546
04F8
04C4
04AD
04B3
04F8
055B
0523
0385
00AB
FDDD
FC46
FBE3
FBD9
FBAD
FB95
FBC3
FBD7
FB68
FABB
FA7A
FAC8
FB1D
FB12
FAE9
FB0A
FB59
FB6D
FB3F
FB28
FB45
FB51
FB21
FAF3
FAFF
FB16
FAFD
FAFA
FB7A
FC2E
FC18
FAF8
FA2C
FB86
FF32
034D
05B4
05F2
0535
04B6
04A2
0487
044B
0448
04AC
051E
052D
04DF
0498
049E
04CF
04DD
04BB
04A9
04D5
0513
0510
04CE
049D
04AA
04B4
046A
03FD
0405
04C2
05B6
0626
05E3
054E
048C
0328
00C4
FDE1
FBA0
FAB6
FACF
FB0D
FAFB
FAD0
FAF0
FB5B
FBB4
FBB5
FB70
FB2E
FB24
FB48
FB68
FB60
FB3D
FB2F
FB49
FB65
FB4D
FB01
FAC6
FAEC
FB7A
FC04
FBF2
FB1F
FA31
FA16
FB06
FC19
FC3A
FB81
FB60
FD2A
008B
03BC
0550
056C
052F
0539
0541
04E7
0468
044F
04B0
0512
0514
04D3
04A3
0497
0490
0490
04BF
0511
0528
04C1
041D
03D6
0433
04D9
052C
0501
04BA
04B5
04CF
04B6
0485
04B8
054B
0543
0373
FFEA
FC45
FA4C
FA5A
FB37
FB91
FB3A
FAEE
FB28
FB92
FB97
FB29
FAC0
FAC0
FB0E
FB45
FB34
FB0E
FB21
FB7E
FBEA
FC1A
FBE3
FB51
FAB0
FA73
FADA
FB95
FBED
FB7A
FAB3
FA7B
FB09
FB90
FB5B
FB18
FC56
FF8F
0338
053F
0533
0471
0452
04C2
04DF
047A
0440
0498
0512
052D
0519
053C
0567
0517
0460
03F7
0442
04CF
04F6
04BC
04AA
04EE
0518
04CB
0460
0476
0512
0587
0542
047B
0404
045F
0501
0482
01F1
FE10
FAF1
FA10
FAF1
FBD3
FBB2
FB25
FB2D
FBB6
FBCB
FB13
FA5B
FA6E
FB11
FB82
FB8C
FB88
FB93
FB6B
FB11
FAF7
FB4B
FB88
FB28
FA86
FA87
FB51
FBFA
FBC2
FB1F
FB0D
FB9A
FBC9
FB05
FA26
FAC1
FD78
013B
042C
053B
04E0
0467
049A
0534
0571
050E
048C
047F
04D7
0507
04D3
0495
049F
04C6
04B8
047F
0465
0477
0489
049F
04F0
056E
0595
0511
045B
0446
04DE
0547
04E7
0458
04A0
05A4
05E7
040A
0061
FCBD
FABF
FA8A
FB06
FB33
FAFD
FAE4
FB1F
FB61
FB54
FB12
FAF2
FB14
FB3D
FB3D
FB39
FB66
FBA2
FB9B
FB5C
FB4C
FB91
FBC6
FB90
FB35
FB3D
FB9A
FB9F
FAF4
FA37
FA3C
FADF
FB1B
FA78
FA00
FB51
FEBF
02C3
055A
05CA
0510
04A5
0503
0571
0519
042F
03BA
045B
0584
061B
05AC
04C3
0429
040E
0420
042E
0456
049B
04C2
04B4
04A7
04B7
04A9
045C
0430
048F
0533
055D
04EF
04C2
0575
0632
0542
0208
FE04
FB61
FAD7
FB52
FB7C
FB21
FAE6
FB22
FB6F
FB4A
FAD1
FAA0
FAFD
FB79
FB7C
FB0F
FACC
FB17
FB9B
FBBE
FB70
FB38
FB69
FB9E
FB5C
FAEA
FB00
FBA7
FC06
FBA1
FB25
FB72
FC23
FBEF
FAA5
FA04
FBEC
0002
03D0
055B
0502
047D
04B4
051C
04F7
0466
0416
0460
050C
05A8
05E3
0592
04C9
03F1
039D
0406
04CD
0556
055D
0516
04D0
04A9
0494
0481
047A
0490
04B2
049D
043B
03F5
0466
056F
05DB
0450
00D3
FD15
FAF0
FAB0
FB14
FAF7
FA7A
FA6D
FB02
FB97
FBA5
FB62
FB51
FB83
FB9A
FB66
FB27
FB2D
FB5E
FB5F
FB20
FAFD
FB3A
FB9C
FBB8
FB87
FB72
FBB3
FBE3
FB7A
FAA5
FA4A
FAD6
FB7F
FB3D
FA7E
FB1B
FE3E
02A4
05AF
061E
0521
04A7
0526
0595
0535
048E
0470
04BF
04CB
0470
043F
0493
0509
051A
04D6
04B6
04EC
0520
04F7
0483
0425
040E
042C
0463
04B0
04FA
050D
04CA
0467
0462
04FC
05A8
0529
02A6
FEC9
FB73
FA10
FA57
FAE0
FAD4
FA9E
FAF5
FBB5
FC16
FBCF
FB64
FB45
FB38
FAF1
FABF
FB11
FBA6
FBBC
FB29
FAAE
FAEF
FB88
FB96
FB01
FAA6
FB15
FBB6
FB97
FAC1
FA3B
FAAC
FB7C
FB9F
FB05
FAF2
FCC3
006A
0436
0646
062C
051F
0499
04E3
0529
04CA
0436
044C
050F
0598
054A
049F
0473
04D3
050A
04BE
0473
04B9
054A
0566
04E2
045D
045C
04A1
04BB
04C8
0531
05CB
05DF
053C
04B5
0502
0572
0453
00FA
FCDA
FA37
F9E5
FAC2
FB44
FB11
FAD3
FAF4
FB27
FB15
FAED
FAFD
FB24
FB0F
FAD5
FADF
FB37
FB53
FADB
FA4B
FA76
FB65
FC2C
FC02
FB37
FAC1
FB02
FB6B
FB5B
FAFA
FAEC
FB4C
FB68
FAB2
F9D6
FA6F
FD6D
01D0
0550
0667
05A4
04CF
04F6
058A
0582
04DB
0489
050C
05B1
0593
04D3
045D
04A4
0527
054B
0530
054E
0595
0577
04D1
043F
0449
04A7
04BC
0480
0478
04CE
0505
04C2
047C
04E3
05B7
0599
0364
FF87
FBD6
F9F0
FA04
FAF3
FB84
FB53
FAD7
FAA6
FAD2
FB02
FAF7
FAD1
FAC7
FADC
FAF1
FB07
FB31
FB57
FB3B
FAE2
FAB6
FB08
FB86
FB94
FB22
FACF
FB0A
FB70
FB64
FB0F
FB27
FBBA
FBD6
FAE9
FA11
FB51
FF27
0393
05F6
05B9
049A
0473
0549
05D0
0555
0487
0465
04FA
0580
0579
0533
052D
0563
0572
052F
04D8
04A9
048A
0452
042A
046F
051D
05A7
058B
04F5
0480
0473
0476
0444
0444
04FA
05E2
0562
0269
FDF8
FA85
F99C
FA7F
FB4A
FB1F
FAB1
FAD9
FB53
FB49
FAA7
FA36
FA75
FAE8
FAE7
FA94
FA91
FAFF
FB4D
FB1F
FAE1
FB18
FB96
FBAF
FB40
FAEB
FB29
FB9A
FB96
FB35
FB27
FB9B
FBC5
FAED
F9BC
FA02
FCE2
0167
052D
067C
05B3
0498
0475
0513
0572
052C
04D6
050C
0592
05A8
051F
0492
048E
04E5
051B
052C
0571
05E1
05E8
0541
048E
0496
052A
0556
04B6
0410
043D
04EF
0531
04D9
04C3
0557
0578
039E
FFDA
FC25
FA73
FAC3
FB77
FB4C
FA7C
F9FF
FA39
FAB8
FAFC
FB09
FB37
FB93
FBCE
FBA5
FB3C
FAEB
FAD8
FAE7
FAFE
FB23
FB59
FB69
FB1A
FA93
FA55
FAB2
FB54
FBA2
FB80
FB5E
FB70
FB40
FA78
F9EA
FB28
FEB1
02EC
0574
057C
0482
0468
0569
0642
060F
055B
0523
0574
0588
0507
0480
0489
04DF
04D9
0474
0454
04C0
0519
04AF
03CE
0373
0404
04CE
04FB
04A3
0484
04D9
0516
04DE
04B9
054F
0617
057E
02A3
FEA0
FBA0
FAC4
FB3C
FB81
FB09
FA7B
FA80
FAD9
FADE
FA74
FA2B
FA65
FAD6
FAF8
FAC9
FABF
FB0D
FB5A
FB4E
FB1E
FB47
FBCB
FC18
FBD3
FB62
FB5F
FBB8
FBD3
FB88
FB70
FBED
FC53
FBB2
FA6A
FA47
FC9E
0099
03E4
0510
04C8
0494
04FD
0561
0537
04D1
04C1
0508
053F
053E
0549
0582
05AA
0585
053D
0527
053E
052F
04D6
047A
0477
04D1
052D
052C
04BD
042D
03DF
03F3
043C
047D
04AD
04D2
0492
0340
0097
FD6F
FB3B
FAB6
FB2D
FB69
FB07
FA9B
FAAB
FAF5
FAF6
FAB9
FAB8
FB09
FB29
FAC1
FA36
FA23
FA7D
FAAE
FA7E
FA66
FACE
FB60
FB77
FB15
FAEF
FB6B
FBFD
FBE3
FB43
FB01
FB77
FBDA
FB66
FACA
FBB6
FED2
02A0
04E2
04E5
040A
03EA
049E
0526
0511
04F9
056A
05F8
05E4
0543
04E1
051C
057C
0584
056F
05B4
0616
05E3
050C
046C
04A8
0540
0545
04A1
042C
0465
04C6
049B
0415
0400
048C
0504
04D5
046A
046E
0491
039E
00FC
FDA0
FB32
FA73
FAC7
FB34
FB63
FB8A
FBB4
FB8F
FAF9
FA52
FA0E
FA26
FA3D
FA33
FA4D
FABD
FB42
FB6F
FB36
FAEA
FAC5
FAAD
FA82
FA6C
FAAF
FB39
FBAE
FBE1
FBED
FBE2
FBA5
FB48
FB32
FB94
FBE1
FB63
FA70
FA8F
FCE6
00A9
03AD
04A2
044A
043F
0501
05B1
058B
04EA
04AC
050B
057D
0588
0542
04F8
04C3
04AF
04E6
056F
05D9
059E
04DB
0447
0457
04B5
04CB
0497
049C
0505
054B
04FB
0475
047D
050F
0544
0497
03D1
0412
0515
050B
0295
FE8A
FB47
FA47
FADD
FB6A
FB45
FAF3
FAEE
FAE5
FA7D
FA19
FA63
FB43
FBE4
FBC7
FB5A
FB40
FB6B
FB54
FAE8
FAA8
FADE
FB25
FB0F
FAD8
FB0F
FBA3
FBE4
FB6F
FABA
FA73
FA9F
FAD4
FB08
FB99
FC6A
FC97
FB9B
FA80
FB32
FE64
028C
055B
05FD
0589
055E
05A4
05A2
0513
048D
0498
04F6
0511
04CA
047C
0455
042B
03FB
0424
04D9
0599
05AB
0503
045C
0452
04B2
04F4
0500
0522
0556
0534
04B0
046C
04D8
0564
0527
0448
03FC
04C8
0544
036E
FF2D
FADE
F904
F9C7
FB36
FBA6
FB33
FAE3
FB16
FB4C
FB1F
FAD6
FAD5
FB13
FB56
FBA2
FC0B
FC4C
FBFE
FB4C
FAF3
FB50
FBCA
FB8F
FAB8
FA3E
FAAA
FB5A
FB67
FADF
FAA4
FB0C
FB67
FB14
FA93
FADF
FBE5
FC74
FBF7
FBA8
FD4B
00E7
0469
05D1
0545
0488
04C4
0571
0583
04ED
0484
04BA
0518
0504
0492
043E
0437
0444
0449
0470
04C7
0503
04E3
0498
0485
04B4
04D8
04DA
04FC
0552
0575
0507
045C
0427
047C
049D
0415
0394
041F
0558
0555
02A2
FE2C
FAA3
F9CB
FAE7
FBDA
FB8D
FAB6
FA83
FB1D
FBBA
FBC6
FB71
FB35
FB3A
FB58
FB70
FB77
FB59
FB03
FAA2
FA8A
FAD6
FB43
FB84
FB92
FB89
FB62
FB17
FAEA
FB37
FBE1
FC37
FBCE
FB2F
FB43
FC02
FC45
FB5A
FA5D
FB64
FF0C
036B
05DC
05A0
0453
03D4
045C
04DB
04AE
0453
0475
04F0
052A
04FB
04CB
04DC
04FA
04EF
04ED
052C
056E
0541
04B4
0461
04A3
0512
0515
04B3
0475
048C
0492
0441
03FC
043E
04C9
04E7
0486
0470
0502
0528
0351
FF76
FBA2
F9FA
FA94
FBA7
FBBD
FB19
FAD2
FB34
FB8A
FB4E
FAE3
FADB
FB1B
FB1C
FAD1
FABE
FB29
FBA2
FBA0
FB48
FB29
FB6B
FB9B
FB66
FB19
FB24
FB6E
FB83
FB47
FB1A
FB2E
FB2B
FACC
FA73
FAAC
FB3E
FB54
FAD7
FB1A
FD8B
01C2
057B
06BA
05B5
0451
0408
04B5
0560
0591
058B
058F
057D
0532
04DA
04AC
0492
045C
0428
043D
0497
04D0
04AC
0464
044C
045F
045F
0457
049D
053B
05B9
05B8
057D
0585
05B1
055A
0465
03BC
0431
0514
0484
018C
FD78
FAAE
FA41
FB18
FB77
FADE
FA1C
F9F4
FA3B
FA67
FA6B
FAA5
FB29
FBA2
FBC7
FBB2
FB96
FB6E
FB2C
FB05
FB41
FBBF
FC03
FBD3
FB7D
FB5F
FB5D
FB19
FA9F
FA65
FA98
FAD8
FAD4
FAE5
FB89
FC60
FC59
FB31
FA61
FBCD
FF8E
038F
059B
0582
04DE
04FE
05A8
05E8
0587
051E
0511
050D
04AD
0430
0425
049B
050E
0515
04E0
04D4
04FD
050D
04DA
0493
0473
048A
04CC
052B
057C
0573
04FE
047D
046E
04C1
04D2
0452
03D7
0433
0527
0535
0320
FF6E
FC12
FA94
FABC
FB37
FB29
FACB
FAAC
FAD4
FAE3
FABD
FAB6
FAFF
FB5E
FB7D
FB61
FB48
FB3C
FB0D
FAB7
FA8A
FAC0
FB23
FB45
FB17
FAF2
FB19
FB61
FB7C
FB63
FB46
FB30
FB10
FB0D
FB79
FC33
FC76
FBB5
FAAB
FB03
FD9D
0163
0439
050C
04A8
047C
04FD
0588
0592
0558
054D
055B
0514
047A
041E
0465
0501
0563
056E
0578
05AC
05C2
0571
04E3
0486
0489
04C2
0500
053F
056A
0549
04D8
0478
0484
04C2
04A6
042C
0418
04E2
059F
0494
012E
FD07
FA7E
FA59
FB34
FB59
FAA9
FA4D
FAE7
FBBA
FBBD
FB02
FA7E
FAB7
FB33
FB4B
FB12
FB08
FB3F
FB48
FAF2
FAA8
FAD5
FB43
FB60
FB06
FAA4
FA99
FAC8
FAEB
FAF7
FAFF
FAE7
FA9A
FA66
FAB7
FB58
FB7D
FAEA
FAC5
FC91
004A
03FB
05A2
0531
0452
0458
0508
057A
0579
058A
05D5
05C9
050B
0427
03F4
0473
04DF
04C4
0485
04AA
0508
050B
04A4
0472
04E1
0590
05CE
057D
051D
0512
053F
0562
056D
0561
0518
049B
047B
0538
062F
05B6
02C4
FE6C
FB1E
FA43
FAFA
FB69
FAE1
FA40
FA62
FAF8
FB2D
FAF4
FB03
FBA4
FC37
FC10
FB69
FB03
FB18
FB2C
FAEE
FAB2
FADA
FB24
FB10
FAB0
FA91
FAD9
FAF5
FA81
F9FC
FA2C
FAF3
FB66
FB22
FADE
FB4A
FBDE
FB8F
FAA4
FAF3
FDCE
0226
0563
0612
052A
048B
04D5
053E
0512
049C
047D
04B9
04D9
04B5
049A
04AE
04B3
0480
045F
04A7
0529
0566
0545
053A
0592
05F9
05ED
0572
050F
050D
0527
050B
04D9
04D4
04DA
048F
0423
044A
052C
059C
0404
0049
FC52
FA50
FAA1
FBB2
FBE9
FB3A
FAB6
FAF1
FB6C
FB7B
FB34
FB2C
FB91
FBEF
FBDC
FB87
FB59
FB5D
FB3F
FADB
FA74
FA5D
FA90
FACB
FAE4
FADC
FAC3
FAB3
FAD3
FB30
FB87
FB7B
FB1E
FB02
FB79
FBF3
FB93
FA8E
FA7D
FCCC
00F0
049C
05F3
053E
0445
0448
04F4
054F
0517
04D8
04F9
052A
04F5
046B
0411
0437
04A7
04F7
04F8
04C1
047B
044B
0458
04B0
0521
0557
0535
04FA
04EF
0512
0526
050F
04F3
04EC
04DE
04AE
0497
04E6
054B
04C2
0288
FF1E
FC13
FA92
FA67
FA83
FA57
FA42
FABB
FB75
FBB6
FB54
FAE7
FAEF
FB32
FB2C
FAE0
FAD6
FB4D
FBD8
FBF3
FBA8
FB6A
FB67
FB5D
FB22
FAEF
FB05
FB44
FB5E
FB52
FB5A
FB7C
FB78
FB34
FAF1
FAD7
FA9E
FA1A
F9FB
FB79
FED9
02B0
0512
056F
04E5
04C2
0520
0546
04F3
04B9
050E
0591
0594
050F
04A2
04B0
04EA
04D6
047E
0453
0485
04D0
04E1
04B8
048B
0477
047F
04A4
04D6
04DA
0485
041B
0423
04B3
0529
04F4
0471
0496
0588
05F2
0442
008C
FCBE
FACA
FAD7
FB83
FBA2
FB44
FB0E
FB27
FB33
FB16
FB1C
FB5F
FB7B
FB1C
FA99
FA92
FB0C
FB59
FB09
FA84
FA80
FB08
FB8A
FBA0
FB86
FB98
FBC1
FBAE
FB5B
FB13
FAFA
FAF7
FB0C
FB73
FC19
FC6D
FC0F
FB71
FB54
FBAB
FB91
FABF
FA7A
FC63
0059
0428
05BA
051E
0418
03F5
0479
04D0
04D3
04F2
0544
0559
04FB
049A
04B3
0524
0569
0549
0501
04CA
04A3
0492
04C0
051F
0547
04EC
0461
0443
04A2
04DD
0484
03F6
03E2
0449
0489
044F
0406
0427
0476
0472
0447
04A6
0583
0581
034A
FF54
FBC4
FA57
FAC5
FB71
FB5B
FAE6
FAD2
FB1D
FB31
FAE4
FAA8
FAD5
FB25
FB2A
FAED
FAD5
FB0B
FB54
FB81
FBA7
FBD5
FBD5
FB83
FB2B
FB3D
FBA8
FBE0
FB99
FB37
FB40
FB95
FBA7
FB52
FB19
FB5B
FBBE
FBBF
FB7E
FB7A
FBA7
FB6B
FACD
FB1A
FD9D
01C3
0539
0635
053B
0440
0469
0530
0592
0563
0527
0523
051E
04FA
04EC
0508
04FE
049B
0434
0440
04A2
04CB
0487
043D
044A
0479
046C
0445
047B
0512
0571
0530
04A2
0460
047F
04A1
04A7
04CE
0519
0522
04C6
049E
052D
05BA
04A8
0155
FD35
FA97
FA54
FB39
FBA7
FB42
FAD3
FAE1
FB1A
FB03
FAB5
FA9E
FAD2
FB03
FB14
FB3D
FB9D
FBEB
FBDC
FB93
FB7B
FBAA
FBD1
FBAE
FB71
FB66
FB87
FB8D
FB66
FB4A
FB5A
FB6E
FB59
FB35
FB30
FB32
FB0B
FAE2
FB17
FB91
FB9A
FADC
FA51
FB9D
FF2C
034E
05BA
05CB
04DE
048A
04F4
053D
0503
04CF
051C
0591
058A
050C
04AF
04B7
04CA
0496
0456
046D
04C4
04F4
04E5
04DE
0502
0510
04D6
048E
0488
04A6
0491
0452
0451
04A7
04E2
04B5
047D
04AB
04F5
04B9
0420
042F
053D
05E0
042F
0022
FC00
FA10
FA59
FB19
FB11
FAA0
FAA7
FB23
FB65
FB30
FAF8
FB10
FB32
FB0C
FADA
FB02
FB5E
FB6E
FB1C
FAE5
FB1D
FB75
FB77
FB33
FB18
FB3C
FB3E
FAE9
FA9F
FACE
FB4A
FB95
FB93
FB98
FBC3
FBC4
FB78
FB51
FBB5
FC29
FBCD
FACA
FAB7
FCFF
0100
0471
05AB
0531
04AF
04F3
0564
054B
04E5
04DE
053D
056D
052B
04E8
050D
0554
0538
04C4
0487
04B7
04ED
04C8
0489
04A4
0507
0532
04FB
04C6
04DD
04FF
04CA
0469
0454
0493
04AA
0469
043A
046B
049B
0456
040C
048D
0589
0543
0279
FE3E
FB27
FA87
FB38
FB61
FAB4
FA51
FACB
FB58
FB21
FA88
FA89
FB37
FBA6
FB50
FACD
FADB
FB48
FB5C
FAFC
FAC2
FB02
FB57
FB58
FB40
FB7A
FBD8
FBCB
FB49
FAF1
FB1D
FB62
FB48
FB15
FB51
FBD3
FBE4
FB65
FB24
FBA0
FC18
FB8A
FA85
FB03
FE1C
0263
0540
05B3
0507
04E6
056F
05A6
052A
04AE
04D5
0545
0552
0504
04F1
053F
056F
0528
04CC
04D6
051D
0509
047C
0408
041C
0478
049C
0484
0487
04B2
04AD
0466
044D
04AE
051C
04FA
046B
0434
0499
04F3
04B1
044F
0494
0510
041D
00E9
FCDB
FA59
FA34
FB05
FB28
FA98
FA64
FAE8
FB5E
FB2E
FACB
FAE6
FB55
FB60
FAF9
FAD8
FB57
FBD8
FBAD
FB1F
FB00
FB70
FBBD
FB82
FB38
FB6F
FBDB
FBCA
FB40
FB03
FB75
FBFD
FBF0
FB84
FB64
FBA1
FBB2
FB6C
FB49
FB82
FB81
FAE2
FA98
FC41
0009
03FE
05F5
05C1
04FC
04EB
054A
054B
04F0
04DE
0537
0561
04FD
0481
0483
04DD
04F7
04B6
049B
04E5
0524
04E3
045B
0427
046C
04B3
04A9
0490
04C4
051E
0530
04E6
049F
0498
049F
0489
0481
04B5
04E0
04A3
0443
0477
053B
053F
0328
FF55
FBDC
FA7D
FAF0
FB88
FB46
FAB2
FAB2
FB37
FB79
FB31
FAE7
FB0E
FB5B
FB4E
FB02
FB06
FB78
FBD3
FBAC
FB4C
FB35
FB6F
FB91
FB70
FB4D
FB61
FB82
FB77
FB58
FB5C
FB73
FB5E
FB30
FB41
FB93
FBB1
FB63
FB24
FB72
FBE6
FBA2
FACC
FAFC
FD88
01A7
04F5
05E5
0536
04A6
04D5
0504
049F
0428
0458
04FB
0544
04F2
049D
04BC
0500
04E8
0491
047C
04BB
04E3
04BA
0490
04AF
04E2
04CA
0482
047C
04CB
0500
04D2
048A
048D
04BA
04B2
047D
047F
04BB
04B4
0438
03ED
0474
0539
04A2
01DB
FDFD
FB13
FA1F
FA74
FAE0
FAF1
FAEF
FB07
FB0D
FAF8
FB11
FB7C
FBD8
FBB4
FB37
FAF9
FB38
FB84
FB60
FAF3
FACA
FB0D
FB4F
FB3A
FB0B
FB2E
FB88
FB91
FB1E
FAB5
FAE3
FB7A
FBCD
FB97
FB42
FB3C
FB6E
FB88
FB86
FB89
FB69
FAF7
FABA
FBE2
FEFA
02E0
0592
0622
057D
0516
0547
0562
04FC
0480
0476
04C9
0508
0519
052E
0541
0514
04C5
04D8
0565
05BB
0535
0442
03FA
04B2
0584
0577
04BD
044F
048B
04DD
04C3
0491
04CC
053B
053B
04BE
0469
0499
04E0
04C9
049F
04D7
04EF
039C
0073
FCD5
FAAA
FA6A
FAE7
FAF4
FAA2
FAA7
FB18
FB51
FAFD
FA99
FAC0
FB4E
FB99
FB52
FAD4
FA97
FAAE
FAE8
FB2C
FB6F
FB7D
FB2E
FABD
FAA7
FB06
FB60
FB42
FAE1
FAD4
FB38
FB8B
FB6E
FB36
FB61
FBC5
FBC8
FB57
FB1C
FB6E
FBB7
FB5A
FB06
FC49
FF9F
037C
05C4
05F4
0553
0524
055A
054C
04FB
04F3
0543
0550
04D3
045F
0498
053F
0581
0519
04A9
04CF
0559
05A3
0572
051A
04E5
04D1
04D0
04F7
0530
0523
04B0
0447
0473
0507
053F
04C5
0432
0439
04A4
04B7
0462
0472
0525
0536
0311
FEF8
FB30
F9BE
FA67
FB56
FB53
FAB6
FA61
FA82
FAB3
FACD
FAFD
FB34
FB1D
FACB
FAC6
FB3D
FB98
FB4B
FAB4
FAA4
FB2F
FB91
FB45
FABB
FAA1
FAE7
FAF6
FAAE
FA98
FB00
FB79
FB8B
FB70
FB9B
FBE4
FBC5
FB52
FB42
FBCB
FC20
FB81
FAA3
FB47
FE42
024B
052A
05DC
053A
04B6
04EC
0572
05A1
054D
04CD
049B
04E5
0562
058F
052E
048E
0450
04B5
0553
0582
0521
04B1
04A7
04E6
0505
04F1
0501
0559
058F
052C
046A
0417
049D
0569
0592
04E9
041B
03CA
03F2
0446
04B9
053E
053C
03D4
00EB
FD9D
FB5A
FA9E
FAB8
FACA
FAAB
FAB4
FB14
FB87
FBA9
FB5E
FAE0
FA9B
FAD0
FB4F
FB8E
FB3B
FAAC
FA8C
FB0B
FB98
FB91
FB0C
FAB1
FAD6
FB1F
FB18
FAE5
FAFE
FB66
FB96
FB41
FADB
FB0C
FBC1
FC30
FBCD
FB01
FAA8
FAFF
FB6B
FB5F
FB44
FC33
FEC0
0231
0503
0627
05CA
04F2
0485
04A3
04E3
04FB
050F
054D
057C
0533
047F
040B
0466
0533
057B
04D5
0400
0406
04EB
05A7
0570
04A0
0426
0459
04CF
050F
0517
050D
04E6
048F
0447
046C
04EF
0541
04FB
0469
0444
04DE
05AB
0589
0394
0000
FC41
FA15
FA11
FB20
FBB4
FB53
FACC
FAE8
FB58
FB4A
FAAC
FA5A
FAE0
FB9F
FB99
FAD8
FA6D
FB0C
FC17
FC5F
FBA0
FAC4
FABF
FB71
FBEA
FB93
FAD1
FA76
FAD3
FB7A
FBCF
FB97
FB19
FACD
FAFB
FB7F
FBE3
FBCA
FB51
FAF3
FB03
FB5C
FBA5
FBB1
FB85
FB36
FB0A
FBAD
FDC6
0117
043A
05C3
05A5
0520
0535
05A5
05A6
052A
04E3
0521
055F
0512
0488
0487
052D
05AB
0549
0456
03D9
045F
0565
05F2
0596
04C6
0459
04B4
0564
0593
04E9
03F8
03AC
0451
0539
057B
04EA
0441
0446
04E6
0550
04F7
0436
03D0
0409
047C
04C3
04DB
04B4
03C2
017F
FE52
FB8B
FA31
FA21
FA7B
FAC3
FB15
FB69
FB4E
FAA4
FA1D
FA70
FB55
FBCE
FB66
FABE
FAAD
FB36
FBA1
FB75
FAF2
FAA9
FAD7
FB50
FBB2
FB9E
FB03
FA5D
FA6A
FB48
FC17
FBE8
FAF6
FA82
FB44
FC76
FCBA
FBCA
FAC3
FABB
FB79
FBF4
FBB7
FB45
FB27
FB39
FB2F
FB76
FCED
FFBA
02D2
04F3
05B9
05A2
0542
04DF
04B4
0502
05A2
05ED
056B
048A
0436
04B9
0561
0576
0508
04A7
0499
04BC
04EB
0516
050E
04B5
045D
048F
0537
0579
04C1
03BB
03B0
04CA
05B8
0556
042B
03B6
0477
0570
058B
04E2
045A
0468
04B2
04CB
04CC
04F6
0511
0472
02AD
FFFA
FD17
FAE1
F9EB
FA2C
FAED
FB4A
FAF3
FA63
FA3F
FA9D
FB06
FB1B
FB08
FB1F
FB55
FB55
FB14
FAF5
FB3B
FB94
FB80
FB12
FADD
FB23
FB76
FB66
FB2A
FB40
FB99
FB9B
FB13
FAA2
FAF3
FBBC
FC0A
FB81
FACF
FABD
FB3B
FBA3
FBA5
FB7D
FB67
FB4F
FB1C
FAFC
FB43
FC39
FE09
00B1
03A7
05D1
0655
0587
04B0
04AB
0515
0514
04AC
04A9
054F
05C2
052A
040A
03C5
04D0
05FC
05E0
0496
0395
03EA
0517
05E2
05BB
050F
0475
042C
0444
04C7
0567
0581
04DB
0416
03FB
0486
04F6
04DF
04A1
04AF
04DA
04B2
0465
0491
053D
05A7
0543
0458
032E
015E
FE96
FBB2
FA31
FA6B
FB17
FAFC
FA82
FADF
FC03
FC6D
FB4C
F9E4
FA0B
FBB6
FCF6
FC5E
FAAD
F9BC
FA5B
FBA9
FC4E
FBE2
FB03
FA81
FAB2
FB55
FBDA
FBD1
FB56
FB02
FB42
FBC2
FBCC
FB41
FAD0
FB10
FBA9
FBBC
FB1D
FA9D
FAF5
FBC8
FC1A
FB96
FAE6
FAB9
FB04
FB97
FCEC
FF94
02EB
0537
0581
04C2
049C
054D
05A0
04DC
03EB
0410
0516
0597
04F2
041B
0433
0500
056F
0513
0488
0479
04DF
0548
0563
0520
04A8
0459
0498
053E
0589
04F5
0416
0407
04EA
0595
0522
0434
041A
04FD
05B8
0569
048B
0422
0468
04C8
04EC
051A
0556
04C6
028F
FF1C
FBFE
FA7B
FA7C
FB07
FB66
FB88
FB93
FB77
FB21
FAD2
FAF0
FB71
FBC2
FB79
FAEE
FADD
FB67
FBDE
FBA2
FAF0
FA8A
FAD0
FB60
FBA0
FB62
FAEF
FAAF
FAD6
FB4E
FBB4
FB91
FAE8
FA6E
FAD0
FBC0
FC23
FB7C
FA94
FA7A
FB2C
FBCC
FBD4
FB86
FB36
FAC7
FA46
FA75
FC27
FF14
01F1
03D0
04DE
0591
05C6
053A
0462
041F
0494
0501
04D8
0478
048B
0503
052A
04AD
0421
0449
051F
05DA
05CC
0503
0432
0416
04DA
05D1
05FB
050E
03E1
03A3
048A
059F
05CE
050D
0438
0406
0463
04D6
0523
0544
0511
0466
03A8
03B0
04D6
0639
0669
04CA
0221
FFA2
FDC5
FC43
FAF7
FA48
FA82
FB2F
FB84
FB55
FB24
FB42
FB4F
FADC
FA44
FA57
FB43
FC2C
FC15
FB05
FA09
FA1B
FB2B
FC37
FC45
FB45
FA27
FA01
FAFC
FC18
FC2D
FB36
FA59
FA89
FB68
FBDA
FB85
FB25
FB60
FBC3
FB7C
FABC
FAA5
FBB0
FCC6
FC83
FB03
F9DF
FA53
FC17
FE2F
004B
02AD
04FF
0631
05CC
04C6
0470
04EC
0542
04E7
047A
04C3
0578
0595
04CA
03F8
041C
0519
05E3
05B0
04BA
03F5
0424
0529
0603
05B8
046E
0374
03E6
054E
060E
0545
03EE
03AF
04C7
05C9
057B
0464
03F3
048F
0529
04C9
03DC
0395
0456
0553
059E
0512
03F1
0221
FF66
FC4A
FA22
F9D1
FABA
FB6E
FB45
FAD6
FADB
FB2E
FB36
FAEF
FAFB
FB9B
FC29
FBDF
FAE6
FA43
FAA1
FB95
FC1B
FBA6
FA99
F9E8
FA4A
FB89
FC82
FC2D
FAD5
F9F8
FA9C
FC03
FC81
FB92
FA82
FAB7
FBDE
FC6C
FBB9
FACE
FADE
FBAC
FC18
FBB5
FB23
FAF2
FB06
FB4E
FC68
FEEA
0242
04EB
05E6
05A0
0526
04EA
04B1
046B
0476
04F2
0563
053A
049C
0439
0476
04FD
052E
04DB
0466
0450
04C0
0569
05C8
057F
04BD
0436
0484
055A
05B3
04F1
03C4
0377
0464
0570
055F
0458
03A8
0413
04F1
0529
0498
0406
03FB
043B
047A
04DF
0563
052A
0345
FFFE
FCD4
FB09
FA8E
FA97
FABF
FB1F
FB85
FB61
FAAA
FA3B
FABE
FBAF
FBF5
FB4F
FAA2
FABD
FB66
FBC9
FB88
FB02
FAB5
FAC0
FB02
FB5D
FB9D
FB81
FB16
FADD
FB3A
FBDA
FBFD
FB6C
FAC7
FAC6
FB5C
FBD9
FBC1
FB51
FB0D
FB26
FB6A
FBAE
FBF0
FC0F
FBB7
FAEF
FA80
FB6C
FDE2
00FD
039F
0547
060C
060B
055E
0483
0442
04D3
0572
0541
047A
042C
04BF
055D
052C
047C
044A
04D7
0569
055E
04E7
049D
04BB
0506
053C
0544
0505
0488
042D
0460
04ED
051E
04B6
044B
0460
04A8
049F
0471
049F
0505
04EF
0441
03D8
0473
0593
05F0
04F3
0324
011F
FED3
FC2D
F9FA
F948
FA12
FB24
FB6A
FAFD
FAB4
FB01
FB7C
FB87
FB21
FAEB
FB4C
FBD7
FBC5
FAFB
FA49
FA77
FB57
FBF5
FBAA
FAC2
FA24
FA62
FB3B
FBED
FBE4
FB32
FA81
FA88
FB50
FC09
FBFB
FB6E
FB42
FB97
FBA4
FB17
FAC7
FB71
FC5F
FC34
FAEB
FA10
FACA
FC75
FDD3
FEFD
011A
042F
067C
068F
052E
044F
04AD
0555
0559
0502
050C
056E
0576
04D8
0426
0423
04DA
058F
0580
04A1
03AD
0392
0493
05DC
0627
051B
03CE
03A7
04C2
05D4
05B5
04BD
0432
04A7
0554
0534
046B
040E
0493
051C
04AE
03B2
0382
048A
05AD
05B6
04CA
03C2
029C
0080
FD4B
FA58
F939
F9F3
FB26
FBAC
FB8C
FB49
FB08
FAC2
FAB8
FB15
FB7E
FB7C
FB27
FAEE
FAEC
FAE8
FAEB
FB3F
FBBE
FBBA
FAF6
FA55
FADE
FC2A
FC9F
FB8D
FA40
FA5F
FBB2
FC6B
FB9A
FA65
FA6A
FB94
FC4F
FBB3
FAA8
FA91
FB76
FC1A
FBB8
FAED
FAAC
FB00
FB5D
FBE3
FD73
005F
0398
0597
05E2
053B
0497
0457
0482
0512
05CA
0606
0565
0472
042A
04C1
055D
0540
04BD
0496
04DF
0509
04DC
04C0
04F3
050D
04B2
0448
047A
0517
0537
048D
0403
047A
0572
059C
04B2
03E6
044F
0568
05C1
04E6
03EB
03F6
04D5
0572
053A
049B
0437
0430
0451
0487
04D8
050E
04BD
0395
0190
FEE8
FC27
FA35
F9C7
FA96
FB73
FB79
FAED
FAA6
FAE6
FB2C
FB15
FAD8
FAD4
FB00
FB16
FB18
FB39
FB5B
FB23
FAA5
FA88
FB1B
FBB7
FB7C
FA8C
F9FE
FA8D
FBB1
FC3F
FBB4
FAB1
FA3F
FAC1
FBA8
FC1A
FBBE
FAF5
FA6F
FA98
FB4F
FBFE
FC0E
FB72
FAC4
FAAE
FB36
FBB7
FBA8
FB3E
FB0A
FB1E
FB00
FAC1
FB89
FE59
0252
0526
0598
04C8
048D
0532
0595
051A
0484
04A8
053A
0562
0512
04F5
052E
051C
0484
0439
04E8
05E3
05E2
04C3
03BF
03E2
04E3
05A9
0589
04C5
0419
0409
048E
0533
0568
04F3
043D
0403
0490
055B
0590
0506
045E
0441
04AA
050C
050B
04D9
04CE
04D6
0489
03EA
03B7
048D
05CB
05D7
03C8
006B
FD65
FBA8
FAF7
FAB9
FAAC
FAD1
FB0E
FB32
FB2F
FB1B
FAFE
FAD4
FABE
FAE8
FB3D
FB67
FB4A
FB1E
FB06
FAE7
FACE
FB08
FB8F
FBC1
FB2E
FA64
FA6B
FB5C
FC1C
FBB8
FAAA
FA41
FAF4
FBD3
FBD7
FB2A
FAC4
FB0E
FB7C
FB84
FB59
FB76
FBCD
FBCE
FB37
FA8B
FA8C
FB48
FBFC
FBF2
FB4A
FAB6
FAAA
FB37
FC86
FEDA
01DF
0475
05A1
058D
0530
051F
051A
04D7
04AD
0506
0584
0564
04AB
043C
048D
04F7
04C4
0455
0483
053A
0580
04E3
042E
0448
04F3
052F
04B3
0449
049A
053D
055B
04E7
0494
04BE
04FA
04D2
0478
0471
04CD
050D
04D8
0470
0459
04A8
04F3
04E3
049B
0470
0478
0485
0488
04B0
0504
0501
03D9
013F
FDE6
FB20
F9E0
FA1A
FAEE
FB7A
FB6E
FB0B
FAB9
FAB1
FAF0
FB47
FB67
FB1F
FA9D
FA63
FAC0
FB69
FBB3
FB57
FAC9
FAB4
FB26
FB8F
FB7C
FB1D
FAE5
FAF2
FB05
FAF7
FAE9
FAFF
FB25
FB31
FB1B
FB0C
FB23
FB53
FB6E
FB5C
FB37
FB25
FB24
FB1D
FB11
FB1C
FB44
FB5D
FB44
FB1D
FB30
FB67
FB5A
FB20
FBCE
FE6E
025D
0571
0627
052D
045C
0490
0522
054E
0538
054E
055C
04F3
0465
0485
0550
05B1
0509
0430
0453
054A
05D2
0557
04A3
04AE
054D
0596
0528
0490
0471
04BB
04F3
04EA
04D2
04D1
04D4
04D3
04E1
04F5
04E6
04AA
0479
0490
04DD
0511
04F4
04AC
0491
04BB
04DD
04B5
0481
04C5
0576
0594
03F2
0089
FCCC
FA7D
FA1F
FABD
FB20
FAFB
FAC8
FADB
FB02
FAF3
FAC8
FAC4
FADD
FAD8
FAB8
FAC9
FB1D
FB45
FAE1
FA44
FA32
FAE7
FBAC
FBA2
FAD7
FA41
FA98
FB77
FBE0
FB70
FAC7
FAB7
FB4C
FBD5
FBC1
FB42
FAFD
FB32
FB7B
FB66
FB1D
FB23
FB84
FBBB
FB6D
FAEF
FAD8
FB36
FB90
FB8F
FB51
FB12
FAE5
FB24
FCA7
FFCD
0370
0598
059B
04D5
04DC
0596
05D0
052F
04A9
04F7
0586
056B
04CF
0498
04F3
0513
049D
045A
04F6
05C3
059D
049E
0411
04A6
0583
0576
0489
03DE
0430
04FD
0549
04E3
0478
048C
04DE
04E7
04A6
048E
04D7
0524
04FE
047F
043E
048B
04F5
04DD
0459
040D
043E
048C
04B6
0500
0573
0529
031D
FF9C
FC59
FAC4
FAAD
FAD3
FA8C
FA47
FA84
FAFC
FB17
FAD9
FAC0
FAFE
FB40
FB43
FB2C
FB30
FB40
FB27
FAE7
FAC2
FAE5
FB2F
FB56
FB3B
FB0A
FB06
FB44
FB8F
FB9F
FB5A
FAFF
FAE1
FB0D
FB43
FB4D
FB3C
FB35
FB38
FB37
FB47
FB8B
FBDB
FBD4
FB59
FADD
FAF1
FB86
FBF9
FBDA
FB68
FB1B
FAFB
FADD
FB2D
FCD9
0020
03B9
05CE
05D8
0510
04DD
0553
0593
0544
04F1
050F
0541
04FE
0483
0485
0515
0571
051C
049E
04B6
053E
0564
04DB
044E
046C
04FC
053D
04EB
0484
048C
04E5
0513
04EE
04B8
04A6
04A5
049E
04AD
04E1
04FE
04BF
0449
0422
048B
0514
051D
04AA
0467
04B7
0510
04BA
03FB
03E6
04BB
0510
0333
FF47
FB77
F9D3
FA52
FB47
FB71
FB04
FAC4
FAD6
FADC
FAC5
FADC
FB28
FB48
FB07
FABD
FAD5
FB34
FB59
FB0D
FAAA
FAA0
FAED
FB35
FB3D
FB16
FAF7
FB05
FB3A
FB65
FB4F
FB07
FAE5
FB22
FB80
FB92
FB46
FB04
FB28
FB7D
FB87
FB31
FAEC
FB18
FB8C
FBD1
FBAC
FB47
FB00
FB2A
FBB9
FC1D
FBB8
FAC9
FAB9
FCDC
00D3
047E
05FD
0588
04DC
0512
05A5
05AF
0548
0520
0551
0554
0502
04DA
0522
055F
050E
047F
047A
0515
0584
0532
048A
0459
04B2
04FF
04E6
04A8
04A5
04DB
050D
0513
04FE
04F9
050F
051C
04F1
0498
0461
048A
04EE
051B
04D6
0468
0444
0474
049F
049B
0491
048D
046D
045E
04CF
0584
052D
02AC
FEA0
FB28
F9DB
FA5D
FB1F
FB2F
FAD3
FAA4
FAB7
FAD9
FB07
FB3D
FB40
FAF8
FAC1
FAF4
FB51
FB54
FAFC
FACA
FAFD
FB3F
FB2E
FAF4
FAFC
FB43
FB5D
FB25
FAF7
FB1C
FB59
FB55
FB1F
FB00
FB05
FB14
FB32
FB66
FB81
FB56
FB1C
FB32
FB8E
FBA8
FB41
FAD2
FAEB
FB56
FB6E
FB32
FB49
FBC1
FBB8
FADF
FA9F
FCBE
00F6
04CD
0628
0574
04B6
0502
059B
0586
04FE
04D7
0529
0556
0517
04D5
04E4
0510
0506
04DB
04D6
0501
051D
0506
04DF
04D0
04D1
04C7
04B9
04B8
04BA
04AC
0499
0496
049E
04AC
04C4
04DD
04D8
04C1
04C6
04E8
04E4
049C
045D
0482
04D8
04D3
0460
041F
0479
04E1
0497
03FD
0437
053C
0535
0293
FE3D
FAD5
F9E5
FA85
FAF3
FAA6
FA5E
FA97
FAE3
FACE
FAA0
FAC8
FB1D
FB32
FB10
FB12
FB3D
FB3D
FB00
FADE
FB0F
FB59
FB6C
FB4A
FB32
FB34
FB2B
FB0F
FB0B
FB2B
FB40
FB2E
FB24
FB42
FB60
FB51
FB38
FB41
FB55
FB4A
FB36
FB42
FB57
FB42
FB19
FB32
FB92
FBC0
FB77
FB2C
FB6C
FBDD
FB9D
FAD7
FB26
FDD1
01EE
051B
05F4
0544
04B4
04E8
0548
053A
04F1
04E4
0516
0529
0502
04D7
04D1
04DF
04EB
04F5
0501
0506
0502
04F5
04DF
04CD
04D1
04EC
04F6
04D6
04A4
0498
04BA
04D5
04C4
04AF
04CE
0500
04F6
04AF
0489
04AE
04D6
04C7
04B7
04E0
0508
04D2
0470
0472
04DC
04F1
044E
03C0
0449
055D
0504
021A
FDF2
FB03
FA59
FADC
FB1B
FAE2
FAE1
FB4C
FB8E
FB40
FAC6
FAB7
FB0E
FB53
FB4F
FB38
FB39
FB33
FB07
FAE0
FAF5
FB3B
FB70
FB6F
FB57
FB52
FB5B
FB51
FB2E
FB13
FB15
FB21
FB18
FB00
FAF8
FB03
FB0C
FB09
FB16
FB49
FB81
FB87
FB68
FB74
FBB5
FBAD
FB08
FA86
FB9F
FEE5
02EF
057E
05AC
04AF
044B
04E3
0579
0549
04BB
0494
04E3
051D
0509
04F5
0515
0527
04E8
048D
0479
04AA
04C4
04A0
0484
04AA
04E2
04E0
04AE
0493
049A
0490
0469
045C
0488
04B3
049D
046B
0473
04B6
04D8
04B6
04A3
04E6
052D
04F5
046B
045B
04FF
0533
0377
FFC3
FBF3
FA09
FA3F
FB18
FB35
FAAC
FA68
FAC4
FB36
FB34
FAF0
FAE9
FB28
FB4C
FB2D
FB10
FB2E
FB58
FB3F
FAF7
FAE0
FB1A
FB5F
FB63
FB39
FB1D
FB1F
FB22
FB20
FB2E
FB46
FB41
FB19
FB0B
FB3E
FB8B
FBA8
FB97
FB91
FBA1
FB8A
FB3E
FB1D
FB6B
FBBE
FB66
FA9B
FAC3
FD1D
011E
04A9
060B
058A
04C4
04CE
054E
056D
050E
04C5
04E9
0523
050E
04CD
04C1
04EC
04F5
04BC
048C
04AD
04F6
0508
04D4
04A0
049C
04AD
04AB
04A2
04A7
04A8
048F
047D
049F
04DA
04E6
04B3
048F
04AB
04CD
04A5
045B
045D
04A5
04AA
043E
040E
04BA
058C
04CE
01AD
FD7B
FA91
FA06
FADE
FB77
FB4C
FAFC
FB0C
FB39
FB13
FABF
FAB2
FAFE
FB38
FB19
FADC
FADB
FB0F
FB21
FAF6
FAD0
FAE8
FB1D
FB2D
FB16
FB0C
FB27
FB43
FB45
FB40
FB4E
FB56
FB3B
FB13
FB16
FB46
FB69
FB60
FB5A
FB82
FBA7
FB7C
FB28
FB27
FB7F
FB8A
FAE8
FA7C
FBD7
FF60
0375
05DB
05F0
0507
04B0
0515
055C
0517
04C1
04DB
052D
0535
04F4
04DF
0526
0566
0543
04EE
04D3
0500
0521
050B
04F2
0509
0533
052F
04F6
04BD
04A8
04A9
04B5
04D4
04F9
04F3
04B1
046D
0465
047E
0472
0447
0456
04B9
04F9
04A9
042E
045F
0537
0557
0353
FF73
FBBD
FA06
FA46
FB06
FB25
FACD
FAAE
FAE8
FB09
FAD6
FA97
FA96
FAB3
FAB2
FAA9
FAD9
FB3E
FB7F
FB64
FB1F
FAFD
FB05
FB10
FB12
FB21
FB37
FB37
FB21
FB1F
FB3D
FB4B
FB23
FAFB
FB24
FB8A
FBB9
FB7C
FB35
FB51
FBA2
FB9C
FB32
FB02
FB69
FBD6
FB79
FAA9
FAFD
FD9A
01AB
04EE
05EF
0542
048D
04A8
051B
0530
04F0
04DA
050E
0539
052B
0523
0552
057E
0553
04ED
04BA
04E0
050D
04FA
04C9
04B9
04BD
049F
046B
0468
04A5
04D1
04B5
048E
04AC
04F0
04EE
049B
046F
04A6
04DD
04A8
0444
0444
04A8
04CA
046A
0439
04DA
0592
04A7
0165
FD3B
FA77
F9FD
FABF
FB3B
FB0D
FACB
FADC
FB02
FAEA
FAB5
FAB2
FAD8
FADE
FAB8
FAAF
FAF0
FB42
FB55
FB2A
FB08
FB13
FB2B
FB2B
FB20
FB28
FB3B
FB3E
FB38
FB49
FB72
FB86
FB72
FB61
FB7A
FB9A
FB80
FB3A
FB23
FB5C
FB8A
FB5A
FB11
FB34
FBA7
FB9D
FACD
FA63
FC08
FFE8
040B
0630
05F3
04E3
048C
04FC
0550
0524
04EF
0517
0555
0537
04DB
04BC
04FB
0539
0522
04DB
04B4
04C0
04D4
04DE
04F2
0513
0528
0526
0523
0523
0500
04B4
0483
04AA
04F6
04F1
0485
042D
0453
04BA
04D4
048B
0463
04AB
04FF
04E0
0493
04D2
0583
054D
02EC
FEE7
FB63
FA17
FAB4
FB7F
FB52
FA90
FA3E
FAA8
FB31
FB45
FAF6
FAB6
FAB4
FACE
FADF
FAE8
FAF3
FB00
FB12
FB2D
FB3E
FB28
FAF2
FAD9
FB01
FB38
FB32
FAF5
FADA
FB0E
FB4C
FB41
FB06
FB01
FB4E
FB9A
FB98
FB69
FB52
FB45
FB09
FAC2
FAE9
FB8A
FBE5
FB53
FA7B
FB08
FDF1
0221
054B
0615
052D
0446
0450
04F0
055D
0559
0528
0503
04EB
04DF
04F4
051F
052C
0507
04E9
0507
0541
054B
0515
04E8
04F5
0513
04FC
04BF
04A6
04CA
04ED
04DA
04AA
048E
0480
0465
0455
047C
04BE
04C1
0474
0447
049B
051E
052A
04BE
04A4
053F
0593
040D
006D
FC66
FA1D
FA20
FB2B
FBBE
FB89
FB2A
FB13
FB17
FAF0
FABE
FAC3
FAF7
FB14
FB05
FAFB
FB14
FB2C
FB15
FAE6
FADB
FAFD
FB1C
FB16
FB07
FB17
FB3E
FB5A
FB67
FB79
FB8B
FB82
FB60
FB4F
FB5D
FB5A
FB1F
FAE6
FB0B
FB7F
FBB7
FB68
FB02
FB24
FBA1
FB9F
FAEC
FABD
FC95
0068
0447
0635
05FD
050C
04AE
04E9
0512
04EF
04D7
0502
0531
0524
04FE
0503
052C
0536
050F
04EB
04E9
04E6
04C0
049A
04AA
04E3
04FF
04E0
04B2
04A2
04A5
049C
048F
04A0
04C4
04CD
04B5
04B1
04DF
0506
04E4
0499
0487
04C2
04E1
04A1
0467
04C2
055B
04DC
0246
FE4C
FAF7
F9C2
FA58
FB33
FB51
FAEB
FAAD
FABD
FAC6
FAAB
FAB0
FAFC
FB48
FB44
FB0C
FB00
FB30
FB4D
FB23
FAE5
FADF
FB05
FB15
FB03
FB07
FB44
FB8E
FBA8
FB90
FB68
FB3F
FB0C
FAE5
FAEE
FB1A
FB29
FB07
FAF7
FB2B
FB6F
FB6C
FB3B
FB4E
FBAC
FBB3
FAFF
FA66
FB78
FEC1
02D7
058D
0602
0539
04B4
04EA
0546
0544
050F
0505
051B
0504
04C0
04A2
04D8
0520
052B
0500
04E4
04F8
0516
0519
050C
0505
04FB
04DD
04B9
04AD
04B8
04B5
049C
0491
04B2
04E5
0501
0504
050C
0510
04EB
04A7
0494
04D8
051D
04F1
0486
0494
0548
0587
03D5
001B
FC22
FA01
FA20
FB1B
FB7B
FB20
FADC
FB15
FB55
FB21
FAB6
FA9C
FAE0
FB0D
FAEB
FAC5
FAED
FB3B
FB4B
FB16
FAF6
FB1B
FB4A
FB43
FB22
FB29
FB4F
FB4F
FB15
FAE1
FAEF
FB23
FB41
FB3E
FB3E
FB44
FB38
FB24
FB33
FB56
FB3C
FADA
FAA9
FB0B
FB8F
FB5A
FA7F
FA79
FCBB
00D6
048E
0602
0572
049F
04B5
0557
0596
0546
04FD
0517
0545
0524
04D3
04B5
04D8
04EF
04D2
04B7
04D8
0513
051B
04E0
04A3
049C
04BA
04CB
04C1
04B4
04B9
04CA
04D7
04D3
04B8
048E
047B
04A9
0503
0532
0502
04AB
0496
04CB
04E2
04A7
048B
050B
05AC
04FD
0210
FDDC
FA9F
F9C4
FAA0
FB6B
FB39
FA9C
FA7C
FADD
FB19
FAEC
FAC5
FAFB
FB45
FB31
FAD6
FAB2
FAF3
FB3C
FB3C
FB19
FB28
FB5C
FB63
FB27
FAF9
FB1B
FB63
FB84
FB6E
FB50
FB3F
FB31
FB26
FB32
FB44
FB25
FADC
FAC4
FB18
FB83
FB7F
FB19
FAF0
FB44
FB7B
FB0C
FAAA
FBDC
FF34
034B
05FA
066F
05B2
052C
052E
0526
04D2
049D
04DC
053B
0532
04C4
0472
048A
04CC
04DD
04C1
04C2
04F8
0529
051F
04E7
04B9
04B8
04DD
0508
0514
04F1
04BC
04AF
04DD
050B
04EA
0486
044D
0489
04FB
0524
04EF
04C5
04EA
050F
04C3
043D
0435
04C8
04D9
030D
FF72
FBCF
FA09
FA56
FB4E
FB9A
FB38
FAF8
FB33
FB74
FB44
FADD
FAC4
FB11
FB5C
FB5E
FB42
FB49
FB62
FB51
FB14
FAE0
FAD2
FAD2
FACC
FAD3
FAF8
FB22
FB34
FB3A
FB49
FB4A
FB1C
FAE4
FAF2
FB44
FB6B
FB30
FAFB
FB3E
FBA4
FB67
FA9D
FABB
FD25
0156
0503
0658
05AA
04BB
04A4
0509
051E
04D4
04AC
04D5
04FB
04E2
04BE
04C9
04DC
04B6
0472
0462
0496
04C6
04BE
04A1
04A4
04C5
04E0
04F1
0503
0504
04D6
049D
04A3
04E4
04F9
04AC
0463
04A2
053A
0561
04CA
0439
0486
053A
04B8
0202
FE15
FB17
FA3B
FACB
FB49
FB0F
FA9B
FA91
FAE6
FB26
FB22
FB15
FB29
FB39
FB1C
FAF4
FAFA
FB2C
FB4C
FB3E
FB2A
FB38
FB54
FB4D
FB1F
FAF8
FAF8
FB13
FB32
FB53
FB69
FB55
FB12
FAE1
FAFD
FB42
FB57
FB44
FB76
FBFA
FC21
FB57
FA62
FB13
FE4B
029C
056E
05A2
0484
0411
04C0
0581
0577
0500
04E5
0533
0557
0519
04D8
04DE
04F0
04C9
049C
04BC
0505
0511
04D9
04C1
04F7
051E
04E4
0489
0489
04E2
0519
04F4
04C9
04E4
0508
04E4
04AE
04D4
052B
0514
047D
043C
04D9
0559
03F9
0055
FC44
FA13
FA37
FB25
FB57
FACE
FA7F
FAD6
FB4F
FB56
FB07
FAD3
FADA
FADF
FAC4
FAAB
FAAC
FAB2
FAB8
FADF
FB32
FB74
FB64
FB1C
FAFC
FB2D
FB6A
FB67
FB38
FB27
FB49
FB61
FB4F
FB36
FB39
FB3C
FB1C
FB0D
FB55
FBB6
FB8B
FACA
FA9A
FC65
0020
03E7
05B9
0568
048C
0492
0552
05BB
0562
04E6
04E8
053B
054D
050A
04DF
0502
052B
0516
04E9
04E3
04F1
04DB
04BA
04D8
0530
0555
050B
04A4
048E
04BC
04CB
04A6
049C
04C5
04CD
0487
044F
047E
04BD
047F
0402
0435
0536
0582
0366
FF38
FB6A
FA0E
FACC
FBB0
FB88
FAD5
FA8A
FAB5
FAC2
FA8C
FA7E
FAC9
FB0E
FAFB
FAC9
FAD3
FB03
FB0B
FAF5
FB14
FB61
FB6C
FB02
FA92
FA9C
FAFE
FB28
FAF8
FADF
FB25
FB71
FB54
FB03
FB04
FB5A
FB7C
FB3E
FB2F
FBB3
FC2E
FBB3
FA9A
FAB0
FD4C
018D
04F7
05F1
0524
0458
0473
04EE
050A
04D3
04CB
050E
053E
0527
050C
052E
0561
055D
052F
051E
052F
051D
04D6
04B3
04F7
055B
055F
04FC
04AB
04BA
04E2
04C5
0489
049C
04FF
0533
04F9
04AA
049F
049D
0452
0414
0480
0536
04A6
01BA
FD87
FA88
FA11
FB13
FBA5
FB3F
FACF
FB03
FB5C
FB26
FA9E
FA90
FB13
FB6B
FB23
FAB2
FAB3
FB01
FB0D
FACE
FABD
FB02
FB2E
FAED
FA96
FAAB
FB0F
FB32
FAEE
FABE
FAEF
FB2D
FB13
FAD5
FAE3
FB27
FB32
FB06
FB2F
FBC9
FC0B
FB5A
FA9F
FBAC
FF15
0328
0587
0592
04B1
0472
04FC
057B
057F
0557
0556
0550
0509
04B5
04B5
04FC
0526
050A
04E6
04F2
0507
04EB
04B5
04B0
04E9
0522
052B
051F
051E
0514
04E3
04B3
04C7
050C
0520
04DE
04A1
04C0
04FF
04E1
0482
049C
0568
05C4
0423
0063
FC5A
FA24
FA1D
FAD9
FAF7
FA7A
FA3A
FA86
FAE0
FAE0
FAC1
FAD8
FB02
FADF
FA86
FA6E
FABA
FB00
FAEB
FABC
FADF
FB3A
FB5B
FB21
FAED
FAFD
FB15
FAF1
FACB
FB01
FB6C
FB7F
FB24
FAEE
FB3A
FB96
FB78
FB22
FB43
FBBF
FBA4
FABF
FA85
FCA7
00CA
047D
05C4
0514
045A
049A
0532
054F
051E
053B
0594
0594
0526
04E4
0523
056F
0549
04F1
04F6
0545
053F
04BB
0454
048A
0502
050D
04AB
0475
04AD
04DD
04A3
0457
0471
04B8
0497
0421
0417
04BC
053E
04CF
03F9
040B
0522
057D
0360
FF47
FB9B
FA30
FA96
FB22
FB02
FAC3
FB06
FB80
FB81
FB00
FA9B
FAAC
FAE4
FAE1
FAC3
FADE
FB2A
FB4B
FB2A
FB14
FB3A
FB62
FB46
FB09
FB03
FB30
FB39
FB06
FAF9
FB4F
FBA9
FB80
FAF5
FAB6
FB11
FB8E
FBAE
FB9E
FBC0
FBCC
FB2A
FA49
FAD2
FDE2
024E
0576
05F0
04E1
0458
04F0
059C
0579
04E9
04BC
04F2
04EE
0488
0446
0480
04D9
04E5
04C8
04D4
04E2
0493
0417
0414
04BA
0563
0568
0501
04DD
0516
051B
04AF
045A
048F
04EC
04D7
0483
04A5
053E
0564
04A3
03E9
0451
053A
0488
012E
FCC9
FA18
FA12
FB37
FB9E
FB04
FA71
FA8B
FAEE
FB0C
FAFF
FB22
FB5B
FB46
FAEC
FACD
FB2C
FBB0
FBDC
FBA5
FB61
FB3E
FB2A
FB1C
FB37
FB7A
FBA2
FB7C
FB38
FB23
FB32
FB17
FAD2
FAC9
FB2B
FB8C
FB74
FB23
FB4D
FBF6
FC30
FB5D
FA82
FB90
FF26
037F
0613
061E
0516
04B1
051D
0563
050B
04AA
04DA
0557
0575
0521
04E2
0504
0531
0507
04A5
0473
0487
04AB
04C0
04D6
04E3
04BD
0474
045E
049D
04CE
048B
041E
0431
04D1
0543
0502
048C
049C
0505
04EB
042D
03C9
045E
04D8
0360
FFC6
FC11
FA60
FAA3
FB1C
FAB7
FA1A
FA52
FB38
FBBD
FB62
FABB
FA7B
FA90
FA84
FA51
FA59
FAC0
FB3B
FB82
FB97
FB8D
FB54
FAF5
FAC4
FB06
FB83
FBBF
FB99
FB69
FB6B
FB63
FB15
FACD
FAFA
FB71
FB8C
FB22
FAE5
FB5E
FBF8
FBA7
FA9A
FA92
FD0A
0148
04D5
05FB
0551
04B2
050B
05B8
05C6
0537
04D2
0501
056E
059B
0573
052A
04DE
0499
0481
04BB
0522
0554
0528
04DF
04C8
04D9
04D5
04AD
048B
047D
0465
0444
045A
04B8
04FB
04C8
046F
04A7
0575
05E2
0534
041D
03FB
04DA
04E6
0273
FE39
FADE
FA1F
FB1B
FBBB
FB2D
FA64
FA5F
FADE
FB08
FABF
FAA0
FAEF
FB2F
FAFB
FAA8
FAC3
FB3C
FB85
FB6B
FB4B
FB6C
FB97
FB7E
FB3C
FB25
FB3E
FB47
FB3A
FB5A
FBA3
FBA0
FB0E
FA6A
FA61
FAE8
FB4F
FB48
FB46
FBA7
FBE9
FB6B
FABF
FB8C
FEA8
02C1
0582
05EA
0511
0495
04DA
051F
04E4
0494
04C2
0553
05B2
0598
0541
04F2
04B1
047E
047E
04BE
04F9
04E9
04A9
049C
04E1
0520
0502
04AC
0485
04AE
04EB
0503
04FF
04F6
04D8
04A2
0492
04D4
0519
04DF
0441
040D
04AA
051E
03C8
004D
FC66
FA4A
FA77
FB6F
FB9C
FAF8
FA8B
FAD0
FB2C
FB01
FA90
FA83
FAEC
FB3F
FB2E
FB06
FB21
FB4F
FB35
FAF1
FAF2
FB4F
FB99
FB7B
FB29
FB0C
FB27
FB33
FB21
FB2A
FB52
FB4D
FB01
FAD5
FB20
FB8F
FB92
FB41
FB4D
FBE8
FC3C
FB99
FAD6
FBD2
FF33
034F
05C0
05D8
04FE
04C5
0545
05A0
0572
0532
053E
0547
04EF
0476
0461
04AA
04D1
04A0
047C
04C0
0529
0536
04DD
048C
0485
0493
0482
047B
04A8
04C2
0472
03F3
03F7
04A5
0545
0531
04CD
0500
05A8
0546
02A7
FE9B
FB65
FA6E
FAF7
FB52
FAE0
FA6C
FAB8
FB6B
FBB0
FB63
FB11
FB10
FB16
FADA
FAA9
FAEA
FB72
FBA8
FB64
FB25
FB4D
FB90
FB74
FB18
FB0B
FB70
FBC0
FB99
FB59
FB87
FBEE
FBDE
FB47
FAF7
FB69
FBEA
FB7E
FA95
FAFF
FDD4
01E8
04D6
057D
04E3
04A2
051B
0589
056A
0517
0508
0518
04EC
04A2
04A5
04F5
0514
04C8
047E
04AD
0518
0524
04B3
044D
0458
0493
0493
0471
0496
04F8
050B
0496
0427
0451
04CB
04CC
044B
0434
0509
05AE
045A
00BA
FCAD
FA7C
FA8F
FB61
FB71
FACE
FA70
FABA
FB13
FAF0
FA92
FA8E
FAF0
FB3F
FB3C
FB2B
FB4F
FB7F
FB6D
FB30
FB24
FB5D
FB88
FB69
FB31
FB22
FB2C
FB1F
FB1A
FB6B
FBEE
FC0A
FB82
FAFA
FB30
FBDD
FBEA
FB0D
FAAA
FC7B
0069
0449
0600
058D
04A1
048B
050B
053B
04EF
04BF
04FD
0546
0532
04F3
04F8
053A
0546
04F1
0492
0484
04A1
0492
0458
044E
0493
04DA
04DA
04B8
04BC
04E0
04DE
04B0
049D
04BB
04B6
045D
0428
04A8
056C
04FD
025D
FE6C
FB55
FA72
FB1A
FB9B
FB2D
FA75
FA5D
FAE5
FB58
FB56
FB2A
FB32
FB59
FB61
FB52
FB6A
FBA4
FBB8
FB8C
FB5F
FB72
FBA4
FBB2
FB9C
FB97
FBA1
FB7D
FB21
FAEE
FB30
FB95
FB91
FB2E
FB0F
FB7C
FBD3
FB5F
FAA9
FB4B
FE26
021D
0501
05C1
0539
04EB
0544
058E
0532
0483
0430
045F
04AA
04C8
04D7
04FC
0519
0506
04D5
04B4
0498
0459
040B
0402
0457
04AC
049F
0450
0437
0475
04AE
049A
0471
0488
04B7
048F
042D
044B
0522
0595
0412
0070
FC83
FA6D
FA8F
FB6E
FB93
FB06
FAC3
FB35
FBBE
FBB6
FB46
FB0B
FB31
FB4B
FB0D
FABB
FABC
FB0C
FB4E
FB52
FB45
FB5B
FB8E
FBBF
FBE0
FBE7
FBBB
FB60
FB26
FB5D
FBD7
FC05
FBB2
FB5A
FB81
FBDE
FBA6
FAD7
FABB
FCAF
0068
03EE
0582
0537
0489
0491
051D
056C
054D
0527
0537
053C
04FC
04AA
049E
04D0
04F2
04E9
04E7
0504
050D
04D0
0473
0441
0444
044A
0452
0492
0508
054A
0506
0489
0465
049B
0492
0403
039C
041F
050E
04B7
020C
FE10
FB08
FA45
FB0D
FBBD
FB97
FB1D
FAF6
FB1E
FB32
FB1F
FB1E
FB32
FB25
FAF5
FAF4
FB40
FB76
FB2E
FA9C
FA69
FAD2
FB5C
FB7F
FB53
FB4A
FB74
FB74
FB30
FB12
FB66
FBC8
FBB3
FB5A
FB7B
FC22
FC54
FB6C
FA7B
FB86
FF27
0382
0605
05FD
04F7
04A9
052D
057A
0514
0493
0499
04F2
0503
04BD
0499
04D8
0526
0520
04D7
049C
0487
047A
047E
04B4
04F5
04E1
0475
0446
04C6
0588
05A7
04F2
043C
0443
04AD
049D
0419
041A
04F6
0555
0375
FF75
FB98
F9FF
FA86
FB50
FB1F
FA79
FA77
FB2B
FBB2
FB82
FB03
FACA
FAD5
FAD1
FAC6
FB06
FB82
FBB9
FB62
FAE0
FABF
FB08
FB59
FB77
FB8A
FBA7
FB98
FB44
FAFD
FB1F
FB76
FB75
FB12
FAF0
FB6F
FBEF
FB8A
FA98
FAC8
FD62
018D
04EE
05F6
054D
04B8
0510
05B2
05BD
053F
04E0
04DF
04E2
04B2
049D
04EE
055C
055E
04F2
049E
04BA
04FF
0507
04E3
04E8
0514
050B
04A8
044C
0455
0499
04B0
0496
04A0
04D5
04C6
044E
040E
04A0
0560
04B1
01C5
FDD6
FB18
FA84
FB12
FB36
FAA3
FA3F
FAA4
FB4C
FB5F
FACF
FA52
FA68
FAD8
FB2C
FB47
FB51
FB4F
FB27
FAF1
FAFA
FB52
FBA3
FBA3
FB80
FB8E
FBB4
FB88
FB04
FAB9
FB13
FBAF
FBD6
FB85
FB76
FBF6
FC46
FBAB
FAE4
FBC8
FF1F
0351
05D3
05BD
047C
03FF
04AB
057B
05A2
0567
056B
05AE
05B3
0556
04FA
04ED
04FF
04E1
0498
0465
045D
0461
046A
0498
04E4
0506
04D0
0486
0487
04C6
04D6
048F
0456
0482
04C9
04A0
0423
041D
04D2
0523
0383
FFDA
FC0C
FA30
FA7C
FB51
FB41
FA85
FA3B
FABB
FB3D
FB0F
FA84
FA5E
FAB6
FAF4
FACD
FAA8
FAF6
FB79
FBA2
FB61
FB32
FB64
FBAF
FBAD
FB63
FB1F
FAFE
FAEE
FB00
FB55
FBB0
FB91
FAFC
FAB1
FB38
FBEF
FBC0
FAD7
FAFA
FD9F
01E7
0538
05F3
04FD
045E
04D8
057F
0564
04DC
04CF
055F
05D2
05AE
0542
0507
04EE
04B3
0475
048F
04F0
0514
04CA
0487
04B9
0518
0511
04B1
049B
050D
0568
0518
0483
0481
050E
053A
048F
03F1
045E
0531
047C
0160
FD63
FAE5
FA98
FB1F
FB13
FA90
FA82
FB0D
FB69
FB21
FAB7
FAC6
FB1B
FB1C
FAC8
FAA4
FAE1
FB0F
FAE8
FAD3
FB41
FBDC
FBDD
FB2F
FAA5
FADA
FB59
FB49
FAB6
FA84
FB1D
FBCF
FBC3
FB37
FB1A
FB9B
FBD0
FB26
FAA5
FC11
FFB5
03AC
05B6
0574
0477
0441
04D3
053D
051A
04EC
0523
0574
0557
04DF
0490
04A2
04C7
04BD
04B4
04E1
0518
0510
04EB
050D
0566
0564
04C1
040B
0402
0496
04FE
04D8
049C
04C9
050C
04D0
0452
0473
0540
0552
0331
FF3E
FBA0
FA1E
FA7F
FB33
FB37
FADB
FAD7
FB37
FB7C
FB64
FB2C
FB20
FB37
FB41
FB37
FB2E
FB28
FB14
FAFC
FAFF
FB1C
FB28
FB1A
FB24
FB64
FBA3
FB91
FB44
FB29
FB6F
FBAF
FB77
FB03
FB00
FB86
FBC1
FB06
FA22
FAE4
FE20
0270
0565
05E3
04F7
045F
04AD
052B
0529
04D8
04C4
04F8
050C
04DB
04B3
04D7
051A
0521
04D7
047F
045B
0479
04B5
04E1
04D5
048D
044C
0466
04D4
051A
04CE
0435
0412
04B5
0581
0598
04EE
0468
04A9
050A
040E
0110
FD3D
FA97
FA18
FAED
FB94
FB6B
FAFB
FAF3
FB41
FB5F
FB20
FAE1
FAF1
FB27
FB33
FB1A
FB20
FB53
FB75
FB60
FB3D
FB4C
FB89
FBB4
FBA1
FB5F
FB1D
FAFF
FB13
FB42
FB4B
FB04
FAB3
FADD
FB92
FC18
FBAD
FAB6
FAB5
FCD6
008B
03E5
0565
0537
04A3
0493
04E9
0518
04EE
04AB
048F
049C
04BE
04EF
0527
0541
0520
04E0
04C4
04DD
04F3
04CF
048A
0471
049C
04CB
04B9
0477
0455
0477
04AE
04C4
04C3
04C1
049E
0445
040F
047F
0551
0536
02FE
FF21
FBA7
FA48
FAD0
FBA2
FB9F
FB1D
FAF9
FB48
FB6A
FB1D
FADA
FB0E
FB75
FB7E
FB28
FAF7
FB2B
FB5D
FB1C
FAA3
FA94
FB1B
FBB0
FBC8
FB7F
FB4E
FB59
FB51
FB13
FAFC
FB62
FBEB
FBDA
FB2D
FB0F
FCC6
002E
0390
0541
0529
0492
0496
0516
054C
04FA
049F
04A7
04D4
04B2
044B
0418
0458
04C5
0504
0513
0526
0539
051D
04DD
04CC
050E
0543
04FD
0466
0426
0488
04FD
04CE
0428
0405
04D5
0584
0457
00E3
FCD4
FA6C
FA52
FB35
FB84
FB0C
FAB0
FAF4
FB65
FB6D
FB2C
FB2D
FB7C
FB9E
FB55
FB01
FB07
FB3E
FB3D
FB0A
FB08
FB46
FB59
FB04
FAAF
FAE7
FB87
FBD5
FB7F
FB16
FB4C
FBEE
FC14
FB59
FA9A
FB3C
FDCE
015C
0438
055B
0518
0491
048C
04E7
050D
04C8
0475
0479
04C0
04EC
04DC
04C9
04D6
04DE
04BE
04A0
04B6
04DD
04C7
047F
046B
04B5
04F4
04B6
0437
0423
049F
04F9
04A0
040B
0439
0529
056A
0381
FFB1
FBFB
FA42
FA99
FB8C
FBC8
FB48
FADD
FAFC
FB5A
FB7A
FB54
FB2F
FB2E
FB2D
FB13
FB05
FB2A
FB64
FB7B
FB71
FB7B
FBA3
FBAF
FB80
FB52
FB69
FB9F
FB8D
FB29
FAF6
FB52
FBCC
FB94
FAA8
FA4D
FBE8
FF6E
0329
0547
056E
04C5
048C
04ED
053B
0503
0496
0479
04AC
04C8
04A7
0492
04BE
04EC
04D0
048F
0491
04D9
04EA
047A
03FE
0411
0493
04C3
0452
03DD
040C
0495
04AA
043A
042D
050B
05E8
0516
0208
FE1C
FB59
FAA1
FB3D
FBE1
FBD5
FB3C
FAA5
FA79
FABD
FB20
FB4C
FB2E
FAF5
FAD8
FAE5
FB09
FB32
FB53
FB62
FB58
FB4B
FB55
FB6D
FB7B
FB84
FBA4
FBC9
FBBC
FB7D
FB68
FBB0
FBDE
FB56
FA71
FAA4
FD19
0124
0493
05C5
051E
044E
0466
0501
0539
04DA
046D
046A
04BE
051A
0556
0575
0561
050A
04A2
047F
04B4
04E9
04CB
047D
046C
04B7
04FC
04D9
047C
0470
04D8
0528
04DF
0451
044E
04E8
04ED
030C
FF6E
FBE6
FA3C
FA83
FB52
FB6D
FAF2
FAC2
FB2D
FB9D
FB7A
FAF2
FAB2
FAFC
FB65
FB6D
FB21
FAF2
FB14
FB48
FB4A
FB32
FB3D
FB5D
FB52
FB1F
FB19
FB5B
FB7E
FB28
FAB6
FAE6
FBB8
FC2B
FB84
FAB2
FBA1
FEFD
031B
0590
05AA
04D6
04B5
0566
05EB
05AE
0518
04BD
049B
046F
0452
0485
04E0
04EC
0494
044F
0482
04F4
051F
04EB
04C0
04EC
052B
0512
04AE
047D
04BB
0500
04C4
042B
03FF
04B9
0594
04F9
0213
FDF1
FAC6
F9DE
FA8D
FB2B
FAEB
FA5E
FA5C
FADB
FB33
FB20
FB0C
FB4B
FB94
FB7C
FB24
FB0C
FB50
FB83
FB56
FB0A
FB0C
FB50
FB69
FB2F
FB00
FB32
FB89
FB8C
FB40
FB34
FBAA
FC12
FBAC
FAB6
FA9D
FCB2
00A0
0469
0627
05B8
04A3
045E
04F8
0581
055E
04E5
04B6
04E9
0515
04FF
04D9
04DC
04E9
04CD
04A4
04B7
0507
0540
0529
04EC
04CD
04C3
048F
0434
0408
0441
048F
0482
043A
045F
051E
0578
03FD
0074
FC76
FA17
F9F7
FAD8
FB2C
FABD
FA76
FAE6
FB83
FB89
FB0F
FACB
FAFF
FB2C
FAE7
FA85
FA9C
FB23
FB79
FB4B
FAF9
FAF8
FB2B
FB2D
FB0C
FB31
FBA9
FBEF
FBA6
FB33
FB48
FBE0
FC25
FB89
FACF
FB82
FE56
0233
051A
05EB
0544
04A1
04D4
0570
05A0
053F
04E4
04F5
052F
0523
04E3
04DB
0521
0546
04FA
0486
046C
04AD
04D6
04AD
0486
04B0
04ED
04D1
0471
044E
048F
04C0
0480
042C
046A
050F
04DC
02BB
FF15
FBB4
FA22
FA5C
FB1E
FB50
FAF4
FAB7
FAEE
FB33
FB0A
FA97
FA6D
FACD
FB51
FB7D
FB51
FB2F
FB3F
FB4D
FB2F
FB0C
FB14
FB2C
FB1D
FB03
FB35
FBA7
FBD2
FB71
FB03
FB2C
FBB8
FBBC
FAF9
FAA1
FC49
0003
03F2
0607
05E7
04F4
049A
04FC
054E
0512
049A
0478
04BD
04FE
04F7
04CE
04C5
04CF
04B3
0471
0454
0487
04DA
0502
04F8
04EF
04EF
04CC
0482
0466
04B3
0508
04C9
040B
03BB
0472
0550
048F
016D
FD3D
FA4B
F9B5
FA9F
FB66
FB56
FAF5
FAF5
FB54
FB94
FB7E
FB5C
FB86
FBE5
FC13
FBD9
FB6C
FB25
FB1F
FB36
FB45
FB45
FB32
FB07
FADB
FAEB
FB4D
FBB3
FBB5
FB61
FB4A
FBBA
FC23
FBBF
FAE0
FB15
FD97
01AA
050D
0621
055B
0476
047A
04FA
0515
04AF
045E
047E
04C6
04CF
04A2
0486
048F
048E
0467
0443
0450
0487
04C0
04F3
0532
0563
0540
04BA
0441
0454
04D6
050F
048E
03DD
03F3
04D4
050F
0321
FF4C
FBA3
FA0C
FA79
FB4F
FB5B
FAE4
FAD0
FB48
FB9B
FB58
FAE7
FAE4
FB48
FB8F
FB82
FB71
FB9F
FBCF
FBA7
FB3E
FB0A
FB39
FB71
FB53
FB06
FB02
FB5B
FB96
FB5C
FB09
FB38
FBCB
FBEA
FB32
FAA5
FBED
FF6C
0377
05CF
05CA
04C2
045C
04E3
0579
0578
051D
04EC
04F4
04F3
04D7
04CE
04DD
04CD
0490
0470
04A0
04E4
04DC
048F
045F
047B
049F
0484
044E
0462
04D1
0523
04E0
043B
03FC
0495
054F
04AE
01E5
FDEC
FAE8
FA35
FB1A
FBBE
FB41
FA78
FA85
FB4C
FBBE
FB61
FADB
FAE1
FB38
FB30
FAC8
FAB3
FB32
FBA1
FB67
FAE4
FADA
FB4A
FB7B
FB23
FAE2
FB4B
FBF0
FBEE
FB43
FAEE
FB83
FC38
FBDB
FAAD
FA86
FCE2
0110
04B4
060E
057E
04B4
04BD
0527
0508
0456
03ED
0454
050D
0542
04DA
047F
04AC
0518
0533
04FE
04F4
0541
0577
0535
04B8
0480
0497
0498
0460
0451
04A9
04FF
04C2
042D
0423
04E2
053A
039E
0001
FC3F
FA53
FA79
FB47
FB74
FB15
FAFE
FB64
FBA2
FB45
FABC
FAB7
FB25
FB54
FAFB
FAA0
FAD0
FB4C
FB69
FB0B
FACB
FB0F
FB75
FB6D
FB1B
FB23
FB9C
FBD2
FB50
FAAD
FAD6
FBB3
FC1E
FB74
FAB4
FBA0
FEC5
02AB
0537
059D
04D4
0452
049A
0522
0545
0508
04E4
050E
0537
050A
04AF
0497
04DC
051C
0504
04C9
04D6
0526
0546
0504
04BF
04D6
050D
04E8
047B
046B
04EA
0540
04C5
03FC
040A
04F0
0506
02B8
FE99
FB18
FA02
FACB
FB89
FB40
FAA4
FABB
FB6E
FBCD
FB62
FAAD
FA65
FA96
FACE
FAD4
FAD9
FB0A
FB3F
FB47
FB3C
FB53
FB78
FB65
FB1C
FAF7
FB2A
FB62
FB3A
FAE0
FAF1
FB8E
FBFA
FB80
FA97
FAC2
FCFF
009E
03D5
055E
055A
04CB
0484
04B0
0506
053B
0529
04E3
049E
0491
04C0
04FF
0522
0525
0519
050C
0508
0514
051E
0507
04DC
04CE
04E3
04E2
04AF
048F
04CD
0524
04F5
043C
03E4
0495
055C
0453
00E2
FCD2
FA89
FA8E
FB5D
FB7D
FB0D
FAFA
FB75
FBC3
FB77
FB0D
FB16
FB6B
FB80
FB37
FAE3
FABD
FABA
FAD6
FB1B
FB5E
FB50
FAF7
FAC2
FAF3
FB42
FB52
FB4F
FB98
FBE5
FB7C
FA88
FA90
FCE9
00EE
0465
05BF
056E
04EB
04EB
0503
04BF
045A
0444
0471
0486
0472
046B
048B
04BC
04F1
052A
053E
04FD
0495
0487
04F9
0561
0527
0482
0438
0489
04D0
048F
0441
0495
050B
0417
00FE
FD10
FA89
FA4F
FB47
FBDD
FBA8
FB4F
FB53
FB81
FB7D
FB4B
FB24
FB16
FB12
FB21
FB4E
FB6C
FB48
FB05
FAFB
FB28
FB29
FADB
FAA9
FAEC
FB57
FB60
FB24
FB3D
FBAF
FBAD
FAF3
FAD0
FCF5
011D
04D4
0600
0513
0426
045B
04FA
04FD
0488
0461
04A4
04B8
046F
044F
04A2
04E6
04A9
044C
0470
04F9
0539
04F6
04AA
04B7
04E5
04E2
04C9
04D3
04D2
0493
0476
04F6
056E
0449
00F0
FCFA
FAAA
FA88
FB2B
FB39
FACE
FABB
FB16
FB47
FB1D
FB10
FB58
FB84
FB44
FAFF
FB2C
FB8A
FB97
FB71
FB95
FBEA
FBBF
FAE9
FA3B
FA74
FB2D
FB74
FB2F
FB1B
FB65
FB43
FA85
FA9D
FD1C
015E
04CC
05A6
04CA
0444
04C6
0551
0513
0494
04B4
0543
0566
04EA
047E
0498
04D8
04BD
0468
0454
0498
04D0
04C3
04A5
04B6
04E8
0514
0532
0529
04CC
044A
044E
051F
05B9
0476
00ED
FCCE
FA5D
FA3E
FB1E
FB85
FB4D
FB24
FB44
FB43
FAF9
FAC7
FAF8
FB42
FB4C
FB3B
FB68
FBAF
FB99
FB21
FAD6
FAFF
FB34
FB13
FAE0
FB0C
FB61
FB4E
FAE8
FAE0
FB59
FB7C
FADB
FABC
FCEA
012B
04E5
05E9
04D9
040F
04A1
057C
0563
04AE
047A
04E6
0504
046F
03EA
042E
04E4
0545
0535
051B
050D
04D2
048C
04B2
053D
0583
0525
04A1
0497
04D5
04BF
047B
04B8
0535
0463
014D
FD31
FA71
FA07
FAD6
FB61
FB62
FB63
FB89
FB7B
FB3C
FB3E
FB8A
FB89
FAFC
FA8D
FACF
FB54
FB4A
FAC5
FA9D
FB26
FBB7
FBAC
FB49
FB27
FB3B
FB0D
FABC
FAE3
FB72
FB79
FABC
FAAE
FCF4
0118
04AD
05DD
052F
0470
047E
04C8
04B4
048A
04C4
052B
0533
04E6
04C5
04F8
051D
04F3
04BE
04C8
04EB
04DB
04A7
0493
04A1
0496
047C
04A4
0504
050D
0490
0444
04D6
0585
0489
0128
FCFA
FA73
FA5F
FB5B
FBBD
FB55
FB00
FB25
FB56
FB34
FAF5
FAEA
FAEE
FAC6
FA9E
FACD
FB30
FB4B
FB0C
FAF1
FB3D
FB8E
FB77
FB33
FB34
FB64
FB53
FB12
FB2E
FBB0
FBC8
FB16
FAD4
FCBF
00C0
048C
0608
0577
04B8
04D3
0535
0514
04A9
049E
04F5
051D
04EF
04D4
0500
0512
04D5
04AB
04E7
0536
0526
04E5
04E5
050F
04E7
0471
0447
0499
04BD
0442
03E9
049B
0594
04B1
011A
FCBD
FA56
FA72
FB44
FB2D
FA73
FA3A
FAC0
FB3F
FB3B
FB06
FB00
FB08
FAF5
FB05
FB5B
FB8D
FB31
FA9F
FA80
FAD9
FB0F
FAE2
FAC0
FB06
FB5E
FB5B
FB44
FBA5
FC2C
FBEA
FAEC
FADF
FD41
0157
04AF
05B2
050F
0480
04C6
054F
056D
052F
0503
0508
0517
051C
050F
04D4
0475
0455
04B7
0547
0566
0507
04C3
04F6
0538
0503
0496
049C
0505
04FB
043A
03C4
047B
056E
047B
00ED
FCB3
FA6F
FAA8
FB92
FB81
FAAE
FA55
FAC8
FB3A
FB14
FAB5
FAB0
FAF4
FB0D
FAEE
FAF2
FB33
FB60
FB50
FB41
FB5D
FB6E
FB46
FB22
FB43
FB66
FB2B
FACD
FAED
FB85
FBBB
FB2F
FB0B
FCEB
00B6
044F
05CD
0566
04C0
04D5
053A
0545
050B
04F9
051A
052C
052A
0544
055F
0526
04AF
047B
04A7
04AA
043F
03F1
044C
04ED
0505
0499
0480
0500
0548
04C1
0435
04BC
05A9
04D3
0149
FCEB
FA68
FA4E
FAF7
FAFE
FAAF
FAE0
FB62
FB5A
FAB2
FA40
FA85
FB00
FB19
FAFF
FB27
FB71
FB75
FB49
FB5C
FBA6
FBA4
FB3B
FAFB
FB45
FBA3
FB7A
FB0A
FB17
FB92
FB8E
FAD3
FAC7
FCF5
00F0
047F
05F1
05A3
0509
04E8
04F6
04DD
04D8
051F
0560
0534
04C4
0483
0488
0494
0497
04C9
051E
052A
04BE
0450
046B
04E7
0522
04EE
04C0
04DB
04D8
0475
043E
04D0
0576
0478
011D
FCF0
FA53
FA0D
FACD
FB13
FACB
FAAF
FAE8
FAFF
FAE1
FB0E
FBAB
FC10
FBB1
FAFB
FAC3
FB17
FB3F
FAF4
FACA
FB2D
FBA5
FB96
FB3C
FB3B
FB8C
FB95
FB48
FB4C
FBCC
FBE1
FAFB
FA61
FC21
0053
0476
0629
05B1
0517
0558
05A2
051A
0444
041D
04A1
04FB
04DC
04C4
04F6
0506
04BE
04AA
0528
0598
052D
043B
03D4
0452
04F2
0502
04BF
04A1
0481
041B
03F3
04BD
05C3
0502
0198
FD3E
FA92
FA4E
FB07
FB5A
FB54
FB84
FBB3
FB55
FAAA
FA8F
FB1C
FB6A
FAF6
FA77
FAC1
FB7D
FBB1
FB41
FAFA
FB40
FB87
FB52
FB0C
FB46
FBB2
FB96
FB18
FB25
FBDC
FC15
FB2B
FA8B
FC52
007C
0478
05E3
0505
0401
0426
04D9
0512
04D5
04CC
050F
052A
04FE
04EC
0515
0516
04B7
0464
0491
04FD
0509
04A8
046D
04A4
04E6
04D6
04B1
04C8
04D9
048F
0452
04D2
0598
04EC
01D0
FD99
FAD4
FA81
FB45
FB72
FAFA
FAD7
FB44
FB84
FB38
FAF2
FB2A
FB76
FB3E
FAC9
FAD8
FB67
FBA7
FB44
FAED
FB30
FB93
FB6E
FB04
FB0F
FB78
FB80
FB0F
FAFB
FB96
FBDC
FAFE
FA31
FBBD
FFE8
0421
05D2
0538
0480
04CB
0540
04FA
0476
049C
053F
0568
04E7
0488
04BF
0500
04CE
0491
04CC
0521
04EF
0473
0476
0502
0540
04CA
0448
0460
04A7
0469
040F
049E
05B8
054F
021B
FDA0
FAB7
FA71
FB51
FB93
FB1D
FAE4
FB35
FB71
FB37
FAEE
FAF5
FB0D
FAEC
FADC
FB2E
FB88
FB5B
FACD
FA90
FAE0
FB32
FB1B
FAF1
FB25
FB7C
FB72
FB31
FB63
FBEC
FBCC
FAB8
FA3E
FC3D
0074
0462
05E2
054C
0488
04A3
0503
04DD
0470
0470
04DC
051C
0503
04F1
050F
0505
04A7
0468
04B9
0547
055E
04F0
04A6
04DD
0520
04F5
049B
048B
04A6
0484
045B
04C8
057A
04D9
01CE
FD80
FA83
FA17
FB07
FB70
FAFC
FAAC
FB05
FB6F
FB50
FAF3
FAF8
FB53
FB81
FB60
FB4B
FB5E
FB43
FAE1
FAB0
FAFC
FB5A
FB44
FAEB
FAE5
FB40
FB86
FB8E
FBA9
FBE2
FBA7
FAD3
FA93
FC6A
002C
03CF
0587
058C
0540
0544
052A
04B5
046C
04B8
052D
0529
04C4
0495
04B3
04A1
043D
0419
0495
0532
054A
0501
04E5
04F9
04C5
044A
042D
04B0
052A
04F6
0487
04C6
055C
0495
016F
FD36
FA5E
F9F4
FADE
FB7A
FB54
FB0C
FB15
FB3F
FB3D
FB23
FB27
FB3D
FB39
FB27
FB30
FB44
FB31
FAFB
FAEA
FB22
FB74
FB98
FB8C
FB82
FB92
FB8F
FB42
FACA
FAB8
FBC6
FE43
01A7
04B0
0632
0602
050F
047E
04A8
050C
051C
04D7
049E
04A0
04BF
04D9
04EF
0502
04F8
04CE
04B8
04DC
0509
04F5
04B1
04A0
04DC
04ED
047D
040F
046B
0543
04F4
023D
FDF7
FA90
F9A2
FA77
FB35
FB06
FA9F
FAD0
FB57
FB76
FB1F
FAF0
FB2D
FB64
FB2C
FAC7
FABC
FB0F
FB52
FB4D
FB42
FB59
FB4D
FAE9
FA96
FAE6
FBB1
FC0B
FB65
FA7E
FAE8
FD80
0171
04CB
0631
05E2
052D
0506
0546
0542
04D0
0480
04C2
0544
0562
050D
04D0
04F6
0521
04F1
04A6
04B6
0502
04FC
0494
0468
04CE
052F
04D9
043C
0479
0587
059C
0314
FEA3
FAE6
F9B1
FA68
FB24
FAF3
FA77
FA86
FB04
FB3F
FAFE
FAB1
FAB3
FADC
FAE3
FACC
FAC8
FAE0
FAEC
FAE4
FAF3
FB35
FB6F
FB55
FB04
FAFD
FB74
FBD8
FB6F
FA80
FA8C
FCE5
010D
04CB
0637
0584
047B
046E
050F
0562
052B
0501
0539
0578
055E
052B
0552
05B0
05AE
0520
0498
049E
04F6
0501
04A9
0475
04B9
0512
0505
04C5
04EB
0565
0512
02DC
FF21
FBAD
FA1E
FA64
FB26
FB53
FB12
FB0C
FB4B
FB3A
FA97
F9F9
FA12
FABD
FB2D
FAFA
FA92
FA83
FAC4
FAF1
FAFD
FB2E
FB7E
FB85
FB1D
FAC5
FAFA
FB64
FB38
FA86
FAA6
FCD7
00A7
041F
05A7
0567
04C4
04BF
052A
0550
0502
04B5
04CE
0525
054C
0526
04FC
0509
0531
0535
0509
04DB
04C7
04BB
04AB
04B1
04DA
04EC
04B5
047D
04CA
0578
0561
0365
FFC8
FC40
FA66
FA56
FAE8
FB25
FB0C
FB0C
FB29
FB13
FAC7
FAA9
FAE9
FB30
FB11
FAA3
FA6C
FAB3
FB2B
FB60
FB46
FB34
FB57
FB78
FB5F
FB31
FB3A
FB60
FB32
FAB2
FACD
FCA2
0023
03BC
05A4
058E
04C2
0494
0511
0569
052C
04C2
04AD
04E3
0503
04FA
050A
0543
0561
053B
0506
0504
0518
0502
04CB
04BB
04D4
04C2
0469
0440
04C4
0593
0568
0348
FFAC
FC3E
FA71
FA54
FADC
FB14
FAE9
FAD7
FB16
FB55
FB42
FB06
FB04
FB3B
FB43
FAEA
FA91
FAA7
FB0A
FB34
FAFC
FAC8
FAED
FB30
FB2B
FAFE
FB1D
FB71
FB4B
FA8A
FA5B
FC32
0001
03E8
05FA
05F6
0529
04CA
04EF
050D
04F6
04E9
0502
0505
04D1
04AE
04E9
055B
0584
0528
0499
0456
0484
04DC
051F
0551
057B
0569
04ED
045E
046D
0539
05A8
0437
009D
FC7A
FA03
F9EF
FB03
FB9D
FB57
FAF0
FAFB
FB34
FB21
FADD
FAD6
FB14
FB2C
FAF0
FABF
FAEE
FB41
FB42
FAFB
FAE6
FB23
FB3A
FAD2
FA61
FA9F
FB6E
FBCE
FB31
FA93
FBAD
FEFD
02F9
0585
05F1
0549
04E0
04F2
04F6
04B8
04A2
04F7
054D
0521
04A7
048B
04F2
053D
04EC
0461
045E
04F7
0576
0559
04F6
04E8
0522
051B
04C9
04D6
0586
05D7
044E
00BD
FCCA
FA75
FA3E
FAFF
FB64
FB2E
FAF9
FB20
FB4B
FB16
FAAD
FA93
FAE6
FB40
FB45
FB1C
FB23
FB61
FB7C
FB4B
FB16
FB25
FB3E
FAFF
FA91
FA90
FB1D
FB73
FAEF
FA54
FB5C
FEBF
0300
05B1
05DC
04C3
042D
0486
04F7
04E4
04A5
04BE
0510
0523
04F0
04E5
0527
054B
04FD
048A
0478
04C2
04DF
049D
0474
04CA
0541
0523
0476
0428
04CE
0587
04A3
0187
FD94
FAE5
FA49
FAD0
FB2D
FB17
FB15
FB60
FB88
FB3A
FAD5
FAE9
FB5D
FB88
FB22
FAAF
FAC2
FB35
FB6E
FB41
FB21
FB5D
FBA5
FB89
FB32
FB2C
FB82
FB87
FAD6
FA4A
FB66
FEA1
029A
053E
05B3
04F6
0490
0501
058E
0570
04C9
0455
0470
04C6
04E9
04DD
04E9
0518
052E
050C
04D8
04B0
0482
044B
0450
04B9
051A
04D6
0418
03E8
04D8
05E0
0517
01D6
FDA7
FADA
FA42
FAC5
FAF6
FAA2
FA85
FAF1
FB5F
FB46
FAE2
FACF
FB29
FB70
FB42
FADE
FAC6
FB0E
FB50
FB4A
FB33
FB51
FB89
FB8C
FB65
FB7A
FBD0
FBCC
FAFE
FA26
FAE5
FE08
024F
0567
0618
0545
04A1
04DC
055E
0575
0539
0520
0533
051D
04D2
04B1
04E8
051A
04E8
0488
0479
04C5
04EF
04AB
044F
0454
04A3
04B8
047B
047C
0521
05B4
04D0
01D9
FDE7
FAEC
F9FD
FA85
FB23
FB16
FAB0
FA90
FABF
FAD8
FAB6
FAAB
FAED
FB32
FB15
FABA
FAB0
FB2F
FBBB
FBC3
FB60
FB20
FB37
FB45
FB0E
FAF8
FB6E
FC06
FBE6
FB20
FB2B
FD68
0155
04BE
05F3
055A
04AC
04DD
0568
0570
0505
04D6
051C
0557
052D
04EC
04F7
051F
04F4
0495
049B
052A
058F
052C
0465
0433
04C2
0525
04A9
03F0
0422
0523
0530
02C9
FE94
FAF4
F9B5
FA6E
FB5A
FB5A
FACE
FA9D
FAF8
FB4D
FB30
FAE0
FAD6
FB1A
FB48
FB26
FAF2
FAFA
FB2B
FB34
FB03
FAE0
FB00
FB3C
FB5F
FB83
FBD2
FBFE
FB7B
FA83
FA85
FCE3
0125
04FB
0665
05AA
04C0
04EA
0590
0583
04C1
0459
04C9
0550
0524
0498
0494
0527
056E
04EE
0457
048E
0557
05A5
050F
0460
0460
04C0
04B1
0445
0465
053B
055E
033A
FF1D
FB49
F9B6
FA32
FAFD
FAED
FA72
FA80
FB27
FB9F
FB71
FB08
FAFB
FB39
FB41
FAF7
FAD0
FB16
FB6F
FB5C
FAFB
FAE0
FB37
FB78
FB3A
FAE2
FB15
FBA8
FBA9
FADA
FA92
FC85
009F
04AA
0675
05FD
0513
050F
058A
0570
04AD
043D
04A9
0550
0556
04D6
0499
04E0
0515
04BE
0449
0467
0502
0554
0501
0492
049D
04D9
04A0
0417
042E
0522
0592
03BE
FFAC
FB8A
F999
FA04
FB11
FB45
FAC3
FA89
FAE9
FB42
FB15
FABA
FAC8
FB34
FB73
FB4B
FB1C
FB35
FB57
FB1F
FABC
FAC1
FB46
FBAD
FB78
FB0D
FB2A
FBBB
FBD3
FB14
FAB1
FC5A
0026
0415
05FF
05BC
04F4
0500
058C
058D
04E8
0489
04F5
0585
055E
04AC
0453
04AB
0511
04F6
04AF
04DE
055C
055D
04AE
0420
0467
050F
051A
047F
0448
04EF
0549
03A4
FFEC
FC10
FA15
FA28
FAE3
FB18
FAD5
FABA
FAEA
FB08
FAEB
FAD8
FB00
FB2C
FB14
FAD4
FACA
FB10
FB5C
FB65
FB3E
FB1E
FB10
FAFF
FAFF
FB4D
FBE3
FC39
FBC1
FABB
FA62
FBF5
FF75
035C
05CD
0627
0564
04EC
0529
0573
0530
04A8
048C
04F5
054E
052D
04E1
04E5
051D
050A
049E
045F
049C
04F0
04E2
04AA
04CC
052D
0520
0489
0448
04EC
0561
03D2
0004
FC12
FA45
FAA8
FB5D
FB14
FA60
FA68
FB25
FB8D
FB2E
FAB7
FAD9
FB4F
FB6C
FB22
FAEE
FB02
FB15
FB02
FB04
FB3D
FB69
FB51
FB34
FB51
FB5C
FAFB
FAD0
FC3C
FF9A
0354
0556
053D
048E
04BB
059C
0615
05B0
050A
04CA
04E6
04FE
04F4
04DE
04BC
0496
04A3
04F1
0526
04F4
049E
049C
04D3
04AF
0435
0447
054B
05E1
040C
FFCC
FBA3
F9FE
FA9C
FB55
FAF2
FA47
FA78
FB3A
FB70
FAED
FA9B
FAFA
FB6C
FB48
FAE4
FAEB
FB40
FB48
FAF4
FAD2
FB16
FB56
FB52
FB60
FBA5
FB88
FAAE
FA4C
FC40
008D
04A8
060F
050C
0405
046F
0573
05A1
0501
04B4
0527
059B
056D
04FB
04DE
04FE
04F1
04C4
04C9
04EA
04D7
04AE
04D8
0537
052E
04A5
0473
0508
0531
032C
FF1F
FB77
FA49
FB0B
FBAB
FB3D
FAAF
FAEB
FB78
FB66
FACB
FA89
FAD9
FB0F
FACC
FA9A
FAF0
FB5C
FB3F
FADC
FAE4
FB47
FB4E
FAD2
FA8B
FAD6
FB04
FA9A
FAAD
FCEA
011E
04D3
05F0
0512
046D
04F2
059C
055A
049C
0474
04F5
0541
04F6
04A9
04DD
053B
0539
04EE
04C6
04C9
04C0
04C0
04FE
0539
04FC
048D
04CA
05B4
05B1
0322
FEB1
FB0D
FA13
FAF0
FB8E
FB27
FAA4
FACB
FB32
FB29
FAD9
FADA
FB2A
FB35
FAE0
FAB8
FB0B
FB62
FB4B
FB0F
FB1E
FB48
FB21
FAE2
FB16
FB80
FB30
FA2E
FA40
FD1C
01F2
05BC
066C
04FF
03F2
0451
051C
0531
04C1
049A
04E0
0513
04FD
04EF
0515
0527
04F3
04BA
04B9
04C4
04AE
04B3
0501
0536
04E0
0465
04A2
056C
0526
027B
FE49
FB04
FA21
FAC1
FB34
FB06
FAF6
FB60
FBAF
FB63
FAD7
FAB1
FAF1
FB14
FAF3
FAE0
FB0B
FB33
FB31
FB3D
FB71
FB77
FB27
FAFA
FB57
FBB9
FB48
FA70
FAF9
FE07
0252
053F
059E
04B1
0448
04AC
04FA
04D5
04CF
0541
05A1
055A
04BA
0483
04DA
052A
050B
04BC
0496
0493
04A0
04DC
0531
0523
0487
0429
04D3
05CA
050B
0194
FD07
FA35
FA2D
FB5E
FBCD
FB3D
FAC3
FAEB
FB30
FB16
FADC
FAE6
FB0E
FAF9
FAC1
FACA
FB0D
FB24
FB05
FB1A
FB7C
FBAF
FB6F
FB39
FB78
FBA4
FB05
FA43
FB32
FEA5
02F8
0596
05B6
04DC
04A5
0502
0507
049E
0480
04E6
0535
0509
04DC
052A
059A
0583
04FF
04C8
0509
051F
04B5
045A
048C
04D1
047F
0402
0457
0530
04AC
018C
FD21
FA30
F9F5
FB13
FB9B
FB3D
FAF2
FB2E
FB71
FB4E
FB10
FB10
FB16
FACB
FA65
FA60
FABC
FAFF
FAFE
FB0A
FB3F
FB43
FB03
FB10
FBAF
FC19
FB79
FA99
FB82
FF11
037C
0602
05DC
04C1
0485
051C
0562
04FD
049B
04B3
04EC
04E6
04DB
0523
0580
057A
051D
04E5
04F6
04F6
04C6
04BF
04FA
04F6
0471
041F
04A9
0545
0424
00AD
FCA2
FA6A
FA7D
FB43
FB4C
FAD5
FAD0
FB40
FB64
FB00
FAA4
FABA
FAF6
FAFA
FAF3
FB23
FB48
FAF8
FA77
FA80
FB2E
FBBA
FBA1
FB5A
FB75
FB8E
FB11
FAAF
FC15
FFC4
03E0
05F1
058B
047A
0464
0508
053A
04C4
0480
04E4
055F
0544
04BC
0471
04AD
0527
057C
0586
0547
04DE
04A0
04C0
04E7
0487
03DD
03F1
0514
05C8
040F
FFDF
FBA4
F9D3
FA70
FB7D
FB81
FAE2
FAB4
FB1B
FB6B
FB56
FB2F
FB29
FB0E
FAC6
FA9D
FACE
FB1A
FB2C
FB25
FB53
FB8B
FB62
FAFE
FB09
FB91
FBB5
FB05
FAB6
FC82
0060
041C
05A6
0536
04A4
04F7
0579
0532
0462
03FF
0456
04DD
052C
055C
058B
0585
0531
04D9
04BB
04A6
0461
0432
047E
04FA
04EE
046A
0468
0533
055B
032E
FF0D
FB70
FA42
FAEA
FB6F
FB02
FA92
FAFB
FBB7
FBCF
FB4B
FAF8
FB18
FB22
FAC5
FA6D
FA94
FB12
FB71
FB99
FBB2
FBA2
FB37
FAC6
FAF0
FB92
FBAF
FAF5
FAC5
FCD5
00EE
04BC
0636
059B
04B6
04A5
04FB
04F4
04A4
0490
04CD
0504
0512
0517
050C
04D5
0499
04AA
04F2
04F4
0493
045A
04AF
0505
049C
03DF
0416
0555
05AB
0334
FEA5
FADC
F9CE
FAB1
FB69
FB23
FAB5
FAE8
FB54
FB4A
FAF1
FAE8
FB39
FB60
FB28
FAEA
FAE9
FAFD
FAFC
FB14
FB64
FBAA
FB9E
FB80
FBAF
FBD8
FB57
FA88
FB03
FDD1
01D4
04BB
056F
04FA
04E2
0559
058A
0524
04BF
04D1
04FE
04D4
0496
04BD
0522
0539
04EF
04BD
04D2
04D2
048A
0462
04AC
04F3
049A
0408
0445
053C
0527
0289
FE4B
FB03
FA36
FAF9
FB69
FAE5
FA42
FA49
FAC8
FB2C
FB4E
FB5A
FB51
FB24
FAFD
FB05
FB0F
FAEA
FADC
FB47
FBEC
FC07
FB66
FAE0
FB31
FBC8
FB83
FA9F
FAFB
FDDA
0205
04F1
057F
04E0
04BB
054C
05B1
0575
050F
04F5
0503
04FF
050B
0542
0551
04FA
049C
04B0
04F9
04D3
0444
0416
04A7
0534
04F8
0471
04B4
0575
04D3
01B4
FD8D
FAEC
FAA2
FB36
FB20
FA90
FA8B
FB1F
FB5D
FAE2
FA6B
FAA0
FB20
FB35
FAEE
FAD1
FAE7
FAD7
FAB9
FB0B
FBAF
FBC9
FB02
FA58
FADE
FC01
FC21
FB17
FAFD
FDAF
022D
0583
0612
0506
046E
04CE
0539
0517
04DB
04FB
052D
0512
04E9
0517
0561
054F
04F9
04E1
0516
051E
04D2
04A7
04DD
04F1
0479
0419
04B7
05AD
04E7
016E
FD0A
FA85
FAA1
FBA0
FBB3
FAEF
FA7D
FABC
FB04
FAEF
FADF
FB17
FB30
FADD
FA93
FAD4
FB50
FB5F
FB19
FB24
FB8D
FB94
FAF0
FA71
FAD4
FB73
FB32
FA89
FB79
FEEB
0313
0555
0542
04AB
0502
05C7
05C6
0500
047C
04A8
04EB
04D0
04B6
04F8
052F
04EA
047E
047E
04C7
04CB
04A0
04E3
0583
0589
049F
03FB
04C7
05F7
04FF
010B
FC72
FA22
FA65
FB27
FAF5
FA6B
FA9E
FB52
FB89
FB27
FAFD
FB51
FB72
FAFB
FA9B
FAFF
FBB8
FBE3
FB7F
FB40
FB53
FB30
FABF
FAB4
FB5D
FBD1
FB38
FA82
FBB5
FF49
0337
053F
0556
0514
0553
057F
0511
048E
04A1
0501
04FB
04AA
04BD
052A
0516
0444
03B1
0432
0522
0556
04CF
048E
04E3
04F9
0467
0419
04D9
0588
040A
0026
FC3A
FA91
FADF
FB34
FABF
FA68
FAF2
FBAF
FBA6
FB12
FAF3
FB7C
FBD8
FB81
FAFD
FAF0
FB2C
FB33
FB22
FB5F
FBBB
FBA4
FB2A
FB00
FB5F
FB8F
FB20
FB08
FCBB
0024
0365
04E3
04EF
04E4
0540
056A
0509
049E
04A2
04CC
04A2
045C
048E
051D
0545
04B4
0419
0426
049C
04CD
04AA
04B7
050D
0530
04F5
04E6
0542
050F
02F6
FF1D
FB85
FA14
FAAD
FB9E
FBAA
FB13
FAC0
FAFB
FB57
FB73
FB64
FB64
FB72
FB6C
FB57
FB59
FB76
FB84
FB64
FB28
FB0A
FB29
FB5B
FB46
FAE2
FAEA
FC75
FFC2
0389
05E3
060F
051E
04AF
0538
05D4
05AB
04F6
0478
0469
0464
0433
041C
0456
0493
0477
0435
044D
04BC
04E9
048D
0447
04CD
05AB
0561
02F1
FF23
FBE6
FA8E
FACB
FB5C
FB6E
FB24
FAFC
FB10
FB1A
FAF5
FADD
FB13
FB7F
FBC0
FBAB
FB7D
FB7D
FB98
FB83
FB3E
FB2D
FB82
FBC7
FB62
FA9D
FAD1
FD1E
00FF
0476
05D8
0551
046B
0454
04D2
0507
04B1
0464
0499
0504
0510
04AD
045E
046E
0490
046A
0437
0473
0508
0536
0499
03E1
0412
0505
051A
02E3
FEEB
FB6A
FA1E
FAB4
FB76
FB52
FABC
FAAF
FB51
FBE0
FBC3
FB3D
FAF1
FB16
FB5C
FB83
FB9F
FBC1
FBB6
FB50
FADA
FAEB
FB9E
FC35
FBDF
FAE8
FAD6
FCFC
00EE
0493
0608
055B
0448
0447
0525
05A2
051F
0448
040C
0477
04DA
04D8
04C0
04E6
050E
04D6
046E
0464
04BE
04D3
0447
03C9
043F
054A
0531
02AF
FE97
FB36
FA19
FAB8
FB72
FB64
FAFF
FAFA
FB50
FB78
FB46
FB1D
FB46
FB7E
FB56
FAE5
FAB1
FAFC
FB63
FB65
FB1E
FB21
FB9A
FBEC
FB79
FAB8
FB1B
FD98
0168
048D
05AE
053F
04B5
04DA
0535
050D
0482
0455
04CE
0554
053F
04BA
047D
04C9
051B
04F4
0495
049B
0509
0538
04CE
045C
04A4
0546
04CB
022F
FE46
FB24
FA24
FAC2
FB73
FB5A
FAE3
FACF
FB29
FB5F
FB22
FAC5
FAB9
FAF7
FB2A
FB39
FB5E
FBA3
FBB2
FB45
FAB2
FA9E
FB20
FB80
FB19
FA74
FB0D
FDC6
01BC
04E3
05E8
0549
048B
048F
04FB
0518
04DB
04C9
0518
0560
053F
04E3
04BD
04D0
04B4
0455
0436
04BB
056B
0566
04A6
043A
04EE
05F3
0568
026A
FE48
FB4E
FA8A
FB11
FB5B
FAFA
FAA0
FAE0
FB5F
FB73
FB0D
FAC0
FAE5
FB31
FB33
FAFE
FB06
FB69
FBB2
FB78
FB00
FAE8
FB4D
FB7E
FAEB
FA2E
FAC5
FD87
0178
0483
0569
04D1
0459
04C4
056A
0560
04B7
044D
0497
0516
0524
04D8
04C6
050B
051A
049F
041E
044F
0508
0559
04D4
0445
04A1
057B
051D
026E
FE69
FB50
FA73
FB1F
FBB7
FB80
FB00
FAE8
FB26
FB39
FB02
FAEB
FB2D
FB77
FB5F
FB08
FAFB
FB5C
FBAC
FB72
FAF4
FAE5
FB65
FBAE
FB1B
FA55
FAFF
FDF1
0201
04F2
0598
04D5
0455
04B9
0543
052A
04B1
049D
050F
0559
0504
047D
0476
04E1
050B
04A0
0428
0448
04CD
04FB
04A8
048B
0529
05BC
04B8
0191
FD9D
FAF6
FA7C
FB36
FB9C
FB35
FAB5
FAD2
FB57
FB88
FB26
FAB1
FAAE
FB04
FB34
FB1E
FB1E
FB75
FBCE
FBA4
FB0B
FAAE
FAED
FB4E
FB24
FABF
FB7D
FE4A
0247
054D
05FC
04FF
0425
0463
0516
0530
04AA
0462
04D6
0582
05A2
052D
04BB
04A0
049C
0479
0482
04FE
0588
0566
04A2
0435
04C7
057C
04A1
0190
FDA2
FAF0
FA52
FAE7
FB5C
FB49
FB23
FB3D
FB5E
FB35
FADD
FAB3
FACD
FAF0
FAF3
FAFA
FB2D
FB5D
FB2F
FAAE
FA69
FAD3
FB93
FBBB
FAF0
FA31
FB25
FE60
0281
054F
05D2
0513
04BB
0540
05B8
054E
045F
03F7
0478
0539
0576
0533
04F8
0507
0523
0514
04FA
04F9
04F1
04B4
0480
04CC
058D
05CB
0461
012E
FD7A
FAF1
FA3C
FAA0
FAF4
FACF
FAA9
FAF7
FB76
FB8D
FB2C
FAE4
FB17
FB69
FB4E
FAD9
FAA6
FAEE
FB2E
FAF6
FAA6
FAED
FB98
FB9F
FAA4
F9ED
FB43
FEDD
02EF
055E
05AD
04FE
0498
04C7
051F
0549
053E
050D
04C9
04A2
04C7
051B
0542
0509
04AC
049B
0501
057F
057F
04D7
041E
0434
053B
0601
04D5
0143
FCFA
FA6D
FA73
FB97
FBEC
FB22
FA71
FABA
FB72
FB9A
FB1F
FAC0
FADB
FAFE
FACB
FAA4
FB02
FB8B
FB7C
FAD1
FA71
FAFA
FBCA
FBC3
FAD0
FA51
FBB7
FEF3
0276
04A2
051B
04B9
047D
04B0
04ED
04D6
0491
0489
04D5
051C
051B
0503
051A
0545
052C
04D6
04BB
050F
054B
04D7
0410
040B
050B
05BB
0469
0105
FD5E
FB5B
FB38
FBB9
FBC1
FB4E
FB01
FB1B
FB47
FB2B
FAE1
FABB
FAE1
FB29
FB4D
FB34
FB05
FAEA
FAE1
FAD9
FAED
FB44
FBAA
FB90
FAD2
FA65
FBBC
FF25
0301
0521
04F6
03FC
03E5
04C4
0574
0551
04ED
04FC
0550
0543
04CD
0495
04EB
054C
0529
04C2
04C0
0529
054A
04C7
0442
049C
05A0
05DE
0409
0068
FCBD
FABC
FAA3
FB4E
FB85
FB13
FAA1
FAB7
FB1C
FB44
FB10
FAE7
FAFD
FB06
FAB2
FA4E
FA71
FB26
FBC1
FBB4
FB42
FB0A
FB1B
FAE5
FA4E
FA59
FC41
FFEC
03A5
059B
0586
04AD
0466
04DB
053C
0500
0484
047C
0506
0591
05A2
055A
0525
051D
04FE
04B3
0493
04D9
0529
0504
0499
04AC
0560
0586
03B6
000F
FC6D
FAAB
FAE2
FBA3
FBB1
FB28
FAD7
FB08
FB48
FB25
FAC0
FA84
FAA1
FAE8
FB18
FB25
FB22
FB19
FAFD
FADB
FAE8
FB41
FB9D
FB77
FAC5
FA7E
FC00
FF8D
0388
05BD
058C
046A
0418
04B8
0521
04BB
0445
049D
0564
0591
04FF
04A3
0511
0594
0541
0468
0429
04CA
054D
04E2
0432
047C
05A9
05F9
03E7
FFF4
FC39
FA62
FA6C
FB2E
FBA8
FBA5
FB75
FB5C
FB58
FB43
FB13
FAE8
FAE3
FAF7
FAFF
FAF3
FB01
FB3D
FB75
FB6E
FB50
FB72
FBB3
FB6F
FA89
FA28
FBD7
FFAD
03BE
05CB
0572
044C
03FF
0499
050E
04D3
0466
0464
04B4
04E0
04E2
050E
0561
0557
04B8
041D
0447
0507
0552
049D
03C2
040D
0570
0616
0430
000A
FBFF
FA3D
FAC9
FBDB
FBED
FB25
FAA8
FB07
FBB6
FBEA
FB8D
FB26
FB10
FB24
FB27
FB25
FB45
FB61
FB32
FAD6
FAD4
FB5B
FBD1
FB73
FA85
FA7A
FC91
0054
03CC
0560
053A
04BC
04C7
0502
04C9
0447
0435
04BA
0523
04DF
0459
0464
050E
057E
0521
0477
045B
04D2
0509
0496
0421
0486
0572
056B
0353
FFAE
FC3A
FA64
FA40
FAE6
FB71
FB8E
FB65
FB32
FB13
FB0B
FB15
FB22
FB20
FB11
FB0D
FB2B
FB5A
FB68
FB44
FB21
FB44
FB9F
FBBC
FB46
FAAC
FB07
FD1A
0072
039D
0558
0581
04FA
04B4
04EC
053D
0540
04F9
04B3
049C
04A2
04A0
0497
04A3
04CC
04F4
0507
0518
052E
0518
04B9
046A
04AB
0542
04F2
029E
FEC4
FB6F
FA4C
FB02
FBC9
FB7C
FAA8
FA70
FB00
FB93
FBA4
FB7C
FB7D
FB7D
FB2D
FAC2
FAB5
FAF4
FAF4
FA9E
FA9D
FB52
FC05
FBC8
FB15
FBBB
FEC9
02F7
05C8
0618
050D
0476
04D0
0542
051A
049F
0464
0477
048E
04A1
04DF
0532
0544
050D
04F5
052A
053F
04CE
044D
0485
0534
04C3
0202
FDE3
FAD4
FA3C
FB1E
FB8B
FAEB
FA4F
FAAA
FB8D
FBF1
FBA0
FB4B
FB58
FB66
FB17
FAB6
FAAD
FAD9
FAD7
FACB
FB22
FBA0
FB70
FA8B
FA7E
FCDF
011D
04A7
05A1
04C5
0427
04A1
054A
0536
04BF
04B2
04F5
04D6
0450
042E
04BD
0540
050A
0494
04B3
0536
0525
046B
0436
052E
05F4
0461
0048
FC10
FA35
FAC2
FBCA
FBE5
FB63
FB21
FB2E
FB14
FAD9
FAFD
FB83
FBBE
FB53
FADB
FB0F
FBAF
FBD7
FB58
FB07
FB69
FBC5
FB2D
FA3E
FAEC
FE3A
02A8
0580
05A4
0474
03EC
0475
0504
04E2
0481
0488
04CD
04C2
046A
0454
04A7
04DA
0493
043E
0462
04B9
04A2
0446
0484
0564
055C
02EC
FEB8
FB41
FA4A
FB19
FBAF
FB3E
FAAA
FADD
FB82
FBBF
FB85
FB72
FBB0
FBBB
FB50
FAF3
FB23
FB8B
FB88
FB34
FB48
FBDC
FC12
FB63
FAD9
FC27
FF8B
033D
053E
0559
04E7
04F7
0549
052A
04A3
0457
0482
04B1
048F
0466
0493
04E2
04D7
0483
0476
04D5
0503
0485
03EB
0423
04EA
048F
01DA
FDCB
FACE
FA31
FAF1
FB4E
FAE4
FAA4
FB25
FBC2
FBAE
FB27
FAFF
FB51
FB70
FB1B
FAEA
FB52
FBC7
FB94
FB0C
FB19
FBB4
FBBD
FAD1
FA80
FCB7
0118
04E2
05EC
04E4
0418
0491
0555
054A
04C5
04B4
0519
0523
049E
044C
04AF
052F
0508
0478
0453
04B1
04D0
0473
0469
0532
05AC
040C
0033
FC4E
FA96
FB06
FBCA
FB9F
FAFD
FAD5
FB10
FAF3
FA76
FA6A
FB30
FC04
FBFA
FB42
FACF
FB03
FB4B
FB2F
FB0B
FB50
FB94
FB23
FA77
FB38
FE45
0244
04D6
051B
0469
046A
0527
057F
0506
0490
04D5
055D
0541
0487
040F
044B
04B5
04BF
04A0
04D0
0518
04E3
045B
0464
0526
053D
0322
FF3E
FBD3
FAA4
FB31
FBA8
FB28
FA74
FA7F
FB1E
FB78
FB48
FB0B
FB1C
FB44
FB48
FB5D
FBB7
FBFF
FBC6
FB48
FB3F
FBB7
FBCD
FAFE
FA60
FBBC
FF59
0346
0547
051E
0470
048F
052D
054C
04DA
049D
04E9
0526
04D8
046E
048F
0505
0500
045B
03E4
0424
0491
046C
040C
0465
053F
04DB
01F9
FDC5
FAE1
FA8E
FB7E
FBC2
FB17
FAB0
FB24
FB9F
FB44
FA86
FA79
FB3A
FBCD
FB98
FB26
FB35
FB9B
FBAD
FB74
FB8E
FC02
FBF4
FB1C
FAD0
FCCA
00D1
0485
05D0
050F
0447
049C
0556
0557
04B8
046E
04D1
0542
0530
04D3
0499
047C
0449
0438
0497
0505
04C3
03E9
03A4
049D
058C
044D
007A
FC49
FA44
FAAA
FB96
FB81
FAC0
FA77
FAE0
FB44
FB3D
FB2C
FB59
FB71
FB2D
FAFB
FB62
FC0B
FC17
FB70
FB0A
FB7C
FC00
FB8A
FAA1
FB3B
FE63
02A1
055B
0593
049F
0445
04CB
0544
0526
04D9
04D5
04E5
04A2
0444
0453
04C7
04FB
0496
0410
0408
0467
049E
049C
04DA
0555
04F5
029E
FECA
FB77
FA3D
FAC4
FB6E
FB4A
FAD6
FAE3
FB5F
FB97
FB58
FB2E
FB80
FBEE
FBE5
FB78
FB38
FB56
FB76
FB62
FB5F
FB90
FB7C
FAD4
FA7C
FC00
FFAB
03A7
05B2
0576
04AA
04C8
056E
055F
047D
03ED
0460
051F
0519
0463
03FB
0450
04CE
04DD
04AA
049D
048D
0432
03FB
0497
058A
0508
01F3
FD93
FA93
FA32
FB26
FB78
FADF
FA8C
FB26
FBE7
FBD8
FB34
FAEF
FB4B
FB99
FB5F
FB01
FB0C
FB5F
FB86
FB87
FBBF
FBFD
FB94
FAA2
FAA5
FD08
0138
04D4
060D
055F
049C
04B8
0521
050D
04A7
0486
04AB
04A2
0467
0481
0509
054B
04C9
0417
041D
04BE
04F4
046A
0425
04EF
05A6
0431
0030
FBEB
F9F2
FA6E
FB61
FB51
FAB1
FA9B
FB16
FB53
FB1B
FB0F
FB74
FBA6
FB37
FACB
FB30
FC05
FC1C
FB45
FAAC
FB2A
FBE6
FB8B
FA83
FAF5
FE23
028B
0570
05C8
04FC
04CB
055C
05B0
0551
04D6
04D2
0511
0510
04C9
0496
0490
047F
0465
0486
04DC
04E9
046F
0408
0472
0559
0539
02E9
FF11
FBB3
FA42
FA70
FAEE
FAF8
FAC9
FACC
FAF2
FAEE
FACD
FADC
FB2A
FB67
FB66
FB58
FB6A
FB69
FB26
FAF6
FB55
FBFF
FC03
FB1A
FA8A
FC0A
FFB1
0392
059D
059C
04F4
04C5
04F4
04FF
04FC
0542
0598
056E
04CD
046E
04AF
04FF
04BC
043B
044F
04F3
052B
047A
03D4
0454
055D
04DC
01B9
FD67
FA82
FA23
FB12
FB8D
FB29
FAB6
FAC4
FB02
FAFC
FAD9
FAF8
FB43
FB59
FB32
FB33
FB7C
FBA3
FB59
FB09
FB44
FBC6
FBA3
FAC5
FAAB
FCF3
0135
04FF
0643
0562
0464
048A
053E
0568
04F4
04AC
04E3
0521
0504
04D2
04DF
04F4
04BD
046F
047A
04BA
04A5
044D
0488
0592
060C
042D
0002
FBD0
F9D6
FA22
FB03
FB38
FAF7
FAED
FB1E
FB1D
FAEA
FAE8
FB27
FB3E
FB03
FAE5
FB3E
FBB2
FBAA
FB43
FB28
FB7E
FB83
FAB6
F9FC
FB02
FE55
027E
0553
0601
057A
050A
0504
04F8
04C1
04BF
051C
056F
054A
04E0
04B8
04DC
04D3
0473
0448
04BC
054A
0525
0484
0485
056D
05B3
0391
FF5C
FB83
FA06
FA7C
FB0D
FADB
FA9A
FAF9
FB7D
FB57
FAB8
FA7D
FAE4
FB50
FB5F
FB66
FBA9
FBAF
FB09
FA50
FA88
FB83
FBCF
FABE
F9D5
FB48
FF44
0376
058A
056D
04CB
04D7
0545
0556
0510
04FD
0535
0547
04F9
049A
0477
0477
046E
0487
04F6
0571
056B
04E7
04B5
055C
0609
050D
01C5
FD9E
FADE
FA72
FB41
FBA9
FB35
FAA5
FAA0
FAEB
FB07
FAFF
FB2F
FB85
FB8D
FB38
FB04
FB32
FB4F
FAEB
FA73
FAAA
FB61
FB81
FAB5
FA7D
FCA8
00E6
04AD
05E2
0505
0430
047D
0530
054A
04EE
04DE
0524
051F
04A8
0459
0498
04F5
04EE
04C4
04F9
054D
0503
043B
041C
052E
060C
049C
009D
FC50
FA36
FA8E
FB87
FB9A
FAF9
FAA8
FAED
FB32
FB10
FAD9
FAF9
FB4F
FB76
FB60
FB55
FB5F
FB3C
FAF0
FAF3
FB74
FBC6
FB2D
FA3B
FABD
FDCE
023F
0579
060C
04F7
0439
048D
051E
0515
04B2
04A0
04E3
0501
04DC
04CA
04E1
04C8
046C
044F
04C4
053D
0508
048A
04D1
05BA
0579
02A8
FE58
FB39
FAAE
FB91
FBEF
FB56
FAC3
FADE
FB30
FB24
FAEC
FAFA
FB33
FB38
FB1D
FB37
FB72
FB71
FB42
FB49
FB78
FB3D
FAA5
FAFD
FD83
0186
04B6
058A
04C8
0436
047A
04EF
0500
04DE
04D8
04D4
04B6
04B8
0509
0552
0526
04B3
0488
04A9
0497
0455
0489
0521
04B0
0204
FE05
FB0D
FA66
FB18
FB7A
FB2E
FAFC
FB42
FB71
FB21
FACA
FAEF
FB49
FB54
FB2A
FB2E
FB4F
FB3B
FB0E
FB1E
FB43
FB04
FABC
FBC6
FEE1
02C3
052A
0554
04A7
04A1
051A
051E
04A2
0477
04E1
0542
0524
04DA
04D7
04F8
04DD
049F
049C
04CA
04DB
04F8
0572
05A3
040A
0049
FC42
FA48
FA9F
FB84
FB8A
FB01
FAE7
FB52
FB86
FB3B
FAED
FAF4
FB10
FB07
FB08
FB28
FB15
FACC
FAD6
FB52
FB66
FA92
FA16
FBE5
000E
0422
05BB
0511
0445
048A
0514
04ED
047A
048A
04EC
04F1
04B0
04CC
053E
054F
04D8
048D
04D9
052C
04F3
04B6
0520
055C
0395
FF96
FBB4
FA46
FB03
FBD2
FB9A
FB17
FB29
FB8A
FB88
FB33
FB1D
FB4C
FB44
FAEC
FAC2
FAEF
FB03
FAD8
FAE6
FB4A
FB4A
FAA4
FAA8
FCE8
00F8
0477
05A1
0506
046F
0494
04CA
048B
044D
0489
04E6
04E6
04BC
04D1
04FB
04E6
04C6
04FE
0548
0519
04AF
04E6
05A5
0549
0277
FE30
FB11
FA6B
FB0A
FB38
FADB
FADD
FB60
FBA7
FB72
FB49
FB70
FB70
FAFF
FA9F
FAD8
FB41
FB23
FAB5
FACF
FB57
FB37
FA68
FACB
FDE4
026F
0578
05B5
04AF
0473
052A
0598
052F
04AA
04A8
04CF
04A7
0470
0491
04D2
04DD
04E3
0522
053A
04CE
046C
04E4
05A6
04CB
0160
FD05
FA6B
FA61
FB3F
FB56
FACD
FAA0
FAE4
FAF6
FAC9
FAE8
FB5D
FB96
FB5F
FB36
FB68
FB82
FB25
FAD5
FB2F
FBAB
FB41
FA77
FB68
FF0D
0371
05BE
0578
0494
04B5
056C
058D
0509
04BE
04EF
0500
04A4
045E
0486
04B3
0493
048A
04DA
04FD
048D
043F
04DB
057A
0415
002D
FBF8
FA1E
FABF
FBAD
FB62
FA91
FA7D
FB09
FB43
FB09
FB00
FB52
FB83
FB64
FB5D
FB97
FBAB
FB62
FB35
FB77
FB90
FAEC
FA84
FC3C
0048
0452
05F5
0564
04A4
04D7
0553
053A
04C5
04A1
04D4
04E4
04BD
04B3
04C7
049E
044C
0454
04AC
04A5
0436
045A
0562
05B1
0368
FF07
FB48
FA23
FAD3
FB4C
FADB
FA71
FABF
FB39
FB46
FB33
FB66
FB83
FB2F
FAEB
FB4A
FBD7
FBBB
FB29
FB23
FBBA
FBC2
FACD
FA8C
FD01
018E
0532
05FA
050D
04A5
052E
0587
0530
04D8
04EF
04FA
049C
044F
0493
04FE
04DB
045E
0455
04C1
04D3
0472
0492
0557
0509
0222
FDB5
FA90
FA13
FAF2
FB45
FAC7
FA77
FAC1
FB0C
FAFC
FAFE
FB55
FB86
FB40
FB04
FB3F
FB83
FB4E
FB10
FB66
FBD5
FB62
FA7E
FB26
FE7E
02EF
05A7
05C1
04E8
04D8
0566
0588
052C
04FF
0518
04FB
04A0
048A
04CE
04E6
04A1
048A
04F3
0538
04BB
0424
0489
0559
0471
00E3
FCA3
FA68
FA97
FB54
FB32
FA9D
FA8A
FAEA
FB0F
FAE3
FAE7
FB30
FB48
FB1A
FB28
FB87
FB8F
FB0C
FAC9
FB4D
FBBF
FB38
FA9F
FC04
FFD8
03EC
05C3
0551
0490
04C5
054D
0535
04C6
04C7
051E
052B
04EA
04DC
0505
04EE
0493
0480
04DA
04FE
0496
0458
04EA
054F
03A4
FFBA
FBDA
FA46
FABC
FB4A
FAF7
FA85
FAC6
FB5D
FB7E
FB1F
FAD6
FAE0
FAF9
FAFE
FB20
FB4D
FB31
FAEA
FB0C
FB95
FBA4
FAF4
FAEA
FD21
0121
0487
059B
050C
04AD
0520
058A
0540
04BB
049F
04CA
04D6
04DD
0516
0535
04EE
049C
04C2
0518
04E8
045A
046C
0539
0518
0268
FE03
FABE
FA35
FB25
FB73
FACC
FA5E
FAB9
FB35
FB3E
FB23
FB4C
FB76
FB3F
FAEC
FB01
FB52
FB4A
FB05
FB2E
FBAB
FB7F
FAA4
FAE7
FDD4
0254
058A
0603
0506
0497
0511
056A
0524
04D5
04EC
04FC
04AA
0467
049D
04E9
04D6
04B8
0501
0546
04E2
0442
0478
054F
04D8
01B3
FD37
FA46
FA0E
FB05
FB52
FAF7
FAF3
FB53
FB5B
FAF3
FACE
FB2A
FB77
FB57
FB32
FB64
FB83
FB1E
FAB0
FAFC
FB9A
FB68
FAAC
FB6E
FEDC
0341
05CD
05C8
04ED
04D2
0533
0519
0495
047C
04F2
053C
04FF
04BF
04D4
04D5
047F
045B
04C5
051D
04D0
0476
04EB
0578
0435
0086
FC5A
FA31
FA5C
FB19
FB13
FAB8
FADF
FB4E
FB5E
FB29
FB2F
FB5A
FB3D
FAFF
FB20
FB7E
FB74
FAFF
FAEA
FB7F
FBC4
FAF7
FA54
FC07
0036
0448
05D6
054A
04B8
0502
0559
0519
04BC
04D3
0507
04D0
0475
0495
0509
0513
04A7
0487
04DF
04E5
0454
0431
0511
0584
0385
FF4B
FB7A
FA2E
FAD4
FB65
FB08
FA93
FAC5
FB34
FB48
FB3A
FB6D
FB9B
FB5F
FB08
FB0F
FB40
FB21
FAEC
FB3E
FBD4
FBA9
FAAF
FA9D
FD17
0157
04B1
058D
04EA
0495
04ED
052B
050A
04F6
0509
04E3
047F
0467
04C8
0510
04DC
04A5
04F7
0559
04F4
0436
0474
0599
0578
026E
FDDD
FACB
FA6D
FB40
FB70
FAF7
FAD8
FB39
FB58
FB05
FAEE
FB58
FB93
FB2C
FAC5
FB00
FB65
FB3A
FAD5
FB05
FB88
FB50
FA7C
FAEA
FDFF
0276
0574
05BD
04C6
047C
04FB
053A
04ED
04AE
04C4
04D1
04AE
04AF
04F4
0519
04E8
04C4
0501
0532
04DB
0479
04E4
0593
0498
0118
FCD6
FA6F
FA76
FB49
FB69
FAF8
FACD
FB02
FB1C
FB08
FB26
FB72
FB6F
FB0F
FAEA
FB38
FB62
FB0D
FACD
FB23
FB6C
FAE7
FA62
FBC2
FF89
03B5
05C5
0572
0491
048F
050C
051E
04D7
04D3
050F
050C
04CA
04B7
04D9
04CE
0491
0492
04E8
0508
04B5
04A1
0551
05B4
03F3
FFED
FBED
FA3B
FAAD
FB62
FB45
FADC
FAE7
FB3F
FB5B
FB34
FB20
FB21
FB01
FADE
FB0C
FB67
FB6A
FB1E
FB22
FB7D
FB51
FA61
FA34
FC81
00D1
0492
05D6
0534
0498
04DF
0555
053D
04DC
04C0
04D4
04C8
04B4
04D2
04F4
04E6
04E6
0528
0548
04D5
0451
04B2
05BC
0596
02C9
FE56
FAF1
FA1D
FAD8
FB5F
FB3F
FB13
FB19
FB04
FAD3
FADE
FB1C
FB1E
FADB
FADB
FB55
FBA5
FB40
FAB7
FAEE
FB8B
FB57
FA67
FABE
FDCF
0243
0543
05AE
04EC
04B2
0513
0526
04C8
04B0
051D
056A
052A
04CD
04CD
04EA
04C4
0497
04BB
04E3
04AA
047A
0501
05B2
04D5
018F
FD55
FA9C
FA44
FB02
FB4F
FB0D
FAE5
FAFC
FAFA
FAE4
FB08
FB4B
FB45
FB02
FB03
FB60
FB8B
FB37
FAF7
FB5C
FBD4
FB63
FA80
FB2A
FE7D
02EC
05BF
0603
0527
04D3
051D
052A
04C2
0480
04B8
04F9
04E0
04B7
04DD
050D
04D1
045C
0452
04C0
04F8
04A6
0470
0509
05CE
0513
0200
FDD2
FAD8
FA31
FAF2
FB7B
FB3D
FADC
FAF5
FB4E
FB5F
FB20
FB02
FB2C
FB44
FB10
FAE5
FB1F
FB76
FB5A
FAE5
FACF
FB46
FB83
FB04
FAD1
FC98
0075
044C
05E8
054E
0464
0476
0504
050B
04A5
04A3
0520
0566
051B
04CD
04F6
0534
04F5
047F
0495
052E
0558
04A8
040D
047A
052F
0441
00FA
FCF8
FA8F
FA6B
FB40
FB94
FB38
FAE5
FAF4
FB09
FAD2
FA8F
FA9C
FAEE
FB2E
FB39
FB31
FB33
FB28
FB0D
FB18
FB6A
FBA8
FB56
FAC0
FB2E
FDAE
019F
04EA
05F0
0520
0445
047F
053E
056B
04EF
04A0
04EE
054F
052F
04CA
04BA
0508
0537
0512
04E5
04D5
04A1
0441
0449
04FC
0541
0375
FF92
FBC5
FA3F
FAE0
FBAF
FB63
FAA2
FA9B
FB37
FB77
FB0F
FAC2
FB12
FB74
FB3F
FAC7
FACE
FB42
FB59
FAEA
FAC8
FB71
FC10
FBA1
FAC9
FB89
FECC
02EC
055A
055D
0483
046C
050C
0558
04FB
04A3
04CD
0514
04F4
04A2
04AD
0506
0511
04A6
0466
04BD
0523
04DA
0432
043D
0514
0524
02CD
FE9C
FB14
FA16
FB00
FBC1
FB5C
FAA6
FAAB
FB35
FB60
FB02
FAC9
FB12
FB60
FB39
FAEF
FB12
FB7E
FB91
FB41
FB2F
FB84
FB78
FAAA
FA56
FC46
0070
0479
0611
055C
0465
0482
0520
0529
04B7
04AA
052A
0574
0518
04A4
04B6
0509
04F6
0488
0468
04C2
04F4
04A0
046D
04FF
058F
045D
00D7
FCAD
FA40
FA3C
FB36
FB8E
FB16
FAB1
FAD4
FB16
FB04
FACF
FAE3
FB2C
FB47
FB2A
FB28
FB55
FB53
FAF3
FAAB
FAFF
FB9A
FB9E
FB0B
FB50
FDC3
01C7
050F
05FA
0529
047C
04D4
0577
0578
04FE
04C7
04EF
04EF
049E
047A
04CB
051D
04F4
049B
04A9
04FD
04ED
0471
0463
0515
0540
033B
FF45
FBAC
FA60
FAEB
FB63
FADF
FA36
FA64
FB21
FB7B
FB45
FB21
FB59
FB76
FB22
FAD3
FB0F
FB85
FB85
FB22
FB27
FBC2
FC02
FB37
FA6A
FB8C
FF16
031E
0548
0539
0494
04C2
0575
059D
0510
049C
04BE
0502
04E3
0499
04A2
04E5
04DA
047F
0471
04E2
0519
047F
03C5
041C
0546
0542
0291
FE46
FB18
FA7C
FB50
FBA4
FB07
FA83
FAC8
FB49
FB4C
FB00
FB00
FB46
FB4D
FB0F
FB1C
FB99
FBDD
FB6C
FADA
FB10
FBD8
FBFD
FB1D
FAAF
FC7E
005D
040D
0595
0522
0460
046B
04F1
0525
04EA
04B9
04D0
04F8
0503
050D
051E
04F4
0475
040B
0434
04BF
04F3
0494
0453
04CF
0550
042F
00CF
FCC2
FA68
FA7B
FB8B
FBDF
FB52
FAED
FB34
FB8E
FB5B
FAE3
FAC9
FB08
FB20
FB02
FB2C
FBB4
FBEE
FB78
FAF3
FB25
FBAB
FB73
FA9F
FAFA
FDEB
025A
0584
05F2
04DD
0454
04CD
052B
04BB
0421
0434
04C6
0512
04EB
04D3
0502
050F
04B8
046E
04AC
0517
04F5
0462
044C
04F5
0518
0324
FF4A
FBA4
FA1E
FA97
FB63
FB60
FAF3
FB01
FB91
FBE2
FB97
FB18
FAE4
FAEC
FAEC
FAF5
FB3A
FB86
FB62
FAE7
FACF
FB68
FBE7
FB77
FAC9
FBBB
FF14
0331
0594
058B
04A0
0479
0503
0527
049C
0434
047B
04F4
0502
04DA
04F8
052E
04E9
0454
0447
04F7
056E
04DF
0405
043A
0549
0522
024E
FDFC
FAE2
FA4F
FB19
FB7B
FB1E
FADE
FB2E
FB85
FB62
FB0A
FAFE
FB27
FB20
FAF7
FB1B
FB8B
FBB5
FB56
FAFD
FB46
FBD0
FBAA
FACE
FAA9
FCA8
006D
03F1
0581
0543
04A1
0492
04E6
0504
04D8
04BC
04D7
04F5
04EF
04E8
04F0
04D5
0479
0436
046D
04E4
04F3
0480
0453
04F6
0587
0453
00DD
FCD0
FA7B
FA78
FB5A
FB9C
FB2B
FAE9
FB23
FB53
FB1E
FAE4
FB0A
FB49
FB2C
FAE9
FB1C
FBB8
FBEF
FB5F
FAC9
FB04
FBA2
FB7E
FAA6
FADF
FDA2
01FC
0544
05EB
04F0
044E
04A5
0511
04E2
0493
04D0
0550
0550
04CC
048A
04E2
0538
04F0
0469
0468
04D9
04EE
0474
0449
04EF
0544
0382
FF99
FBBF
FA2D
FACF
FBB9
FB9B
FAF4
FAD2
FB35
FB4B
FAD7
FA89
FAD8
FB55
FB69
FB3A
FB48
FB82
FB63
FAF9
FAF9
FB98
FBEB
FB2F
FA59
FB70
FF0F
0345
0585
0553
0461
044C
04F5
0553
0516
04D5
04F3
051B
04FE
04D8
04EA
04EC
048D
042A
046D
052A
055C
0498
03DB
0450
0568
0516
022A
FDF7
FB07
FA79
FB34
FB97
FB44
FAEB
FAF4
FB0C
FAE9
FAD0
FB12
FB68
FB5E
FB13
FB1E
FB98
FBDD
FB78
FAEE
FB0B
FBA5
FBBB
FB01
FAC7
FCA7
0078
0423
05BE
0564
04AA
049E
04EF
04F3
04BD
04CD
051B
0521
04B8
0468
0494
04DF
04C0
0460
045F
04C7
04E8
047C
043E
04D3
0566
0436
00C0
FCBA
FA6B
FA60
FB34
FB7F
FB3B
FB1C
FB45
FB43
FB00
FAF4
FB4F
FB95
FB5F
FB0F
FB40
FBC5
FBD9
FB52
FAFD
FB67
FBD9
FB51
FA51
FACE
FDED
0252
055E
05E3
0508
048A
04C4
04F5
04C3
04B1
050E
054D
04E4
0445
044E
04F6
0543
04BB
041E
044A
04E1
04DE
043D
042E
0527
059C
038F
FF3D
FB4C
F9F5
FAC1
FB91
FB53
FAD0
FAF2
FB5F
FB3F
FAB4
FAA5
FB48
FBC3
FB7F
FB02
FB15
FB81
FB80
FB14
FB0E
FBA7
FBE8
FB24
FA78
FBDA
FF9C
03A4
05A4
0573
04BB
04AD
04F1
04CB
046E
048E
051F
055A
04EB
046F
0487
04ED
04F5
04A6
04A8
051C
054C
04C6
0435
047C
0527
0483
019E
FDAD
FAEF
FA5B
FAF6
FB5C
FB51
FB6F
FBD2
FBE2
FB55
FAC2
FACC
FB37
FB4B
FAF5
FAD9
FB3E
FB8C
FB30
FA9B
FAB3
FB65
FBA1
FB01
FAD8
FCCE
00B2
0455
05CF
0554
0487
0464
048F
0470
0434
045B
04D1
050E
04F5
04EA
0519
0524
04D3
0496
04E3
0560
0546
0499
045F
0525
05C9
046E
00BF
FC9E
FA50
FA49
FB24
FB83
FB5B
FB5F
FBB7
FBDF
FB8E
FB29
FB1C
FB39
FB1A
FACE
FAC4
FB0E
FB38
FB02
FAD6
FB1F
FB7A
FB25
FA6A
FADD
FDAB
01E3
0519
05DE
050A
046A
04A4
04FE
04D9
048F
04A3
04D2
0493
041E
043B
04FF
0583
052A
048E
0495
0513
051C
0498
0487
054F
0587
0369
FF44
FB95
FA5C
FB11
FBB6
FB5E
FACB
FAD5
FB3C
FB57
FB33
FB5D
FBCE
FBE5
FB73
FB17
FB49
FB92
FB45
FAAD
FAB3
FB70
FBD7
FB31
FA70
FB69
FEAC
02AA
053A
05A9
0506
04A6
04D5
050A
04DF
048E
047E
04B7
04DF
04BA
0470
0452
046F
0490
0497
04B1
0504
0554
053B
04CC
04A6
051A
055D
0411
00DB
FD1E
FACA
FA82
FB32
FB7E
FB22
FAD6
FB19
FB94
FBB0
FB60
FB0C
FAFB
FB11
FB24
FB37
FB53
FB5D
FB39
FB0A
FB1B
FB71
FB9E
FB2D
FA5A
FA3A
FBE2
FF4B
0302
053F
0571
04A8
0459
04D7
0544
04EC
0448
0448
0503
0591
0548
049A
0464
04B7
04E1
048F
0450
049F
0508
04D5
0448
0475
0598
062C
0469
006F
FC78
FA97
FAC6
FB65
FB53
FAE4
FAE3
FB54
FB8A
FB37
FAD3
FAE5
FB49
FB74
FB3A
FAFF
FB1F
FB6C
FB7D
FB44
FB28
FB65
FB97
FB2A
FA48
FA26
FC00
FFB0
037A
0576
054D
0458
0417
04BD
0556
052F
04A5
047A
04CE
0515
04F4
04B2
04B6
04E8
04E1
0496
046C
0497
04BF
048C
044E
04AC
058D
05BA
03F2
005D
FCB3
FAB7
FAAD
FB5E
FB8B
FB19
FAC3
FAF0
FB3F
FB30
FADF
FAD4
FB32
FB80
FB5A
FB10
FB30
FBA9
FBCF
FB5B
FAEB
FB2E
FBC1
FB96
FA8B
FA21
FC06
FFFE
03CF
0572
0502
0440
0471
0540
05A3
0548
04C6
04A6
04C1
04B2
047A
046E
04A1
04C1
0495
045F
0480
04E2
04FD
048F
041D
046B
055C
059C
03C7
0002
FC2D
FA3B
FA67
FB3A
FB52
FAC3
FA8E
FB19
FBAF
FB96
FB15
FAFA
FB6F
FBCC
FB95
FB2B
FB33
FB98
FBB1
FB48
FB04
FB69
FBF2
FBA7
FAA0
FA62
FC5C
002F
03D4
0587
0553
04A9
04A7
0524
0555
04FB
0496
049C
04D4
04C1
0462
0439
048C
04EF
04CF
044A
0412
0477
04E7
04BB
0437
0446
0516
0562
03A6
FFF4
FC36
FA61
FA9C
FB6D
FB7F
FAE6
FA8A
FAD6
FB4B
FB58
FB15
FB0B
FB60
FBA7
FB8A
FB46
FB52
FBAD
FBD9
FB94
FB40
FB5A
FBA6
FB65
FA8B
FA5B
FC4E
003C
0417
05CD
0547
0446
044A
051D
058B
051B
0488
0492
04FB
0502
048A
0432
0461
04B5
049E
043F
0436
04A9
04FF
04BD
045B
04AB
0589
0589
035F
FF79
FBDD
FA50
FABF
FB9B
FB9D
FAED
FA86
FAD7
FB56
FB61
FB1A
FB1C
FB91
FBF4
FBCE
FB61
FB41
FB7C
FB8C
FB30
FAE3
FB24
FB96
FB67
FA9D
FA97
FCB3
0093
0429
05AD
0540
0477
047E
051C
056D
0525
04BC
04A1
04AE
048C
044C
044A
049B
04E2
04D0
0497
049E
04E5
04F6
0494
043A
0494
0564
054C
0316
FF30
FB9F
FA2E
FABB
FB92
FB64
FA91
FA56
FB0E
FBCD
FBB0
FB09
FADA
FB66
FBE1
FB9A
FAF2
FAC4
FB31
FB86
FB5C
FB35
FB92
FBFE
FB96
FA93
FA9B
FD08
0124
049E
05CE
052D
046E
0490
0522
054B
04ED
0499
04B0
04F6
0504
04D0
04A7
04B5
04D0
04C3
049D
0497
04B6
04B6
0471
0438
0485
0524
04E8
02B2
FEDE
FB58
F9E8
FA81
FB7C
FB81
FAD6
FA97
FB18
FB93
FB5E
FAD9
FACB
FB37
FB6D
FB20
FADB
FB22
FBA5
FBAE
FB3F
FB1F
FBAF
FC30
FBB8
FAAF
FAC9
FD3E
0150
04CC
0613
056D
0479
046E
051C
0586
052E
048C
045F
04C8
0537
0533
04E8
04C8
04E5
04E9
04AE
047B
0483
0481
0435
03FB
0471
0549
0509
0280
FE6F
FB27
FA43
FB1F
FBD5
FB6F
FAA6
FA8A
FB12
FB63
FB13
FAA6
FAB3
FB1B
FB57
FB42
FB32
FB58
FB73
FB4D
FB2D
FB7B
FC0B
FC1D
FB50
FA6F
FAFD
FDB6
019A
04A7
05A0
050A
046D
04AA
054E
0570
04F5
049B
04E4
0562
0560
04DA
0477
0490
04BF
048D
043C
0461
04E9
050C
0475
03F1
046C
0566
0518
0266
FE5A
FB45
FA68
FAEF
FB41
FAD2
FA61
FA9D
FB38
FB6E
FB1D
FAD7
FB08
FB65
FB6C
FB22
FB08
FB53
FB98
FB6D
FB11
FB2D
FBD3
FC34
FB94
FA8A
FACC
FD73
0197
04F1
0601
0553
049B
04BF
0538
0529
04A7
047C
04F1
0561
0526
0483
044D
04C1
053E
052A
04C1
04A3
04DA
04C7
042F
03CB
0459
054D
04F0
0235
FE1F
FAF9
FA26
FAEC
FB8C
FB34
FA90
FA91
FB2B
FB8A
FB45
FADC
FAEE
FB52
FB5F
FAE8
FA8C
FAD6
FB78
FBB8
FB77
FB59
FBB4
FBEB
FB4E
FA79
FB23
FE3A
027B
0576
05F2
04F5
0453
04AB
0531
0524
04CA
04D1
0533
054C
04DD
0472
0498
050E
0521
04AE
0456
0493
0506
04F9
046A
0428
04B3
0545
0467
0180
FDB6
FAFE
FA5B
FB15
FBAE
FB66
FAC0
FA99
FB0A
FB6C
FB49
FAEC
FAE6
FB3D
FB70
FB3B
FAF6
FB11
FB65
FB74
FB37
FB30
FB95
FBC8
FB33
FA80
FB52
FE72
028F
0554
05B7
04CF
0453
04B8
052E
0512
04BE
04CD
0522
0521
04B1
0469
04AE
051B
0515
04B1
0497
04F9
053B
04CE
0419
0416
04F5
0590
046E
0157
FDA5
FB16
FA59
FAC5
FB39
FB2B
FAE1
FAD9
FB2D
FB80
FB7D
FB33
FAF4
FAF4
FB1E
FB4E
FB7B
FB9F
FB90
FB38
FADF
FAF5
FB68
FB88
FAF5
FA7C
FB9A
FED3
02C4
0548
058B
04AE
0452
04D6
0556
051B
0488
046B
04DE
0533
04F2
0472
045B
04BA
04FD
04C8
046E
0475
04D6
0505
04C5
048F
04E5
054F
0475
0191
FDA3
FAC3
FA25
FB04
FBA8
FB54
FAC1
FAD5
FB61
FB89
FB19
FAC7
FB1E
FBAC
FBAE
FB34
FB0A
FB84
FBFA
FBB4
FAFF
FABC
FB1B
FB4C
FAD0
FA81
FBCD
FEF3
0285
04CA
0552
04FF
04C7
04DA
04E7
04D3
04CD
04E9
04FA
04DE
04B3
04A5
04AA
0491
0455
0434
046A
04D3
0504
04C5
0476
04AC
0566
05A2
0426
00D3
FD1B
FAE0
FAB9
FB83
FBBA
FB0F
FA6D
FA9B
FB48
FB95
FB47
FAF5
FB1E
FB81
FB90
FB48
FB28
FB66
FB9A
FB67
FB16
FB36
FBAD
FBB4
FAFA
FA80
FBCD
FF2F
0316
0570
0593
04A1
0420
047C
0510
0538
050C
04F2
04F9
04E2
04A2
0485
04B1
04DC
04B5
046A
0473
04DA
050F
04A8
0418
043E
0527
0595
0420
00BF
FD0A
FACB
FA7B
FB1F
FB89
FB65
FB20
FB16
FB29
FB1E
FB05
FB17
FB4C
FB4F
FAFE
FAB5
FAE5
FB78
FBD4
FB9B
FB31
FB37
FB9E
FBA2
FAEA
FA6F
FBC0
FF39
034A
05C4
05E3
04CC
0420
0464
04F5
0528
0500
04DC
04D7
04C7
04A7
04A3
04CD
04F4
04F2
04E5
04F4
04F6
04A7
042A
0410
04B8
05A0
0593
03A8
002E
FC99
FA79
FA53
FB52
FC18
FBE9
FB25
FAA0
FAB2
FB01
FB24
FB20
FB28
FB2B
FAFA
FABA
FAD9
FB65
FBCA
FB94
FB28
FB4E
FBF3
FC11
FB25
FA5B
FB8C
FF19
0334
059E
05C6
04EE
0477
049A
04D0
04D9
04E9
0514
0524
04FA
04C9
04CA
04F4
0512
050A
04E7
04B5
048B
048F
04C4
04DC
0499
0455
04B6
0597
05A1
038C
FFBA
FC2B
FA91
FACB
FB6E
FB79
FB1C
FAE9
FAF5
FAFD
FAF1
FAEF
FAEB
FAC2
FA9C
FAC6
FB33
FB6F
FB45
FB16
FB44
FB8F
FB75
FB13
FB08
FB62
FB58
FA95
FA47
FC0D
FFE0
03B5
058A
0566
04D8
04EB
0549
0548
0507
0509
0541
0536
04DA
04AA
04E9
0538
0527
04CB
048A
0484
0499
04CA
0521
054D
04EA
0453
047F
0586
05DD
03C3
FF89
FB9B
FA0A
FA85
FB28
FAE8
FA6A
FA9D
FB49
FB91
FB33
FAB8
FA96
FABF
FB05
FB56
FB8A
FB59
FAD5
FA8E
FAE6
FB75
FB8A
FB2D
FB06
FB2C
FAEA
FA26
FA4E
FCEC
016B
052C
062E
051D
042F
0484
054A
0569
0500
04DF
052F
0563
0530
04E2
04C4
04C3
04C1
04DA
050F
0514
04C4
0485
04C2
0524
04FC
0479
0495
056E
056A
02E9
FE95
FB12
FA2F
FB16
FBAC
FB2B
FA8B
FAAA
FB14
FAFB
FA88
FA7F
FAFB
FB58
FB3D
FB10
FB33
FB70
FB68
FB30
FB17
FB0C
FAD8
FABA
FB2E
FBE6
FBE1
FB00
FAD8
FD14
0134
04B8
05CC
0515
0484
04E9
0572
0549
04C2
04A5
04FA
0533
0517
04EF
04E1
04CC
04AD
04B7
04E4
04DF
049B
0494
0512
0577
0504
0427
0422
0510
0519
0282
FE22
FACA
FA31
FB45
FBD8
FB43
FAA1
FAD2
FB53
FB4A
FADB
FAC5
FB2D
FB81
FB6C
FB34
FB20
FB19
FAFC
FAF6
FB29
FB53
FB34
FB13
FB55
FBAA
FB5E
FABC
FB4D
FE17
01FF
04B8
0543
04BD
04AF
0534
0560
04EB
0491
04CE
051A
04CF
0432
0404
0463
04C9
04EB
0502
0526
050A
049C
045D
04AA
050B
04D0
044C
0481
055D
0523
0265
FE16
FAD4
FA1F
FB00
FB98
FB4E
FAE3
FAEC
FB1C
FB0E
FAFD
FB3B
FB85
FB6C
FB16
FB03
FB49
FB81
FB74
FB60
FB6B
FB53
FAFC
FAD6
FB3C
FBA7
FB4C
FAA6
FB6F
FE93
02AF
0550
0590
04B8
0460
04BA
04F8
04C8
049E
04BF
04D9
04B8
04B8
0514
0552
04EF
0442
0417
0492
0506
0501
04D4
04DA
04CF
0466
0426
04BA
0574
047C
010E
FCE7
FA98
FAB7
FB90
FB83
FAC7
FA8F
FB20
FBA0
FB7F
FB2E
FB37
FB68
FB4F
FB0C
FB09
FB33
FB27
FAE8
FAE4
FB32
FB5E
FB32
FB24
FB8C
FBD5
FB4C
FA9F
FB9A
FEEC
02EB
0539
054B
0496
047B
04DF
0507
04E6
04F9
053F
0526
0499
0444
0493
050B
0513
04E5
050F
056D
0556
04BC
045C
049C
04EE
04C4
0493
050E
0585
0434
0091
FC7F
FA6F
FABB
FBA5
FBAE
FB09
FAAE
FAD7
FB10
FB2E
FB70
FBB7
FB7B
FAB8
FA3E
FA9B
FB44
FB60
FB09
FAF9
FB55
FB7A
FB22
FAE8
FB33
FB5E
FABE
FA38
FBB3
FF96
03C2
05C6
0581
04C8
04DF
0549
0517
0479
0448
04AF
0506
04F2
04D4
04F7
0506
04BF
048C
04D3
0531
050C
049B
049F
051E
053C
04A4
044D
0505
05B0
0424
0009
FBCB
FA09
FAB6
FBA5
FB6A
FAAB
FA9B
FB33
FB8C
FB53
FB14
FB2A
FB44
FB1C
FAFA
FB23
FB4D
FB2C
FB0A
FB48
FB95
FB57
FAC4
FABB
FB62
FBB0
FAFC
FA7E
FC36
003B
0430
05CB
0542
047E
048C
04D9
04B6
047B
04BD
0530
0517
0484
044A
04BC
052E
050A
04AD
04B0
04EB
04DA
0494
04A0
04F2
04E4
0469
0466
0541
0598
038A
FF49
FB6B
FA2E
FB18
FBF8
FBA8
FAEC
FACB
FB26
FB48
FB1D
FB20
FB67
FB7E
FB40
FB1B
FB4C
FB6E
FB36
FB06
FB48
FB9A
FB5D
FAD2
FADB
FB87
FBBD
FAEB
FA6C
FC3D
0058
0448
05D9
055B
04BB
04EA
0531
04CB
0424
0416
049E
0503
04F6
04D9
04F5
0506
04D6
04AD
04CB
04E8
04B8
0482
04B2
0504
04DA
045E
047C
055E
0582
0340
FF0E
FB6C
FA38
FAD6
FB6A
FB36
FAF8
FB49
FBB2
FB94
FB24
FB05
FB3B
FB3E
FAEB
FAC1
FB09
FB60
FB65
FB51
FB71
FB7D
FB1F
FABB
FB00
FBAE
FBAD
FAC6
FA9E
FCFF
015C
04FC
05E2
04DC
041C
0486
052D
0520
04AD
049D
04F4
051F
04F2
04D1
04ED
04F4
04BB
0494
04B9
04DA
04A8
046F
0497
04DE
04B7
0457
0496
056D
0548
02AE
FE60
FAF6
FA22
FB05
FBA9
FB5D
FAF2
FB0D
FB48
FB1B
FAC6
FAD6
FB39
FB65
FB40
FB42
FB90
FBB0
FB55
FAEC
FAF4
FB39
FB40
FB26
FB5F
FBB5
FB71
FAB6
FB08
FDAB
01C1
04E1
05AF
0523
04E4
053A
0545
04B3
043B
046E
04DB
04DE
0499
04A1
04F6
0501
049D
045F
04A5
0500
04EF
04B2
04BD
04DC
0497
0436
0489
055A
04FF
0232
FDFE
FAF3
FA57
FAF9
FB10
FA77
FA4C
FB01
FBCB
FBE8
FB95
FB70
FB83
FB72
FB42
FB42
FB57
FB16
FA9D
FAA0
FB48
FBBB
FB54
FAB6
FAED
FBBC
FBDF
FB1E
FB2D
FDAF
01DA
0510
05CC
0518
04C5
0528
0552
04DC
0470
0493
04E5
04D8
0490
0488
04BF
04CB
04A9
04C2
0521
0540
04E7
049D
04C6
04F3
04A8
0462
04ED
05B6
04D7
015D
FCE7
FA32
FA29
FB3B
FB9D
FB45
FB2B
FB81
FB9A
FB34
FAE2
FB0E
FB52
FB36
FAFA
FB1D
FB76
FB6F
FB06
FADA
FB1F
FB40
FAF6
FAE2
FB79
FBEA
FB34
FA19
FADE
FE8B
0334
05DB
05BA
04B6
04AD
055A
0572
04C8
045A
04A1
04FC
04D5
0484
049A
04EA
04E2
048A
047A
04DB
0524
0502
04D7
04EF
04E3
0461
0408
0499
056C
04A9
017C
FD68
FAD6
FA83
FB1B
FB34
FAD8
FAC7
FB14
FB34
FB02
FAE6
FB11
FB3B
FB3E
FB5F
FBC0
FBEF
FB86
FAEA
FAD5
FB41
FB72
FB31
FB2C
FBBB
FBFF
FB2A
FA36
FB44
FF02
0371
05E1
05BB
04AE
0458
04B2
04E6
04C5
04BD
04DF
04D0
048B
0480
04D1
0507
04C7
046C
0477
04C1
04BC
046A
0462
04C6
04F5
049F
047E
052F
05C0
0458
008D
FC57
FA25
FA58
FB3E
FB58
FAD0
FAA5
FB15
FB87
FB91
FB6B
FB62
FB6E
FB73
FB7D
FB8A
FB73
FB33
FB1B
FB60
FBA3
FB67
FAE2
FAD5
FB5D
FB95
FAF4
FA8D
FC23
FFE6
03D3
05B1
054E
0458
043E
04DE
054F
0542
0512
04F7
04C3
0469
0437
045F
049F
049F
0469
0455
0493
04F9
0543
054B
04FF
047C
0437
04A2
0568
0548
033B
FFBB
FC7F
FAE4
FACD
FB33
FB61
FB67
FB71
FB5D
FB0D
FAC1
FAC9
FB0C
FB34
FB32
FB48
FB8B
FBBC
FBAC
FB7C
FB59
FB30
FAF7
FB02
FB97
FC3C
FBFE
FADC
FA5F
FC31
0013
03CD
0567
0507
045E
048D
052E
055D
0506
04C6
04E3
0502
04DB
04A7
04B8
04E6
04CD
046F
043E
047D
04DC
04E8
04A9
0481
0494
049C
046B
0453
04BA
0550
0500
02E8
FF6E
FC28
FA88
FAA8
FB60
FB91
FB21
FAC3
FAEF
FB5A
FB79
FB3C
FB0E
FB2B
FB58
FB51
FB33
FB48
FB80
FB80
FB32
FAFA
FB2E
FB97
FBB9
FB89
FB6D
FB85
FB64
FAE0
FAD4
FC7B
FFE3
0375
055D
0553
04A7
0493
050A
053F
04F0
04A2
04C0
0503
04F9
04B4
04A2
04CD
04C8
0461
0408
0436
04B2
04D7
047F
0440
048E
0500
04E6
0462
045D
0524
057E
03C4
FFED
FC04
FA40
FAD9
FC04
FC0E
FB04
FA34
FA6C
FB34
FBA1
FB78
FB2A
FB0F
FB13
FB19
FB43
FBA0
FBE4
FBB5
FB3B
FAFF
FB32
FB6A
FB40
FAF8
FB21
FBA6
FBC2
FB2B
FAEC
FC80
0003
03B9
05A5
0576
0490
0456
04CD
0513
04BD
044F
0460
04CF
0506
04CC
0477
045B
0461
0457
045C
04B1
0531
055E
0505
0497
048F
04C4
04A1
041D
03F5
0490
0502
03B5
004A
FC6C
FA50
FA83
FB90
FBD0
FB21
FA90
FAC4
FB50
FB83
FB5C
FB51
FB80
FB96
FB72
FB69
FBAD
FBDA
FB76
FABE
FA7A
FAF3
FB8C
FB91
FB36
FB3D
FBC6
FC07
FB76
FAF1
FC10
FF45
0312
0563
0592
04C3
0469
04D0
0546
053E
04E8
04B2
04A8
048F
0462
045A
048A
04B4
04A5
0487
049D
04D5
04D9
0499
0473
04B1
0507
04EA
0460
0422
04A8
0531
0442
013D
FD5C
FAAE
FA2B
FAF2
FB77
FB2C
FAC1
FAF0
FB89
FBD4
FB94
FB37
FB22
FB38
FB3D
FB45
FB77
FB9A
FB4D
FAB9
FA92
FB28
FBD2
FBB5
FAF8
FA9D
FB13
FB85
FB17
FA78
FB71
FEBF
02DE
0572
05A0
04A4
041D
0464
04BB
04A6
0474
0492
04E0
04F4
04BF
0492
0498
04AA
04A0
04A3
04E4
0533
052A
04BC
0460
0482
04F6
0530
0504
04E4
052E
0560
0456
018A
FDEA
FB3A
FA81
FB34
FBF8
FC01
FB8E
FB38
FB25
FB19
FAFB
FAFB
FB24
FB3A
FB12
FAF2
FB2F
FB9D
FBAF
FB3E
FAD8
FB05
FB76
FB6F
FAE0
FA98
FB13
FB98
FB20
FA19
FA78
FD89
020F
0541
05A7
047B
03E7
048E
0550
0528
047F
0458
04DF
0559
054B
04FD
04D1
04A4
043B
03E5
041D
04BB
050B
04C5
047B
04C3
0549
0544
04AD
0479
0542
061A
0545
022A
FE26
FB55
FAA1
FB39
FBB4
FB77
FAF3
FABE
FADD
FAF0
FAD6
FADA
FB38
FBB3
FBE4
FBC3
FBAE
FBCF
FBD0
FB5E
FACE
FACB
FB5B
FBB5
FB52
FAB6
FAB3
FB2A
FB30
FAA7
FAFA
FD90
01B6
04F2
05A6
04B4
0426
04B7
0567
054A
04CC
04CF
0537
0526
0469
03D9
0422
04C6
04E0
0473
044E
04BD
0518
04D4
0464
048E
052C
0547
048F
040C
04C1
05FA
05A2
0293
FE19
FACE
FA0F
FAF0
FB9C
FB50
FAC0
FAC7
FB4F
FBA0
FB73
FB33
FB4D
FB96
FB9B
FB55
FB2D
FB57
FB81
FB53
FAFF
FB00
FB57
FB79
FB1F
FAC5
FAFD
FB7B
FB60
FAA8
FAC1
FD13
0124
04AE
05E9
0543
048C
04BD
0537
0514
0486
0463
04C8
04F6
048D
042D
0482
052A
0530
0476
03F5
0461
0524
053E
04B4
047F
0509
0582
0529
0491
04DC
05D8
05B2
0306
FEBD
FB49
FA25
FA98
FB01
FAC9
FA9A
FB07
FBAB
FBCB
FB52
FAD4
FAC5
FB02
FB2B
FB37
FB59
FB93
FB96
FB3C
FADF
FAF3
FB69
FBB1
FB6D
FAF7
FADD
FB0D
FAE2
FA43
FA58
FC81
0087
045F
060F
0597
04A3
0481
04F9
052D
04F6
04E8
0532
054A
04DD
046A
048F
0508
0511
048D
0441
04B3
0557
0554
04BB
046D
04CB
0523
04CB
0445
049A
05A7
05BF
0371
FF5B
FBBD
FA46
FAA7
FB54
FB56
FAF3
FAD3
FB04
FB1C
FAF4
FAD7
FAFC
FB2E
FB22
FAF4
FB07
FB71
FBCC
FBB9
FB60
FB2C
FB31
FB17
FABF
FA94
FAF2
FB75
FB4F
FA85
FA66
FC5C
002E
03E6
05A7
0568
04AC
04AE
053E
0571
0505
0490
0494
04D9
04EF
04DD
04F9
0536
0523
049E
042A
044F
04CD
04FB
04BA
049E
04FC
0551
0504
0471
0490
056C
0595
0395
FFC5
FC31
FA90
FABA
FB4C
FB5D
FB1C
FB04
FB17
FB12
FAFD
FB17
FB58
FB64
FB18
FAD3
FAFD
FB73
FBAD
FB70
FB17
FB0F
FB4A
FB5B
FB1F
FAF8
FB41
FBB0
FB98
FAF6
FAEF
FCD1
007F
042C
05EE
0596
04A3
0476
04F1
050C
0476
03F9
0447
04FF
0543
04EC
049E
04C5
0504
04E6
049C
049F
04DF
04D5
046D
0444
04B6
052B
04E2
042F
042E
0514
056E
039E
FFD5
FC19
FA2C
F9F9
FA40
FA51
FA85
FB38
FBF9
FC14
FB8F
FB15
FB19
FB57
FB5E
FB39
FB3F
FB76
FB86
FB46
FB0C
FB34
FB90
FB99
FB3A
FB04
FB77
FC2A
FC20
FB24
FA77
FBC4
FF46
0346
05A6
05DF
0530
04FF
055F
057A
0502
049C
04D4
0543
0522
0474
040E
0464
04EC
04E9
047F
046D
04E2
0535
04F1
048C
04A5
04F4
04B1
03EE
03CB
04C9
0592
0426
0055
FC4F
FA66
FAB7
FB83
FB77
FAE7
FAC4
FB24
FB5C
FB27
FB03
FB4B
FB9E
FB70
FAF2
FACB
FB24
FB6B
FB2D
FACA
FAE6
FB71
FBAE
FB42
FAC9
FB04
FBB0
FBB8
FAC5
FA23
FB9E
FF6F
03AF
0616
061C
0527
04BF
0508
0521
049F
0417
042C
04A5
04D0
0489
0462
04BE
0535
0530
04CF
04B5
0510
0548
04E7
0457
0450
04BE
04DF
047B
0465
053D
0609
04E1
0137
FCDF
FA57
FA3F
FB10
FB30
FAAC
FA89
FB12
FB7E
FB3F
FAD8
FB09
FBA8
FBE6
FB80
FB17
FB2C
FB60
FB1F
FAA6
FAC0
FB80
FBF5
FB70
FA9B
FAAB
FBA6
FC37
FB7E
FA8A
FB69
FEC0
02D8
054F
056C
047D
041D
04A1
053D
0551
050C
04EF
0512
0531
0522
0504
04F1
04CC
0483
0451
047C
04E0
0502
04B4
0460
0481
04ED
0506
04AB
0484
0511
058D
0465
0108
FCED
FA56
FA29
FB38
FBCE
FB71
FAED
FAEE
FB34
FB2F
FAE8
FAD7
FB10
FB22
FAD6
FA9A
FAE4
FB6F
FB8C
FB1D
FAD3
FB29
FBA8
FB8B
FAEE
FAC0
FB62
FBED
FB6B
FA83
FB25
FE4B
028E
057B
0609
0551
04E2
0513
053A
0505
04E3
052A
0578
054A
04C3
0472
0488
04BA
04CC
04DB
0502
050C
04CD
0489
04AB
051E
054F
04F4
0487
04AB
0543
055D
0412
0152
FDFB
FB41
F9F2
F9FC
FA96
FAF8
FAF6
FAED
FB1E
FB51
FB30
FAD2
FA9D
FAAD
FAC1
FABE
FAE7
FB50
FB95
FB64
FB11
FB2C
FB9D
FBB2
FB39
FAED
FB60
FBE1
FB4E
FA06
FA19
FCF9
0184
050C
062C
05D1
0598
05DA
05DE
0559
04DC
04D9
04F7
04BD
046B
0495
052C
0582
053B
04BA
0487
04A9
04D3
04F1
0524
0557
0533
04AF
043D
044A
04BE
0538
0586
058D
04DB
02DB
FFAB
FC6D
FA6C
F9F8
FA52
FAA3
FABD
FAE1
FB1D
FB49
FB55
FB5C
FB63
FB43
FAFC
FAC7
FAD3
FB05
FB2A
FB43
FB60
FB58
FAF7
FA7F
FA7C
FAFF
FB68
FB3F
FAF1
FB2A
FBAD
FB90
FAD7
FB18
FDC8
0219
0573
063B
055F
04C3
04ED
04FF
0491
045E
04F9
05B6
0591
04B1
0433
048D
04FE
04D1
0461
0467
04D6
0517
0509
0508
0520
04ED
046A
042D
0489
04F7
04DA
048E
04C9
0509
03B1
002F
FC3F
FA30
FA61
FB41
FB72
FB1F
FB0A
FB43
FB4E
FB1C
FB13
FB3C
FB22
FAB8
FA8F
FAE9
FB32
FAE8
FA79
FA9C
FB25
FB55
FB13
FB17
FBAB
FC15
FBB6
FB22
FB43
FBC2
FB6B
FA62
FABB
FDF2
0297
0598
05B3
048B
043E
04EA
053C
04AC
0426
0476
0522
054A
04FB
04F0
0566
05E1
05FD
05D3
058E
0527
04B4
0494
04E7
052B
04D1
041C
03D9
0440
04A2
0483
0464
04D2
0516
03AE
0047
FC89
FA7D
FA7C
FB32
FB6B
FB3A
FB32
FB4D
FB28
FAD0
FABC
FAFB
FB0D
FAA8
FA38
FA38
FA80
FA90
FA65
FA72
FAD5
FB22
FB28
FB47
FBB4
FBF0
FB88
FB01
FB2C
FBC8
FBA8
FAAD
FAAC
FD6C
01FF
0556
05B2
0484
0437
0529
05C9
053C
047B
04B0
0584
05CF
055A
04FF
0538
0585
0570
054D
0572
057D
050A
0484
048E
04F1
04F1
048C
047E
04FA
052F
04A1
0431
04D8
05A5
0461
0086
FC60
FA72
FAA9
FB0D
FAA5
FA44
FAB1
FB4E
FB31
FAA6
FAA5
FB31
FB47
FA88
F9E1
FA25
FAE2
FB35
FB18
FB11
FB14
FAB9
FA44
FA7F
FB60
FBCB
FB23
FA57
FA9C
FB74
FB50
FA2F
FA54
FD80
0256
05AD
061E
052A
04DF
0578
05D1
055D
04C2
04A5
04D9
04EF
04F6
052E
056D
055D
0519
04FD
050D
0502
04E5
050F
057C
05A3
053D
04D9
0519
05AB
05A4
04F8
04BD
0580
05EF
0411
FFD8
FB9E
F9BF
FA37
FB21
FB21
FA96
FA6C
FAAA
FAB3
FA71
FA74
FAFA
FB7C
FB73
FB15
FAF4
FB25
FB3E
FB15
FAF0
FAF7
FAF3
FAC5
FAAF
FACF
FAC7
FA5F
FA1F
FAA8
FB7D
FB6B
FA6B
FA67
FD2E
01DA
0565
0600
04F4
049E
057C
062A
05C0
04F8
04D9
053C
0551
04FC
04D4
0501
04FC
0492
0457
04A9
0503
04DB
048A
04AF
051D
0537
0511
054D
05DD
05D4
04E7
0450
0523
0637
04FF
00D4
FC32
F9F2
FA30
FAE3
FAC9
FA80
FAD9
FB6A
FB5F
FAD8
FAA4
FAF0
FB19
FAD1
FA98
FAD1
FB1C
FB1B
FB26
FB9F
FC10
FBC9
FB0D
FAC3
FB13
FB2C
FAA3
FA3A
FAB0
FB57
FAEE
F9D1
FA3A
FD8E
024C
0579
05DC
04DD
0467
04D2
0535
04FD
048B
0469
049B
04D9
050F
054B
056F
054D
04FF
04C4
04A6
048A
0475
048B
04B7
04B2
047B
047C
04F4
057C
0574
04EF
04C1
054D
0592
0401
0062
FC7B
FA6C
FA98
FB80
FBA7
FB12
FAC1
FB27
FBAB
FB9D
FB19
FABB
FAC4
FAF2
FB0D
FB2A
FB58
FB70
FB5D
FB49
FB49
FB37
FB08
FB06
FB52
FB81
FB23
FA87
FA73
FAFC
FB3B
FAC6
FAD7
FD1A
013B
04BF
05B9
04DD
043C
049F
0515
04DA
0483
04E0
0593
059B
04D8
043B
045E
04C3
04CD
04AF
04D9
0520
0513
04D0
04C5
04F0
04F2
04D9
051E
05B1
05CA
0516
0483
0506
05C7
04A5
00F0
FCB1
FA82
FABC
FB93
FB92
FAF5
FAA3
FAD0
FB10
FB2F
FB52
FB6E
FB46
FAF4
FAE8
FB2D
FB39
FACE
FA7A
FAC5
FB51
FB61
FAFD
FAD7
FB22
FB36
FAA8
FA15
FA55
FB1D
FB48
FAA3
FAA7
FCDC
00CB
0442
059E
0544
04BC
04E0
054B
0552
04F4
04AD
04B6
04C5
04A5
0498
04F9
059F
05ED
0589
04CE
046E
04B6
0548
0589
053F
04C1
048F
04CA
0514
0507
04C4
04E1
0599
0606
04A2
00F2
FC90
F9F4
FA06
FB56
FBE2
FB3E
FA83
FA95
FB1D
FB58
FB32
FB1C
FB2D
FB10
FABD
FAA0
FADA
FAFC
FAC4
FA97
FAD5
FB2B
FB18
FACD
FADF
FB45
FB50
FACD
FA73
FAC9
FB36
FB06
FB10
FD1C
014A
052D
065C
0534
0421
0487
0589
05C5
053F
04F6
0535
0556
04FB
04AA
04E7
0563
058B
055E
0539
0522
04E7
04A7
04A8
04D5
04E1
04E4
0536
05A9
0584
04A2
0415
04C8
05BF
04AE
00D0
FC45
F9E7
FA42
FB68
FB86
FAAF
FA0A
FA17
FA68
FA97
FAB9
FAE5
FAE3
FAA2
FA7B
FAAE
FAF5
FAF8
FAF1
FB48
FBCF
FBE3
FB5D
FADF
FAEB
FB2E
FB0F
FAB0
FABD
FB40
FB67
FADB
FAC9
FCC8
00B8
047E
061B
05AB
04E3
04F6
058D
05C2
057C
0557
059A
05DF
05C1
0565
0527
050F
04E5
04A9
0499
04C8
04F1
04D9
049D
047D
0493
04D2
0526
055B
052C
04A9
0475
0501
058F
047B
010F
FCD0
FA40
FA43
FB4F
FB73
FA88
F9E2
FA41
FAF4
FB0B
FAA1
FA7D
FADC
FB35
FB20
FADE
FACA
FAD4
FAD1
FADE
FB18
FB45
FB2C
FB0A
FB31
FB6D
FB46
FAD5
FAC6
FB41
FB81
FB0B
FAFC
FD10
0130
04F8
063C
0563
0489
04D0
057B
0586
0518
04ED
0510
04F8
04A4
04B5
0559
05D7
059A
050B
04DD
0500
04EC
049E
048A
04C8
04EB
04CF
04D9
0534
0554
04D6
0462
04D4
057D
0461
00BA
FC65
FA00
FA0D
FAD8
FAE3
FA79
FA9A
FB47
FB9E
FB42
FACA
FAC3
FAF8
FAFE
FAE2
FAE3
FAEB
FAD8
FAE8
FB57
FBCC
FBB8
FB36
FAF8
FB3D
FB67
FAFC
FA7F
FAC1
FB81
FB9D
FAE6
FAE9
FD2F
0124
047C
05A9
0541
04D7
0519
0584
057E
0528
04F1
04E7
04D1
04AE
04B7
04F0
0508
04D4
048E
0492
04E7
0533
0524
04C3
046F
0480
04ED
0543
0506
043E
0399
03D8
04E8
058B
0449
00F0
FD0C
FAA7
FA71
FB4A
FBA8
FB25
FA8C
FA95
FB09
FB37
FAFB
FAD4
FB1B
FB83
FB91
FB49
FB18
FB47
FBA7
FBD1
FB93
FB25
FAFF
FB5C
FBD8
FBD1
FB38
FAD0
FB3D
FC05
FBFD
FB07
FAD4
FD25
016D
0502
0603
052F
048F
04E2
0549
050D
04A7
04C4
051A
04EF
045F
043E
04C5
0528
04D2
0439
0415
0446
0441
040C
0428
0496
04C3
0473
0428
044D
0491
0477
0449
049F
050F
0425
012D
FD67
FAD5
FA30
FA94
FAE5
FAD9
FAB9
FAC0
FAF3
FB45
FB90
FBA0
FB73
FB5A
FB8C
FBBF
FB86
FB11
FB0E
FBA1
FC14
FBE8
FB9A
FBDB
FC6B
FC67
FBB0
FB30
FB84
FC05
FBB1
FAD0
FAFE
FD53
00FD
0409
0552
053B
04D1
04BB
04ED
0511
04F2
04B3
0498
04B2
04CE
04C2
04AC
04B3
04B9
047E
0419
03FC
0461
04E0
04DC
045A
03FC
0424
047F
049B
0487
048A
048A
0448
03FF
043B
04E5
04ED
0344
0025
FD08
FB41
FAE3
FB0B
FB06
FAE0
FAF7
FB5E
FBC1
FBBE
FB4F
FADE
FAD7
FB29
FB64
FB57
FB40
FB5A
FB7D
FB70
FB51
FB68
FBA3
FBA3
FB54
FB2C
FB73
FBB4
FB5B
FAC6
FAE0
FBAF
FBFF
FB25
FA65
FBBA
FF5A
033B
053C
053D
04B4
04AE
04E9
04C9
046A
0459
04A7
04E7
04D9
04AB
049D
04B5
04D1
04CB
0499
0460
045C
0499
04D4
04D4
04B7
04C9
050B
0526
04F7
04D1
04F4
0505
048D
03E8
03FC
04B4
0481
020E
FE20
FB0B
FA4B
FB2A
FBE7
FBA4
FAEF
FAA1
FADF
FB36
FB52
FB3A
FB17
FB11
FB39
FB70
FB77
FB44
FB15
FB16
FB23
FB12
FAFB
FAFE
FB00
FADB
FABA
FAE3
FB3F
FB6A
FB4F
FB5C
FBBE
FBEA
FB69
FB18
FC99
0038
040E
05E2
0586
04A3
048A
04F7
050F
04C7
04B9
050B
0530
04D2
0463
0478
04F5
0546
0535
050D
050B
0517
0508
04E6
04DB
04FC
0526
050F
049F
0432
0440
04B8
04F9
04A5
044C
04B7
056E
04A3
0139
FC9A
F9B7
F9E3
FB79
FC07
FB1B
FA36
FA70
FB37
FB75
FB13
FACE
FAF0
FAFD
FAA3
FA46
FA66
FAD3
FB04
FAE9
FAE8
FB34
FB80
FB7E
FB41
FB16
FB22
FB44
FB4F
FB4D
FB6C
FBA0
FB89
FAE9
FA56
FB10
FDD9
01D9
050C
0613
0576
04DC
051A
0591
0578
050B
0505
0571
059D
0533
04B4
04B9
0526
056B
054F
051E
0512
0503
04C6
0493
04B1
04F7
04F6
0494
0440
0467
04F3
0556
052A
04A9
0479
04BC
0487
02A7
FF24
FBAE
FA19
FA83
FB57
FB36
FA6F
FA38
FAD3
FB42
FACD
FA10
FA0C
FAB4
FB24
FAFA
FAC5
FB0A
FB73
FB67
FAFA
FAD3
FB30
FB8B
FB63
FAFA
FAE8
FB3F
FB82
FB6D
FB54
FB8E
FBDC
FBAB
FAF2
FAAC
FC1B
FF78
035A
05C9
0600
0505
0474
04DF
0585
0590
0521
04F1
053A
0579
054F
0504
04FF
0520
0506
04B8
0499
04BC
04CC
04A1
0494
04EF
0553
051F
046C
0417
049F
054F
051B
0415
0381
0431
0530
048F
0185
FD7B
FAC7
FA69
FB42
FB99
FAF7
FA4F
FA7F
FB2E
FB6C
FAFF
FA95
FAC3
FB38
FB48
FAEE
FAC9
FB20
FB79
FB50
FADC
FAB9
FB08
FB55
FB52
FB3B
FB5D
FB86
FB5B
FB00
FB07
FB92
FBED
FB76
FAB4
FB25
FDAC
0172
0486
059D
0518
0464
0470
04FB
0545
0514
04D7
04E8
0511
04F8
04B2
04A5
04EB
0526
0514
04EF
050A
053A
050E
049A
0482
0506
057C
0521
0441
03EF
0495
054B
050D
0435
040D
04E5
0540
0364
FF86
FBCD
FA26
FA7F
FB4C
FB68
FB09
FAF6
FB56
FB9A
FB5A
FAE0
FAB4
FAED
FB2C
FB2B
FB0B
FB07
FB14
FAF9
FAB9
FAA1
FADF
FB30
FB39
FB08
FB05
FB4D
FB79
FB3A
FAE5
FB16
FBBB
FBFD
FB67
FAE3
FC0D
FF57
0339
058E
05A1
04A4
042B
0494
051E
0527
04E0
04CC
04F6
0503
04D6
04C0
04FB
0540
0529
04C5
048D
04BA
04FA
04EC
04AE
04AC
04F3
050A
04AA
0442
046E
050E
054A
04B8
0413
0452
0520
04D1
0231
FE2C
FB17
FA5B
FB27
FBA3
FB10
FA48
FA51
FB04
FB71
FB32
FAD3
FAEB
FB4F
FB6E
FB2D
FB01
FB2F
FB69
FB54
FB20
FB3D
FBA3
FBC4
FB5C
FAE8
FB04
FB89
FBB7
FB43
FACF
FAFC
FB6B
FB36
FA68
FA79
FCC8
00CF
045F
05BE
054B
04B6
04F7
0583
056F
04CC
046F
04BF
0535
052F
04D5
04C2
051D
0563
0529
04B3
0483
049E
049C
045A
0439
0487
04F5
04F5
048C
045D
04C5
0547
052E
0498
046C
050E
0574
0410
009F
FCBD
FA72
FA40
FAEC
FB18
FAA9
FA7C
FB01
FBAB
FBBD
FB3D
FAD1
FAD6
FB07
FAFE
FAC6
FAB1
FACF
FAE4
FADA
FAEE
FB4A
FBA6
FBA1
FB4D
FB2B
FB72
FBBD
FB95
FB29
FB18
FB86
FBC4
FB3F
FA9E
FB76
FE86
0294
055C
05C2
04CB
0444
04C9
0571
0548
0492
044B
04C5
0551
054D
04F3
04E4
0530
0555
0517
04DD
0508
0556
0540
04CA
0488
04BC
04F1
04AC
0438
0440
04C8
0508
0483
03D9
0400
04CE
04B9
0271
FE88
FB2C
FA0B
FACF
FBC1
FBBD
FB24
FAF2
FB54
FB93
FB2F
FA99
FA8B
FAFE
FB3F
FAF5
FA9A
FABB
FB29
FB4C
FB0A
FAE6
FB27
FB6B
FB47
FB00
FB2C
FBAE
FBC1
FB22
FAAE
FB47
FC73
FCC3
FBCC
FB13
FC88
0039
0407
05CD
056A
0475
0441
04B2
04F1
04C6
04B5
0512
0579
0562
04E5
049F
04DB
0535
0531
04E3
04BA
04CF
04C8
047D
0453
04A4
0521
0526
04A4
0448
0489
04F3
04C1
0417
03F8
04D0
0574
0425
0096
FC8C
FA36
FA23
FB07
FB63
FB02
FAC2
FB2B
FBC4
FBC7
FB33
FABB
FACF
FB19
FB10
FAC3
FABA
FB20
FB7C
FB5C
FB04
FB05
FB61
FB8B
FB4E
FB2E
FB92
FC02
FBC3
FAFC
FAAA
FB3B
FBCC
FB57
FA65
FAD6
FDB9
01E0
04F1
05C0
0524
04A3
04CF
0526
0519
04C8
04A9
04DC
0508
04EC
04B9
04CE
0527
055E
052B
04C5
049A
04C0
04DF
04B5
047D
048D
04BE
049F
043C
0431
04BC
0531
04D6
0418
042C
0547
05C9
03D7
FFB1
FBCC
FA51
FB01
FBDE
FB9F
FAC4
FA6B
FAC3
FB14
FAEE
FAB6
FAEE
FB63
FB79
FB0D
FAAF
FADA
FB49
FB61
FB05
FAB9
FAE3
FB45
FB6B
FB58
FB6F
FBB1
FB9A
FAF1
FA6E
FAE3
FBEE
FC29
FB0C
FA15
FB66
FF3A
035F
056F
052D
0453
045C
0513
0566
0508
04A7
04D8
054E
0566
0505
04AC
04C0
050F
051F
04DA
04A2
04C7
050C
0502
04A5
046B
049B
04EE
04FB
04D4
04DF
0522
051E
04A9
0472
0517
05D6
04E5
018F
FD6A
FAE2
FAB8
FB86
FBAD
FB18
FAC7
FB27
FB8F
FB60
FAEA
FADA
FB36
FB6A
FB2D
FADE
FAEB
FB43
FB7F
FB6F
FB3C
FB1F
FB1E
FB23
FB31
FB5D
FB93
FB89
FB14
FA81
FA61
FAE3
FB74
FB54
FAA4
FAB9
FCDA
00B0
0445
05DE
058F
04CD
04AD
04FC
0503
04AA
0479
04C2
0525
051C
04A9
0449
0458
04BF
052B
055F
054E
0506
04AA
045E
043F
0458
0490
04BA
04C3
04CE
0503
053F
0535
04E7
04C7
0512
0510
0388
002B
FC66
FA42
FA62
FB7B
FBED
FB70
FAE3
FADC
FB05
FAE3
FAA4
FAC6
FB44
FB86
FB39
FACB
FAD9
FB5D
FBC0
FBA1
FB45
FB1F
FB3E
FB52
FB38
FB2B
FB5F
FB9C
FB7D
FB12
FAF1
FB62
FBC9
FB6A
FAC0
FB6C
FE61
0270
053D
05AC
04DC
048F
0518
0575
0512
0499
04C9
054D
0553
04D2
048C
04DB
053A
0525
04D8
04CE
04ED
04B7
0433
0410
049D
0539
0521
0482
042F
0474
04C5
049B
0431
0410
0448
0472
0475
04B1
053D
0545
03A6
004D
FCA6
FA6E
FA31
FAFE
FB8A
FB63
FAF9
FAD1
FAE3
FADC
FAB6
FAB7
FAF4
FB28
FB1D
FAF7
FAFC
FB2E
FB63
FB8A
FBB0
FBC6
FBA2
FB4B
FB12
FB2C
FB6B
FB83
FB7E
FB95
FBA8
FB5E
FADB
FAD7
FB94
FC36
FBBA
FA94
FAA2
FD29
013A
0482
059D
0528
049E
04AC
04F4
0505
04EB
04DE
04E0
04DA
04D8
04EE
0505
04F1
04B0
0475
0467
0478
0487
0493
04B3
04D9
04D8
04AB
0488
049A
04BB
04A2
044F
042D
0482
04F4
04D7
0432
03F8
04D9
05E6
051A
019E
FD1E
FA49
FA29
FB51
FBCD
FB3A
FAAC
FADC
FB4D
FB45
FAE2
FAC3
FB0B
FB4B
FB42
FB29
FB32
FB39
FB22
FB27
FB7F
FBE0
FBC7
FB36
FAD4
FB10
FB87
FB92
FB32
FAFF
FB40
FB88
FB70
FB3C
FB75
FBF8
FBF2
FB0E
FA61
FB98
FF11
031A
0576
058C
04BD
049C
053F
0594
050E
045E
0465
0503
0559
0513
04C0
04DA
0516
04F2
048E
0474
04BD
04F3
04D1
04AE
04E3
0529
04FB
046D
041B
0447
0481
046D
045F
04BE
053A
052C
04AB
0493
0521
051C
030F
FF33
FB9E
FA2E
FAB4
FB7C
FB62
FACD
FAB0
FB26
FB77
FB37
FAC7
FAB0
FAE5
FAF1
FAB9
FAA3
FAF6
FB65
FB76
FB30
FB07
FB30
FB62
FB56
FB2D
FB28
FB3B
FB2B
FB11
FB3B
FB9C
FBAD
FB35
FACD
FB16
FBA6
FB74
FA8F
FAA6
FD39
0183
04FB
05F9
0541
04AF
04F5
054A
050A
04B1
04EB
056C
0564
04CA
0474
04DF
057B
0578
04DE
0466
0471
04A8
04AF
04B0
04F5
054E
0544
04DA
049C
04D0
050D
04E0
048D
04B0
053C
0565
04C2
041B
046E
0546
04C3
01B7
FD5A
FA48
F9D1
FAD9
FB7A
FB2E
FAD3
FB06
FB4D
FB0C
FA8E
FA8E
FB04
FB2C
FAB8
FA53
FAA2
FB4C
FB7E
FB1D
FAD7
FB0D
FB50
FB21
FABC
FAAC
FAED
FB00
FACF
FAE4
FB77
FBE4
FB8B
FAD7
FAC3
FB60
FBA2
FAF4
FA76
FBEE
FF90
0377
0593
05B3
0541
0550
059B
056F
04E7
04B9
051F
0584
055C
04DF
04AF
04F2
053C
0535
050B
0509
051D
0504
04CF
04CF
050D
052A
04EC
04A0
04A6
04DF
04D9
0491
0482
04D9
0509
0494
03FF
044B
0556
0577
0332
FF2A
FBAE
FA5F
FAB5
FB0C
FAAA
FA37
FA6C
FAFE
FB29
FAC8
FA78
FAA6
FB0B
FB28
FAF3
FACC
FAF4
FB48
FB88
FB98
FB83
FB4F
FB0A
FADF
FAF0
FB1C
FB25
FB04
FAFD
FB3D
FB84
FB6F
FB10
FAE8
FB37
FB86
FB38
FAA3
FB25
FDC2
01BF
050F
063F
05B6
04F5
04DA
0512
0502
04BF
04C8
0527
055E
0526
04D3
04CB
04F1
04E6
04A4
0485
04B0
04D9
04BD
0486
048A
04C6
04E7
04D3
04C5
04DF
04EA
04BA
0491
04C4
0519
04FE
0478
0457
051D
05D7
04C0
013E
FCEA
FA2A
F9DC
FAC6
FB3B
FAE4
FA9B
FAED
FB64
FB59
FAEA
FAC1
FB13
FB68
FB53
FB06
FAF7
FB31
FB5C
FB58
FB62
FB98
FBB1
FB71
FB19
FB13
FB54
FB66
FB1F
FADF
FAF4
FB17
FAE5
FA9B
FAD8
FB81
FBA1
FAC6
FA21
FB8E
FF59
0390
05EB
0608
0564
0549
0582
0534
0461
03F6
046D
0525
0541
04C6
0470
04A1
04ED
04D5
0479
0456
0490
04CB
04C4
04A4
04AE
04D4
04E5
04E9
050C
0539
0526
04D5
04B2
04F6
0537
04F2
046D
047B
0525
0510
02D6
FEE8
FB77
FA41
FADD
FB8B
FB58
FAD6
FAD8
FB30
FB29
FABD
FAA4
FB33
FBCF
FBC8
FB52
FB20
FB59
FB76
FB25
FAD5
FB04
FB7C
FB9C
FB41
FAED
FB02
FB3B
FB2F
FAFA
FB01
FB3A
FB3A
FAF9
FAF7
FB6B
FBB1
FB24
FA6A
FB33
FE4E
0269
0535
05B7
0505
04AF
0508
054C
0508
04B3
04CD
0517
0502
0494
0461
04AC
050C
0514
04EB
04F2
0511
04DE
045E
0426
048C
051D
0530
04D3
04AA
04F1
052C
04EC
0485
048E
04EB
04F4
0488
046A
0509
056C
03F9
0075
FC99
FA6C
FA4B
FAF3
FB39
FB2A
FB5A
FBC3
FBD6
FB61
FAE3
FACF
FAFC
FB06
FAF4
FB16
FB67
FB7F
FB2E
FADE
FB03
FB7D
FBC8
FBBA
FBA5
FBB9
FBA9
FB36
FABC
FAC9
FB3C
FB5E
FAF1
FAAD
FB3F
FC19
FBFB
FAD3
FA5D
FC5F
0075
043E
05CA
0563
04AF
049F
04C5
0483
041C
0438
04DF
0566
0561
0514
04EB
04E0
04B8
0480
0476
048C
046F
0418
03FD
046F
050E
0537
04DE
0498
04C0
04FE
04E2
04A1
04BE
0520
0513
0467
03FC
04AA
05C1
0559
026A
FE34
FB18
FA3D
FABC
FB19
FAE9
FAC8
FB19
FB73
FB5D
FB05
FAE7
FB0C
FB16
FAEA
FAE5
FB4B
FBCB
FBE9
FBA9
FB7A
FB90
FBA7
FB7B
FB38
FB2C
FB45
FB34
FAFE
FB00
FB55
FB86
FB35
FAC0
FAD8
FB71
FBA5
FB04
FA8D
FBD9
FF33
02FA
0536
0581
050E
0504
0556
0555
04DB
0477
0494
04F0
0516
04FF
04F2
04FF
04E4
048C
043F
0441
0471
0485
047B
0493
04D6
04FF
04E5
04C2
04D6
04F6
04C4
045A
044B
04D5
0562
0538
0489
0449
04D5
0519
0394
0027
FC79
FA5F
FA2C
FABD
FAFB
FAD9
FADE
FB30
FB6E
FB53
FB12
FAFE
FB16
FB29
FB2F
FB49
FB77
FB7E
FB44
FAFA
FAE2
FAF9
FB0A
FB09
FB1F
FB62
FBA2
FBAD
FB8F
FB73
FB53
FB10
FACC
FAEA
FB74
FBCC
FB51
FA74
FAAE
FD15
0106
0486
060F
05CD
0510
04CE
04F2
04FD
04D5
04BC
04D0
04E2
04D4
04D0
04FD
0533
0529
04DE
049F
04A1
04C9
04E3
04EB
04F5
04F5
04D0
049D
049B
04D0
04EC
04B3
0468
047C
04E5
0518
04C9
0478
04C1
0544
04A7
020A
FE3B
FB22
F9F7
FA45
FAC8
FADC
FACD
FB01
FB55
FB6D
FB4A
FB37
FB43
FB34
FAF6
FAD3
FB06
FB53
FB55
FB0F
FAE9
FB15
FB47
FB2D
FAF2
FAFF
FB56
FB85
FB4B
FB00
FB08
FB3E
FB31
FAEF
FB01
FB8A
FBD7
FB53
FAB6
FBA4
FEC9
02C0
0552
05A8
04E5
0497
0505
0560
0525
04C0
04CB
052B
0551
0517
04E0
04F4
051C
04FF
04AC
0479
048C
04BA
04DB
04F3
0506
04F3
04B8
0493
04B8
04F6
04F5
04BD
04B1
04E4
04D9
0441
03BC
043C
0588
05E0
03B0
FF81
FBB2
FA2D
FAAA
FB73
FB73
FB09
FAFA
FB47
FB5C
FB09
FABE
FAD4
FB16
FB22
FAFE
FAF4
FB16
FB2A
FB1A
FB1A
FB4A
FB74
FB57
FB17
FB0C
FB44
FB70
FB5B
FB2F
FB1E
FB10
FAE1
FACB
FB27
FBCB
FC0C
FB9F
FB1B
FB37
FBB6
FBA4
FADF
FAC3
FCCC
00A4
042D
05A6
055B
04E3
0522
058B
0551
04A6
045F
04C5
053F
0538
04D6
04A4
04C8
04F2
04E9
04CE
04CD
04DD
04E2
04E8
0505
051A
04FF
04C7
04BC
04E8
04FC
04C2
0472
0468
049D
04BB
04A6
04A3
04D6
04EA
0496
043C
047C
0513
04AA
023C
FE7E
FB6B
FA53
FAB6
FB2F
FB14
FAD9
FB00
FB55
FB58
FB12
FAFF
FB4A
FB93
FB7C
FB2D
FB04
FB13
FB20
FB17
FB25
FB62
FB95
FB83
FB3F
FB0B
FB00
FB0B
FB2D
FB77
FBBD
FBAA
FB37
FAE2
FB1D
FBA3
FBC3
FB55
FAFB
FB2F
FB7A
FB25
FA9B
FB69
FE7A
02A7
0595
060C
0500
0435
0457
04BF
04C4
0493
04A7
04F6
050F
04D6
04AD
04DC
052A
053F
051B
0501
04FD
04DD
0491
044D
043C
044A
0456
0474
04C4
051C
052D
04F1
04B8
04B3
04B0
0486
0476
04CD
0541
052E
048E
0446
04EB
0595
047C
011D
FD27
FAE5
FAE2
FBA0
FB92
FAC4
FA4D
FAA7
FB2C
FB2A
FACF
FAB7
FAF8
FB23
FB07
FAFC
FB4B
FBB6
FBD0
FB94
FB5E
FB57
FB4C
FB18
FAEE
FB05
FB3C
FB4C
FB36
FB39
FB5B
FB5B
FB20
FAED
FAF9
FB07
FACA
FA84
FACB
FB8F
FBE6
FB49
FAB5
FBF0
FF66
0355
0572
053D
0447
0436
0511
05C4
05BA
056D
0572
05A4
057B
04EC
047D
048C
04DF
0507
04EB
04C4
04B8
04BC
04C1
04CE
04E2
04ED
04EC
04EE
04EF
04D3
049E
048F
04CB
0511
04FB
04A2
0494
050B
057B
0543
04AA
049E
0540
053D
0323
FF49
FBCF
FA7A
FAF7
FB88
FB20
FA4F
FA1D
FAA4
FB20
FB1A
FAE3
FAF4
FB37
FB46
FB12
FAED
FB0B
FB4A
FB73
FB7A
FB63
FB23
FAC6
FA9B
FAE4
FB69
FBA8
FB72
FB2E
FB4C
FBAD
FBDB
FBAD
FB67
FB3E
FB14
FAD9
FADA
FB50
FBC8
FB91
FAE6
FB2D
FD90
016F
04BD
05FC
0590
04F2
04F2
052C
0506
04A4
048D
04D6
0508
04DB
0494
0498
04DE
0510
0500
04D5
04BE
04BC
04C3
04D6
04EB
04E7
04C5
04AE
04BB
04C4
0498
0460
0472
04C4
04D3
0457
03D3
0400
04C6
053B
04E1
046E
04C4
0566
04A2
0194
FD88
FAD8
FA7D
FB4F
FBA7
FB2F
FABA
FAD4
FB19
FB0D
FAE5
FB1B
FB9B
FBD2
FB8C
FB3C
FB51
FB92
FB84
FB25
FAEA
FB17
FB67
FB7F
FB61
FB47
FB3D
FB2C
FB29
FB66
FBC8
FBE6
FB9C
FB54
FB74
FBBB
FBA0
FB31
FB19
FB96
FBEA
FB58
FA94
FB6D
FEB7
02FB
05BF
0602
04FE
0475
04CF
0533
0504
049E
0498
04DA
04D9
0474
0419
0423
0469
048C
0470
0447
043C
0458
049E
0500
0542
0520
04A9
0447
0441
046B
0478
0475
04A9
0501
050B
049A
042B
0446
04B0
04B7
044C
043E
04F4
055B
03C3
FFFA
FBEF
F9E7
FA45
FB7B
FBF6
FB99
FB35
FB2B
FB27
FAF0
FAD9
FB37
FBC6
FBFD
FBC5
FB85
FB80
FB8B
FB6D
FB49
FB5F
FB9B
FBB1
FB91
FB79
FB8A
FB95
FB6B
FB39
FB47
FB89
FBA9
FB89
FB62
FB58
FB38
FAE7
FACA
FB46
FBFB
FC02
FB3D
FB01
FCDE
00AD
0464
0608
0591
0499
046E
04F5
0556
053C
04FD
04E1
04CC
049A
047B
04A3
04E1
04D5
0478
0427
0432
0480
04CE
04F3
04EB
04B1
0454
0415
042E
047A
0493
0459
042F
046B
04D5
04F2
04BF
04B1
04F6
0516
04B2
0449
04AA
0588
0544
02A2
FE76
FB17
FA0E
FABA
FB67
FB41
FACD
FAB7
FAE1
FAD1
FA93
FAA2
FB23
FBA2
FBBC
FB94
FB84
FB87
FB53
FAE5
FAA3
FAD5
FB4B
FBA1
FBB8
FBAE
FB92
FB69
FB5F
FBA7
FC18
FC35
FBC7
FB3C
FB1E
FB5A
FB61
FB12
FAFD
FB7C
FBF4
FB93
FAC3
FB2C
FDEB
0200
0521
05FC
0557
04CC
04FA
054E
0535
04E7
04DB
050D
051A
04E7
04BF
04C6
04C9
049E
047E
04AB
04FA
0505
04BA
0478
048A
04C6
04D7
04B1
0485
0465
043C
041E
0442
0499
04BA
046D
041F
0453
04D4
04DC
043A
03CF
0463
0536
0471
0146
FD2C
FA87
FA42
FB33
FBBC
FB7D
FB28
FB30
FB41
FAFC
FAA7
FAC2
FB46
FBAD
FBA8
FB65
FB2E
FB0A
FAEA
FAE9
FB1F
FB62
FB68
FB39
FB31
FB75
FBB7
FBA1
FB57
FB40
FB6F
FB99
FB93
FB90
FBB5
FBC4
FB86
FB52
FBAD
FC5B
FC63
FB6E
FAB7
FC0B
FFAA
03B6
05F5
05F8
051C
04C3
0501
0530
0512
04FB
050D
04F8
0490
0432
0450
04CB
051D
0506
04C9
04B0
04B0
04AB
04BB
04FC
0531
04FC
0471
0418
043D
048F
0498
0467
0464
04A4
04C4
0497
047A
04BB
04FB
04AA
0407
03FF
04C0
04F8
0316
FF46
FB93
F9DF
FA19
FAC6
FAE2
FAB3
FACE
FB1C
FB21
FAE2
FAE5
FB56
FBB8
FB98
FB31
FB10
FB4B
FB78
FB58
FB25
FB1D
FB27
FB17
FB0F
FB51
FBB6
FBC5
FB60
FAFC
FB08
FB53
FB71
FB61
FB81
FBCF
FBCD
FB4E
FAF2
FB56
FC0A
FC03
FB43
FB5F
FDCA
01DB
0534
0637
0589
04F1
052F
058F
0552
04CA
04B6
051D
055A
051D
04C2
04B0
04C1
04A6
0480
04A7
0512
054E
052B
0502
051F
0541
0503
0486
0452
0489
04B0
0469
0406
040E
0473
04B1
04A7
04BA
0505
04F3
0422
0355
03B2
04F3
0511
0263
FDC2
F9F9
F8F5
FA0B
FB32
FB5C
FB11
FB19
FB5B
FB51
FAFA
FACE
FAEF
FB00
FAC1
FA7E
FA90
FAD8
FAFB
FAF8
FB16
FB52
FB4E
FAEB
FA9A
FAD2
FB61
FBB5
FBA4
FB97
FBCB
FBE9
FB90
FB0E
FAFF
FB69
FBB0
FB84
FB57
FB95
FBCD
FB53
FAA0
FB5D
FE81
02D0
05DA
066A
0581
04D8
04F5
0528
04EF
04AF
04EA
0567
0588
0530
04D4
04C8
04E3
04ED
0502
054C
0593
0580
052B
0509
0541
0566
051F
04AA
0486
04B0
04B0
045C
041F
0455
04B7
04C3
048A
048F
04EE
051A
04C2
0471
04B9
04FC
03C1
0085
FCB8
FA71
FA44
FAEF
FB13
FAAA
FA8B
FAF3
FB44
FB0F
FABE
FAE7
FB71
FBB7
FB70
FAF8
FAB4
FA9E
FA8C
FA9A
FAF2
FB5A
FB62
FB00
FAAD
FAC1
FB02
FB0D
FAED
FB03
FB5F
FBA3
FB95
FB77
FB89
FB91
FB3A
FAC7
FADD
FB7D
FBCE
FB50
FAF7
FC65
FFE3
03AF
05B6
05A9
04F1
04CD
051D
051C
04BC
04A1
050D
056F
0533
0492
0439
045F
04A1
04AF
04AE
04D5
0505
0503
04F0
0520
058A
05BC
0572
04F8
04BC
04BF
04B6
0495
04A4
04F3
0528
04F8
049C
0479
048B
0483
0475
04D8
0586
053C
02CB
FEC1
FB4D
FA25
FACC
FB69
FAFD
FA47
FA62
FB38
FBC4
FB8B
FB1A
FB17
FB5F
FB69
FB23
FB01
FB37
FB73
FB62
FB2C
FB1D
FB22
FAED
FA8A
FA65
FAAF
FB18
FB3C
FB20
FB13
FB25
FB1B
FAE6
FAC5
FAE3
FB0D
FB0B
FB05
FB48
FBB4
FBD0
FB84
FB50
FB90
FBD6
FB79
FAD3
FB54
FDF3
01CD
04C9
05AE
052E
04D3
0534
05A8
0570
04BC
0442
044B
0482
0494
04A2
04E6
0542
0569
054D
052C
052C
052B
050C
04F1
050C
0549
0565
0547
0516
04F3
04D0
04A7
04A5
04E4
0527
0513
04B7
0484
04AE
04DC
04B0
045A
044F
0485
0479
0418
0415
04EC
05B4
04B7
0165
FD4D
FAB0
FA4B
FAFB
FB58
FB23
FAF6
FB1A
FB36
FAFF
FABB
FAC9
FB14
FB3C
FB25
FB0E
FB1C
FB2B
FB18
FAFD
FAFE
FB12
FB18
FB15
FB28
FB41
FB2D
FAED
FAD5
FB22
FB97
FBBE
FB7F
FB38
FB39
FB5F
FB65
FB57
FB79
FBC4
FBD6
FB80
FB2D
FB55
FBB8
FB92
FAC7
FA84
FC34
FFD1
039A
05B2
05D3
053D
051D
056E
057F
051B
04C4
04DD
0528
052E
04F2
04D4
0505
0544
0548
0515
04E1
04C7
04C4
04DC
0511
053A
0523
04D9
04AB
04BC
04CD
049B
044B
0435
0469
049C
04A3
04B0
04EB
0514
04D6
045F
043E
0493
04CD
0488
0445
04C1
05A6
0568
02E3
FED9
FB68
FA0A
FA5C
FAF1
FAF2
FAA7
FA9E
FAE0
FB0A
FAF0
FACB
FADC
FB1E
FB5B
FB69
FB4A
FB13
FAE7
FAE2
FB08
FB39
FB4A
FB3D
FB37
FB50
FB70
FB76
FB6E
FB7E
FBB1
FBE0
FBE2
FBC3
FBA1
FB75
FB22
FABD
FA9C
FAEA
FB57
FB70
FB3B
FB37
FB9C
FBE7
FB87
FAF7
FBA1
FE5A
022B
0507
05CA
0536
04D1
0531
05B0
0591
04F3
0479
0472
04A1
04C5
04EC
0531
056F
0571
053E
050D
04EF
04C9
0491
046A
0469
0472
045F
0438
0427
043A
0459
0475
049A
04C7
04D6
04BC
04AA
04D3
050E
04FA
0481
0408
03FB
0441
0471
047C
04C9
0572
05A1
0421
00C6
FCF6
FA91
FA44
FB19
FBA0
FB57
FAC6
FA95
FAC7
FAF2
FAE2
FAC9
FADB
FB09
FB26
FB30
FB46
FB6B
FB82
FB78
FB66
FB69
FB7D
FB83
FB6D
FB4D
FB3D
FB49
FB6D
FB92
FB98
FB75
FB4E
FB59
FB98
FBC9
FBB1
FB71
FB57
FB73
FB84
FB5E
FB3D
FB65
FB9D
FB64
FAD3
FAFB
FCF1
0076
03E7
05A9
0598
04DF
049E
04F1
0548
0549
051A
04FF
04FA
04EF
04E3
04EE
0504
04FE
04D9
04BE
04CB
04EC
04F8
04EC
04DD
04D6
04CA
04BA
04B5
04BA
04A8
0476
044D
0460
0498
04AD
0487
0469
048B
04C3
04C0
0488
0479
04BD
0500
04EF
04CD
0510
056D
04B0
0205
FE2C
FB16
FA12
FAAC
FB6F
FB79
FB15
FAE5
FB02
FB1C
FB14
FB17
FB34
FB33
FAF3
FAAF
FAB1
FAEE
FB17
FB0D
FB02
FB22
FB4F
FB54
FB39
FB31
FB49
FB56
FB3C
FB1D
FB22
FB42
FB5B
FB72
FBA6
FBE2
FBDB
FB78
FB07
FAF0
FB36
FB7F
FB9D
FBB2
FBCA
FB91
FAD8
FA56
FB60
FE7A
0274
0543
05E1
051C
047E
04AE
052D
055A
053A
052E
053F
052C
04EA
04C0
04D1
04E2
04B7
0483
049D
04FE
053A
051B
04E4
04EB
051F
0533
050F
04E4
04CB
04A9
0475
0463
0494
04D0
04C8
0491
048D
04D3
0509
04ED
04C3
04E5
0524
050C
04AC
04AA
0536
0544
0376
FFCB
FC05
FA07
FA16
FAEC
FB53
FB35
FB21
FB4D
FB6B
FB49
FB13
FAFA
FAE1
FAA8
FA83
FAC1
FB4B
FBA0
FB73
FB0E
FAEE
FB2B
FB72
FB87
FB85
FB95
FBA0
FB77
FB31
FB15
FB35
FB54
FB46
FB35
FB52
FB74
FB4A
FAE9
FAC9
FB1B
FB7A
FB74
FB37
FB39
FB65
FB23
FA7A
FAAB
FD01
010B
049E
05F6
056C
04BD
04F1
0583
0594
052C
04F3
0518
0522
04D4
0499
04D1
052C
0516
049D
045D
049C
04EA
04D1
047C
0472
04C1
04F0
04B0
0444
040F
0414
041E
0436
048E
0509
053D
0506
04BF
04C6
04F6
04E8
049B
0478
04A1
04B1
046A
0447
04D3
057D
04B9
01B0
FD8C
FA93
F9F6
FACE
FB6E
FB31
FAC3
FAD8
FB3D
FB57
FB0E
FAD3
FAE4
FB02
FAEF
FADF
FB15
FB6E
FB81
FB42
FB19
FB50
FBAA
FBBC
FB80
FB50
FB5A
FB73
FB74
FB77
FB9A
FBAF
FB84
FB40
FB3B
FB76
FB92
FB63
FB3A
FB67
FBAA
FB8C
FB2F
FB34
FBB3
FBE6
FB4A
FAD4
FC37
FFCE
03CA
05E1
05A7
04B0
048A
0527
0580
052D
04C0
04BD
04EC
04E4
04B9
04D0
0520
0537
04E9
049D
04B9
050B
051E
04E5
04CA
0501
053A
051A
04C3
049A
04AF
04B5
048A
0471
049B
04CC
04AE
0461
044C
047B
0481
0425
03CD
03EB
0446
0448
03FC
0424
04ED
0517
031B
FF2B
FB75
FA05
FABA
FBB7
FBA8
FAF5
FAB6
FB18
FB5B
FB0F
FAA0
FA9D
FAE8
FB08
FAE4
FAD4
FB04
FB28
FAFE
FAB8
FAB5
FAEF
FB0D
FAED
FACE
FAF3
FB3F
FB6F
FB74
FB76
FB7F
FB72
FB4A
FB35
FB57
FB90
FBAD
FBB6
FBD3
FBF3
FBDD
FB9A
FB8A
FBD8
FC09
FB90
FAD8
FB4A
FDE0
01CB
04F3
05EF
054D
04AB
04E4
056F
0577
0501
04B9
04F4
0553
0563
052E
0509
050A
0506
04F3
04FC
052C
054F
0542
0529
052D
0531
0502
04B8
04A0
04CB
04F0
04D9
04B1
04B8
04D4
04BA
0472
0452
0472
047B
0440
0422
047F
04FA
04DA
042D
03EC
04A2
0549
041F
00BC
FCD1
FA81
FA4D
FAFE
FB46
FAFF
FABE
FACF
FAF0
FAE0
FAB8
FAB3
FAD6
FB02
FB2D
FB59
FB71
FB58
FB20
FB06
FB19
FB24
FAF8
FAB2
FAA3
FAE7
FB40
FB5F
FB3C
FB19
FB25
FB45
FB49
FB2C
FB10
FB05
FAFC
FAFE
FB2F
FB89
FBC2
FBA6
FB73
FB95
FBEF
FBCC
FAF1
FA7E
FC13
FFDB
03EF
061B
0603
052B
04FC
0563
0582
052A
04FF
0559
05C0
05B1
055B
0534
053D
051D
04D6
04C4
04F4
04FF
04AB
045F
0499
052B
056B
0526
04DA
04F7
053F
053E
04FE
04DA
04DE
04C4
0485
0478
04BC
04E6
049D
0434
0447
04CD
0509
049C
042B
0485
054B
0502
02A4
FEDD
FB81
F9EF
FA08
FAA7
FADD
FAA0
FA73
FA9B
FAE5
FAFE
FAE1
FACF
FAEE
FB1C
FB27
FB0F
FAFF
FB01
FB04
FB05
FB16
FB1F
FAE6
FA78
FA41
FA8A
FB0C
FB44
FB20
FB03
FB32
FB71
FB72
FB53
FB5C
FB72
FB3B
FAD7
FADB
FB6C
FBE0
FBA4
FB1A
FAFD
FB3B
FB1D
FAB5
FB62
FE40
026C
0593
0658
0593
04F7
051D
056A
0555
0510
04EE
04E2
04C6
04BC
04F0
0532
0530
04F4
04E0
050E
0522
04DE
0496
04BD
0540
059C
058E
054E
0522
0517
0515
0513
0510
0500
04D0
048D
045D
0456
046D
0491
04B8
04D3
04D6
04D5
04EB
04FD
04DC
04A0
04A0
04DC
04DA
0460
03FD
0455
04F4
0462
01C0
FE0B
FB47
FA73
FACB
FB11
FAF2
FAD6
FAED
FAF8
FADA
FAC6
FADB
FAEE
FAE3
FAE3
FB11
FB3B
FB1E
FADD
FADD
FB2A
FB58
FB1F
FAC2
FAA3
FAB8
FAC6
FAD1
FB09
FB5D
FB8B
FB85
FB84
FB9F
FB9F
FB54
FAF0
FAC5
FAD7
FAE4
FADF
FB01
FB51
FB80
FB71
FB69
FB90
FB9C
FB57
FB22
FB66
FBC9
FB8E
FAF2
FB71
FE26
0222
051E
05E2
0558
0509
0545
054F
04DC
0480
04B6
052D
0557
052C
0505
04FF
04DD
0493
046F
04A4
04F2
0504
04EB
04EA
0506
0506
04D8
04A6
0499
04B3
04EB
0530
055F
0556
0519
04D4
04AB
049F
04A1
04B1
04CC
04D0
04A4
046D
0460
0461
0433
0401
0441
04E9
053E
04D5
0459
049F
052A
044D
0136
FD44
FABE
FA5F
FAD7
FAC1
FA3B
FA28
FAA3
FAFA
FADB
FAB4
FAE1
FB1A
FB00
FAC6
FAE2
FB4B
FB82
FB53
FB19
FB21
FB32
FAF9
FA9D
FA7B
FA9C
FAC1
FAD9
FB09
FB4B
FB66
FB48
FB2B
FB41
FB66
FB56
FB19
FAFB
FB22
FB5C
FB79
FB86
FB96
FB99
FB88
FB7F
FB78
FB49
FAFB
FAF1
FB49
FB7F
FB24
FAE1
FC2A
FF85
0381
05F2
0628
0567
052A
0584
05A7
054A
04EA
04DD
04E0
04AF
047B
0494
04DE
04F9
04D3
04BF
04F2
0533
053C
051C
050C
0514
051A
051C
0525
0528
0514
04FB
04F0
04D9
0494
0438
040E
0431
046E
048F
04A0
04C3
04E4
04D7
04AC
04A6
04CA
04D6
04BD
04C3
04EF
04DA
0467
0432
04B8
052E
03F6
008D
FC93
FA4B
FA46
FB0E
FB28
FA9C
FA52
FA93
FADE
FAE8
FAF3
FB2E
FB4E
FB10
FAB7
FAB6
FB0A
FB3D
FB14
FAD5
FACF
FAE8
FAE3
FACA
FACD
FAE9
FAF6
FAF3
FAFC
FB13
FB1E
FB22
FB3C
FB6C
FB85
FB69
FB33
FB10
FB08
FB03
FB05
FB2C
FB74
FBB0
FBC8
FBC6
FBA0
FB3E
FAD7
FAD9
FB3A
FB55
FAD8
FAAB
FC43
FFD9
03BA
05CD
05A4
04A8
0450
04BD
0531
054A
053C
0532
050E
04C8
04A0
04BC
04F4
0506
04F3
04E9
04F6
04FA
04E5
04CE
04CD
04D7
04E5
0503
0526
0522
04F6
04DC
04F3
0506
04DF
04A7
04AD
04E8
04FF
04CD
0494
049A
04C3
04BE
048A
046D
047D
048D
0494
04C1
0502
04F1
0486
0469
04F9
0548
03C7
0031
FC3E
FA12
FA18
FAEE
FB37
FAF3
FAD6
FB10
FB36
FB11
FAE3
FAE3
FAEE
FAE5
FAED
FB2E
FB7D
FB84
FB36
FADE
FAC5
FADD
FAEF
FAEE
FAEF
FAFE
FB0F
FB16
FB0E
FAF8
FAEB
FB07
FB3D
FB53
FB35
FB17
FB2C
FB56
FB54
FB24
FB07
FB1E
FB3C
FB3F
FB4B
FB81
FBA2
FB5F
FAFE
FB17
FB98
FBA7
FAF8
FAB6
FC6D
0014
03C0
0591
057C
04E4
04CF
0514
0522
04EF
04CA
04C1
04B1
04AF
04DE
0510
04F2
0496
046C
04AB
0502
050E
04E1
04D0
04ED
04F0
04BD
049B
04CA
051F
0549
053D
0523
0507
04DC
04B3
04AD
04C2
04C8
04B2
0499
0495
049C
04A7
04C1
04E0
04D7
0496
0465
0489
04C9
04B1
046B
04AC
057F
0598
038C
FFA3
FBE4
FA25
FA5D
FB1D
FB4D
FB01
FAD2
FAE9
FB09
FB09
FAF3
FAD0
FAAF
FAB8
FAF4
FB23
FB06
FAC8
FAC1
FAFC
FB25
FB0E
FAF3
FB1A
FB5D
FB66
FB32
FB20
FB50
FB71
FB47
FB0C
FB11
FB3A
FB3B
FB17
FB12
FB36
FB49
FB32
FB1E
FB30
FB4B
FB4B
FB4B
FB67
FB6D
FB22
FAD0
FAF5
FB5E
FB37
FA6D
FA66
FCA1
00B5
0467
05EA
058B
04EF
0516
059D
05C1
0575
052A
0512
0508
04FA
04FE
050E
050D
04FF
04F9
04F3
04D7
04BC
04CF
0506
0514
04D5
048A
0487
04BB
04D4
04C5
04D6
0519
0535
04F3
049D
0492
04BC
04C7
04B2
04BE
04F3
0508
04D7
049E
049D
04BD
04CC
04E4
0528
054E
04EF
0464
048F
056A
0566
0309
FEE5
FB4F
FA00
FA86
FB39
FB33
FAD8
FAC0
FAD7
FAC4
FA9D
FAB1
FAF6
FB1E
FB12
FAFD
FAF4
FAED
FAF2
FB1B
FB51
FB5A
FB29
FB03
FB20
FB5F
FB7B
FB70
FB77
FB95
FB8A
FB44
FB0F
FB22
FB51
FB63
FB6C
FB8F
FBA3
FB67
FAFF
FAD4
FB07
FB48
FB5A
FB5B
FB74
FB74
FB2B
FAF3
FB42
FBC2
FB8A
FAA6
FAA9
FD08
011C
0495
05DB
0575
04F4
0516
0565
055F
0530
0531
0546
0529
04ED
04D7
04EA
04F2
04EB
04ED
04E3
04A5
045C
0460
04BD
0507
04E6
0491
047B
04AA
04B6
0473
043B
045E
04AB
04C7
04B6
04B3
04C5
04C2
04AA
04A3
04AD
049F
0474
0463
0485
04A9
04A8
04AD
04E1
04FA
049B
041A
0442
04F6
04B9
0241
FE40
FAF6
F9EF
FA9B
FB56
FB46
FADB
FAC1
FAF2
FB05
FAE9
FAE4
FB17
FB56
FB6E
FB52
FB17
FAEC
FB07
FB54
FB7D
FB50
FB11
FB26
FB7F
FBA0
FB4C
FAE4
FAE5
FB37
FB5C
FB34
FB2C
FB82
FBD9
FBC7
FB72
FB3D
FB2F
FB0D
FAE5
FB04
FB67
FBA4
FB80
FB4B
FB5E
FB87
FB67
FB2E
FB5A
FBB7
FB72
FA92
FAA8
FD2F
0172
04EF
05ED
051E
046C
04AB
0521
0501
0494
0490
04F2
051B
04CD
0476
047A
04AB
04A7
0467
043E
046B
04D3
0526
0532
050C
04E8
04DE
04DD
04C8
04A5
0497
04AF
04CB
04BD
048E
046F
046A
0459
043F
0450
0493
04BB
049D
047C
04AA
04FA
04F8
04A2
047F
04CF
0508
04A9
0432
048B
055E
04E5
01F0
FDB0
FAAF
FA2D
FB18
FBAD
FB63
FAEC
FAD6
FAEA
FAD8
FACF
FB0C
FB52
FB41
FAF6
FADB
FB06
FB29
FB1B
FB13
FB38
FB61
FB50
FB1A
FB02
FB10
FB10
FAEC
FADD
FB0F
FB58
FB74
FB69
FB6C
FB8C
FBA4
FB99
FB7D
FB70
FB7C
FB99
FBAB
FB9B
FB6F
FB50
FB52
FB55
FB2A
FAF3
FB1B
FBB3
FC13
FB96
FACA
FB4B
FE0F
020A
0505
05C6
050A
0467
0497
0523
055D
053E
052E
0559
0589
057E
0536
04DD
04A0
0499
04B9
04DC
04EE
0505
052D
0544
0523
04DD
04B0
04B8
04CF
04C5
049F
0485
0483
047F
0479
0491
04CA
04EB
04CA
0483
044D
043A
0444
046F
04AF
04D2
04B5
0491
04B2
04F4
04D2
0438
03F1
04A6
058A
04BF
017A
FD44
FA94
FA48
FB10
FB49
FABF
FA57
FA87
FAD5
FAC2
FA8D
FAB3
FB1F
FB50
FB1E
FAE3
FAE8
FB09
FB08
FAF1
FAF4
FB09
FAFD
FAD0
FAC9
FB15
FB81
FBB4
FBA1
FB81
FB78
FB73
FB5F
FB57
FB7B
FBB3
FBC5
FB9F
FB6C
FB53
FB45
FB23
FB0C
FB40
FBA2
FBA9
FB21
FAE4
FC50
FFBF
03B6
0613
0617
0501
0482
04F3
0564
0523
049C
048A
04E8
0523
050A
04F7
0522
053D
04FD
04A6
04AC
0500
0520
04E4
04B5
04E2
051E
04F9
049B
0483
04C3
04DD
0486
0412
03FF
0446
047D
047E
048B
04C1
04DB
04AC
0478
0486
049B
0457
03F6
0424
04D7
04CE
02BE
FEF3
FB5A
F9B4
FA01
FAD6
FB13
FACC
FAA5
FAD4
FB02
FAF5
FAE2
FB01
FB31
FB2D
FAF8
FADF
FB02
FB1F
FAF5
FAAD
FAA3
FADD
FB06
FAE6
FABD
FAE3
FB4A
FB8C
FB76
FB4A
FB5C
FB9E
FBBF
FBA0
FB72
FB60
FB60
FB5C
FB60
FB6B
FB5E
FB3B
FB47
FBA0
FBD9
FB6E
FAC4
FB44
FDF1
01FD
053F
0648
05AA
04FB
0502
0546
0530
04E7
04E2
051A
051D
04CB
048A
04A6
04E4
04E8
04C3
04CD
050B
0524
04E7
0491
0478
049B
04BE
04C6
04CE
04DD
04D3
049A
0451
0422
040D
0409
042D
0488
04DA
04C9
0467
0436
0485
04EC
04C9
0439
0418
04CF
055C
041B
00A8
FC95
FA0C
F9BF
FA8C
FAFE
FAC2
FA7F
FAA4
FAEB
FAED
FAC5
FAD0
FB10
FB2F
FB13
FB05
FB37
FB6F
FB59
FB0F
FAEF
FB12
FB30
FB19
FB04
FB32
FB7A
FB80
FB42
FB22
FB52
FB93
FB9C
FB86
FB88
FB87
FB48
FAF8
FB12
FB9F
FBFC
FBB2
FB37
FB5B
FBFE
FC0F
FB2A
FAA5
FC4E
002A
041A
05FA
05B8
04EE
04DC
0546
055D
050A
04E0
051E
055E
0544
0500
04F0
050A
0508
04E9
04F7
0540
055F
0506
047F
0459
04B4
0518
051F
04EB
04D7
04E4
04CC
047C
043E
0449
047B
0499
04B2
04EC
0521
04F9
0481
0442
048B
04F0
04DC
0480
049E
052C
04CF
0238
FDFE
FA70
F955
FA37
FB32
FB25
FA98
FA80
FAE6
FB1D
FAE2
FAAE
FAE4
FB48
FB6B
FB52
FB4E
FB62
FB39
FAC4
FA72
FA9F
FB0B
FB27
FAD6
FA8B
FAA5
FAFD
FB36
FB3D
FB46
FB65
FB76
FB66
FB58
FB60
FB5A
FB2A
FAFC
FB09
FB37
FB39
FB14
FB2C
FB9A
FBCA
FB3E
FAA3
FB8B
FEB8
02EA
05D4
0652
0559
04A3
04D9
0551
054F
04F7
04D7
0507
0526
0500
04D6
04EB
051D
0522
04FF
04F4
0513
0521
04F9
04C3
04B6
04C7
04C7
04B5
04BF
04F2
0521
051D
04F1
04B8
0477
042F
040A
0437
0492
04BF
04A8
04A7
04F4
052F
04D4
041E
03F9
04B9
0537
03C8
0033
FC45
FA20
FA2D
FB0C
FB5A
FB08
FADD
FB26
FB65
FB2F
FAC8
FAB5
FAFE
FB35
FB17
FAD7
FABC
FACA
FADE
FAFB
FB32
FB66
FB61
FB25
FAFB
FB12
FB42
FB4C
FB3A
FB43
FB71
FB92
FB8C
FB7E
FB84
FB7D
FB52
FB3F
FB8E
FC0D
FC1F
FB92
FB04
FB1C
FB8C
FB67
FA9B
FA8C
FCB2
00AC
0455
05DA
0579
04D8
04FC
0572
0559
04B8
0457
04A5
0533
0564
052A
04E9
04E0
04F3
04FE
0507
0510
0500
04CE
049F
049B
04AC
04A2
0481
0480
04AE
04D4
04BC
047A
0444
0421
03F9
03E6
0429
04B6
0511
04E5
0484
0486
04F0
0519
04A8
043E
04A6
056D
04F1
0220
FDFC
FAD3
F9FD
FAB5
FB42
FAE3
FA3F
FA29
FA94
FADC
FABE
FA95
FABF
FB1D
FB57
FB51
FB34
FB24
FB23
FB30
FB56
FB81
FB84
FB54
FB21
FB1D
FB2E
FB1D
FAEC
FADE
FB12
FB57
FB75
FB80
FBA3
FBC4
FB96
FB28
FAF3
FB3E
FBA6
FB97
FB2B
FB0F
FB71
FB93
FAE0
FA30
FB44
FEC1
0311
05CE
0622
0555
0514
05A0
060A
05BB
0522
04EE
051F
0534
0500
04D4
04F3
0532
0547
052F
0518
0503
04D3
0497
0489
04B8
04E7
04E4
04CB
04D2
04EF
04E8
04B9
049B
04A9
04AA
0471
043C
0469
04DF
0519
04D8
047F
0484
04B9
0499
0435
044D
0523
0595
040A
0058
FC57
FA2D
FA36
FAFA
FB0B
FA79
FA42
FAC5
FB56
FB40
FAB1
FA62
FA97
FAEC
FAF7
FAD0
FACC
FAF2
FB02
FAD9
FAA1
FA8C
FAA0
FACA
FB06
FB4F
FB7C
FB6E
FB3D
FB2B
FB45
FB5B
FB54
FB55
FB84
FBB1
FB97
FB4A
FB2C
FB63
FB9B
FB87
FB5C
FB76
FBA4
FB53
FAA2
FAD5
FD24
0116
04A0
0611
05AA
0501
0516
057F
056F
04EE
04B3
050A
0576
0566
04F5
04AC
04CD
051C
0548
0540
0518
04DB
0495
046D
0478
0499
04AA
04BA
04F6
054F
0574
053C
04E4
04BB
04B8
0494
0449
042B
046C
04C7
04DD
04B4
049A
048F
0443
03C3
03C3
04B5
05B8
050A
01E6
FDAA
FAB2
FA0F
FAB8
FB09
FA94
FA30
FA87
FB2A
FB4E
FAE1
FA8C
FAC1
FB35
FB66
FB46
FB2C
FB46
FB6E
FB77
FB6C
FB56
FB1F
FAC6
FA8C
FAB3
FB16
FB4D
FB33
FB14
FB34
FB6F
FB73
FB41
FB26
FB33
FB2A
FAF3
FAE1
FB32
FB92
FB83
FB2A
FB31
FBBB
FBF9
FB53
FABB
FC00
FF9E
03BB
05EC
05B4
04C2
04B7
056E
05B0
050F
0460
046F
04F4
0525
04DD
04A3
04C6
04FD
04F5
04D0
04D7
04FE
04FB
04CD
04C1
04F4
0524
0515
04F7
050E
053B
051E
04B2
045B
045D
0487
0493
049B
04DE
0533
0524
04A5
044B
047D
04C7
047F
03DF
03E7
04D4
0540
036E
FF77
FB8B
F9CC
FA33
FB04
FAFE
FA88
FA9F
FB4B
FBAF
FB56
FACF
FACF
FB3C
FB6E
FB29
FADF
FAF6
FB40
FB4D
FB15
FAEC
FAFD
FB22
FB34
FB46
FB63
FB5B
FB16
FAD4
FAED
FB49
FB76
FB49
FB1D
FB46
FB90
FB8F
FB54
FB55
FBA4
FBC0
FB65
FB26
FB97
FC41
FC0D
FB03
FAE5
FD58
01AC
052E
05FB
04D9
03F9
045E
0526
0537
04BC
0498
0501
0549
04F8
0478
0466
04BF
050B
0519
051D
052C
0511
04BA
047A
049D
04F0
0504
04C8
0493
0495
049C
047E
0473
04AC
04E3
04A2
0406
03BC
041B
04A3
04A1
042E
0403
046C
04DA
04CB
049F
04FD
057B
04A3
019F
FD97
FAC7
FA48
FB26
FBBE
FB87
FB34
FB5A
FBA1
FB6C
FAD2
FA7A
FAB1
FB10
FB1E
FAF3
FAF4
FB32
FB62
FB51
FB28
FB1E
FB29
FB20
FB0D
FB18
FB31
FB26
FAFC
FAFC
FB46
FB8D
FB7E
FB43
FB4B
FBAA
FBF0
FBC4
FB62
FB37
FB48
FB4A
FB3D
FB73
FBD8
FBC2
FAF2
FA77
FBEA
FF86
037D
05A4
058C
04A5
045F
04C7
0511
04F4
04DC
050B
0529
04DC
0462
0440
048C
04E0
04F6
04F1
0504
0514
04FD
04DD
04EF
0523
0530
0506
04E4
04F3
0503
04DC
04A4
04A3
04CE
04C9
047F
044F
0483
04D3
04C4
0465
043B
0476
049C
0452
040F
0490
0583
055C
02E7
FED9
FB5C
FA01
FA68
FB0F
FB0F
FAC0
FACD
FB39
FB81
FB64
FB2C
FB2C
FB52
FB56
FB26
FAEE
FAD0
FAC2
FAC2
FAE4
FB27
FB59
FB4E
FB21
FB1E
FB60
FBAD
FBBF
FB8C
FB42
FB09
FAF7
FB1A
FB59
FB66
FB05
FA86
FA92
FB51
FBF3
FB97
FAAD
FAF6
FDA8
01CF
0507
05E4
0532
04AE
04F9
054C
04F1
044E
043E
04DA
056C
0570
0523
04F5
04EB
04C4
048D
048D
04CD
04FA
04DA
049B
0487
04A5
04C3
04C9
04C9
04C9
04BB
04B2
04D0
04FA
04D8
0462
0415
0460
04E5
04DC
0438
03F1
04BC
05B4
04F8
01C6
FD9D
FACF
FA43
FAE4
FB3C
FAFA
FAC8
FB11
FB73
FB6F
FB19
FAE1
FAF5
FB15
FB0C
FAF4
FB07
FB45
FB7A
FB7B
FB49
FB04
FAD4
FAD7
FB09
FB38
FB30
FAFB
FAE1
FB10
FB5A
FB74
FB5E
FB5A
FB7D
FB7D
FB28
FAD2
FAF3
FB62
FB5C
FA97
FA1F
FB85
FF11
030F
0557
0560
0485
044C
04E2
056A
0562
0527
052D
0550
052A
04CA
04A0
04CB
04EA
04B2
0465
046C
04BD
04FB
04FA
04E5
04DC
04C0
0489
047D
04CA
0528
0526
04D2
04B2
04FE
0544
051D
04C8
04C2
04EF
04C8
0457
0469
054A
05C7
042C
005E
FC5B
FA3D
FA2E
FAC0
FAE2
FAD2
FB24
FB9B
FB88
FAEA
FA89
FAE1
FB80
FBAD
FB5E
FB16
FB16
FB23
FB12
FB0E
FB3E
FB68
FB45
FAF8
FAE6
FB1F
FB47
FB26
FAFD
FB12
FB30
FAFA
FA8F
FA7A
FAE2
FB45
FB2C
FAE4
FB06
FB73
FB65
FAC0
FAC8
FCE7
00CD
045C
05C0
053A
0482
04A4
0517
04EE
0446
040A
049D
055C
058F
0552
0539
055D
0550
04DD
046B
0463
049E
04B1
0490
048A
04B0
04B4
0477
0455
04A5
0521
053A
04E3
049B
04A7
04B0
046B
0431
0474
04EF
04EF
0483
0494
0568
059B
036D
FF23
FB42
F9F6
FAD9
FBC3
FB7C
FAC8
FACD
FB65
FB8A
FAF4
FA70
FA9A
FB0A
FB17
FADA
FAEC
FB5D
FB9F
FB60
FB04
FAFD
FB28
FB25
FB01
FB1C
FB72
FB85
FB25
FADB
FB36
FBEC
FC33
FBCC
FB44
FB22
FB48
FB5F
FB7A
FBCB
FBF4
FB5E
FA70
FAC6
FD94
01E9
0549
0619
0529
0477
04E4
059C
0596
04F6
04A4
04EF
0539
04F8
0473
044B
049A
04EA
04F0
04E0
04FC
0522
050D
04C7
04A0
04B0
04B6
0488
045A
046A
0498
048C
0440
0413
0444
04A4
04DD
04DB
04BC
0488
044A
0453
04DD
054C
0445
0119
FCFB
FA38
F9F3
FB0E
FB9D
FB0B
FA60
FA8C
FB32
FB62
FAF8
FAA7
FAD9
FB1E
FAF6
FA9E
FAAB
FB22
FB7A
FB63
FB25
FB22
FB4B
FB5C
FB52
FB5C
FB76
FB69
FB36
FB2E
FB74
FBB8
FBAA
FB73
FB64
FB6F
FB4C
FB15
FB3F
FBCD
FC01
FB5F
FACE
FBF9
FF5B
0353
05B2
05E5
052B
04E0
0518
0522
04C9
0490
04CC
0528
0532
0500
04F8
052C
0549
0524
04F3
04F0
04FF
04E6
04A6
0473
0462
045D
0461
048F
04DF
0507
04D1
0478
0467
04AA
04E4
04D9
04BE
04CE
04CD
0464
03D7
03E7
04B0
0501
035E
FFC4
FC06
FA1D
FA4D
FB38
FB93
FB4B
FB01
FAEF
FAD6
FAA7
FABE
FB38
FB92
FB45
FA8C
FA29
FA6A
FADA
FAF7
FAE1
FAFC
FB44
FB53
FB11
FAE9
FB24
FB7E
FB89
FB5B
FB5D
FB9C
FBB2
FB73
FB41
FB6A
FBA0
FB78
FB27
FB3B
FB9E
FB8C
FAE2
FAE8
FD13
0106
0490
05E8
0570
04D2
04E0
050B
04C3
0472
04B7
054F
0567
04E8
04A8
052A
05D9
05DF
0553
0501
0536
0562
0512
049B
0491
04DC
04EE
04A7
0487
04DF
0543
052C
04BB
047B
0493
04AA
049E
04B8
050C
051D
0494
0408
045C
053E
04F8
024A
FE23
FAF2
FA2B
FB03
FBB8
FB8F
FB29
FB28
FB55
FB31
FAD9
FACF
FB16
FB1E
FAA2
FA23
FA43
FAE1
FB44
FB10
FAAD
FA9E
FAD2
FAE3
FAC0
FABD
FB04
FB45
FB30
FAEE
FAD7
FAF1
FAF5
FAD8
FAE5
FB37
FB78
FB6B
FB55
FB89
FBB5
FB45
FAA0
FB51
FE5C
02A5
05AB
0615
04F3
043B
0492
0515
0502
04B5
04DC
0554
0577
052C
0505
054A
057E
052D
04AF
04AA
0513
0545
04FB
04A7
04BE
050B
0519
04F8
0516
057D
05AB
0559
04F2
04F3
0533
0532
04EC
04D2
04FB
04F4
0492
0471
050C
058A
043D
00A7
FC7D
FA1B
FA25
FB28
FB7D
FAF3
FA71
FA7F
FACA
FAE0
FADA
FAFF
FB30
FB1A
FAC7
FAA0
FACF
FB06
FAFD
FADD
FAF1
FB2B
FB35
FAFB
FAD3
FAF7
FB2E
FB23
FAEC
FAE1
FB17
FB42
FB38
FB2F
FB51
FB57
FAF2
FA68
FA5D
FAE3
FB3C
FAEE
FAD3
FC66
FFEC
03BD
05D0
05C0
04E8
04A5
04FA
0524
04E8
04C7
0515
0570
0559
04F4
04CA
0501
053B
0537
0527
0546
0569
054C
050D
0507
0537
0536
04D5
0474
047C
04BB
04B3
0463
0457
04CA
0539
051B
04A4
0473
04A2
04BF
04AD
04E6
057C
054A
0302
FF04
FB7C
FA35
FACB
FB6F
FB20
FA82
FA85
FB0F
FB58
FB22
FAED
FB0B
FB26
FAE4
FA8A
FA8D
FADB
FAFB
FACF
FAB9
FAED
FB20
FB04
FAD9
FB11
FB9A
FBDA
FB87
FB0F
FB05
FB5D
FB9B
FB85
FB53
FB35
FB16
FAF7
FB1B
FB93
FBD6
FB54
FA88
FAF1
FD94
0194
04C4
05B9
0501
0441
0461
04F4
0536
0519
051A
0566
059C
056D
0513
04F6
0511
0515
04F6
0503
055A
0595
0546
0499
0428
043D
0483
0489
0459
0450
048A
04C7
04D5
04CB
04CD
04D3
04CF
04D2
04DA
04B1
0453
043C
04D9
058A
04C6
01B5
FD8A
FAA0
FA2B
FB28
FBC8
FB74
FAF0
FAED
FB29
FB1C
FADE
FAE3
FB22
FB14
FA94
FA31
FA6D
FB01
FB41
FB0C
FAD6
FAF2
FB26
FB24
FB07
FB1F
FB68
FB91
FB77
FB47
FB2F
FB23
FB16
FB29
FB5E
FB62
FB04
FAAA
FAEA
FB98
FBC0
FAF3
FA4C
FB8C
FF12
0323
0591
05D3
0527
04E1
051E
0537
04EC
04A7
04C1
050C
052C
0526
0537
055C
0553
0507
04C2
04CB
0512
0551
0565
055D
0541
0501
04A1
0457
044E
047D
04B6
04E6
050C
0514
04EC
04B7
04C5
051B
0549
04F5
047A
049D
0563
058D
03A9
FFD6
FBFE
FA1E
FA61
FB40
FB52
FAAE
FA52
FAAF
FB39
FB48
FAF3
FAC2
FAE5
FB0F
FB08
FAF6
FB05
FB15
FAFB
FAD9
FAEE
FB2B
FB3B
FB04
FAD6
FAF8
FB3A
FB43
FB1B
FB1A
FB52
FB71
FB48
FB1E
FB3B
FB63
FB37
FAE0
FAE6
FB48
FB46
FA92
FA51
FC27
0023
0439
0639
05FA
051D
04FA
055F
0573
0516
04DD
050D
053E
051A
04E6
0508
0556
0558
0501
04BA
04BE
04CD
04AC
048F
04BA
04FE
04F0
0499
047C
04D0
0518
04D9
0464
047A
0524
0586
050E
0464
0492
055A
0515
0288
FE90
FB6B
FA76
FAFF
FB77
FB40
FAF3
FB1F
FB7C
FB74
FB0F
FADD
FB17
FB5E
FB51
FB16
FB0B
FB30
FB35
FB06
FAE9
FAFE
FB0A
FADF
FAC8
FB20
FBAD
FBCF
FB58
FADE
FAF2
FB57
FB67
FB17
FB06
FB71
FBA4
FB02
FA59
FB5F
FEB4
02CE
0559
0586
0493
0426
049B
0525
0523
04D6
04C2
04F4
0518
0503
04DB
04CB
04CC
04CA
04C8
04C8
04B5
048D
047B
04AA
04F7
0515
04F4
04E3
051A
055E
0549
04E2
04A2
04CA
04FB
04BB
0441
0450
050E
055F
03DA
006D
FCBD
FAAD
FA9A
FB4D
FB82
FB21
FAE2
FB26
FB8E
FBA2
FB70
FB4C
FB44
FB21
FADB
FABD
FAF9
FB5A
FB85
FB6D
FB4B
FB39
FB19
FADE
FABC
FAD5
FB07
FB1E
FB25
FB43
FB58
FB1F
FABC
FAC4
FB6B
FBF5
FB7C
FA65
FA79
FD09
0138
049B
059E
04ED
0455
04B2
0556
055A
04D4
048B
04D2
0534
0530
04D9
0497
0491
0497
0488
047C
0493
04BA
04CE
04D5
04F3
0529
054A
0538
050A
04E4
04CC
04C0
04D0
0505
0530
050A
04AE
04A8
0549
05E0
0501
01FC
FDE4
FAD1
F9F0
FA89
FB14
FAF1
FAC1
FB26
FBC8
FBD4
FB34
FAAC
FACB
FB37
FB4A
FAFC
FADC
FB2F
FB99
FBA2
FB53
FB0B
FAF6
FAFE
FB17
FB50
FB8A
FB7C
FB23
FAE1
FAF2
FB08
FAC9
FA7E
FAC2
FB77
FB9D
FAB0
F9DE
FB21
FEF3
0364
05F0
05F3
04F1
0490
04FF
0565
054D
0514
0520
0546
052F
04EE
04D4
04ED
04FA
04EB
04EB
04FB
04D4
0462
0417
0464
050E
055C
0508
04A1
04B8
050F
04FF
0482
0456
04DE
0576
0545
048B
0463
051F
0563
0387
FFAC
FBEE
FA49
FAB8
FBA2
FBCA
FB5B
FB19
FB31
FB37
FAFA
FAD1
FAFC
FB34
FB19
FAD0
FAD1
FB28
FB5E
FB21
FABF
FAB9
FAFF
FB18
FADD
FABC
FB14
FB93
FBAB
FB5C
FB31
FB65
FB92
FB62
FB30
FB6C
FBB7
FB3D
FA2E
FA32
FCBC
0119
04CF
061D
0593
04FB
0524
0569
051B
0492
0487
04EB
050B
04A8
044E
047F
04F4
051A
04ED
04E6
052B
0556
051B
04C7
04D1
052A
0556
051F
04D2
04B4
049A
044E
040E
0440
04C3
04FD
04B9
0498
0525
05AD
049B
0148
FD16
FA58
FA14
FB32
FBE9
FBA0
FB19
FB14
FB61
FB6A
FB24
FB06
FB41
FB73
FB46
FAEF
FAE0
FB1E
FB48
FB2E
FB0E
FB1B
FB2C
FB0D
FAE8
FB0A
FB5C
FB73
FB35
FB09
FB3C
FB80
FB61
FB03
FAFF
FB66
FB7D
FAE2
FA92
FC21
FFCD
03D0
0603
05F0
0501
04AC
0503
0529
04C1
0457
047B
04F0
0518
04D3
0498
04BC
0500
0502
04CB
04BC
04F4
0522
0503
04C5
04BD
04E9
04FA
04D1
049E
0488
0475
0455
045F
04B4
0503
04D8
046C
0480
0536
054F
034C
FF5F
FBA3
FA0A
FA77
FB39
FB2F
FABF
FAC6
FB34
FB51
FAF4
FABF
FB22
FBA2
FB95
FB12
FAC9
FAFD
FB40
FB2E
FB04
FB23
FB6F
FB72
FB1D
FAE6
FB20
FB7F
FB92
FB61
FB4C
FB62
FB4F
FB05
FAF5
FB5E
FBB7
FB50
FA93
FB0B
FDC3
01D1
04FF
05F0
054D
04AF
04C8
0508
04D2
0461
044E
049D
04D4
04C1
04C0
0514
056A
0552
04EF
04C4
04F2
050D
04CB
0481
04A1
04FD
0505
0495
0433
0450
04AF
04D6
04C5
04DC
051A
0506
047D
0431
04B8
055B
0473
0148
FD36
FA85
FA2D
FB1B
FBAB
FB65
FB08
FB2D
FB83
FB74
FB12
FAF3
FB4C
FBAB
FB9D
FB3D
FAE9
FABF
FA9F
FA9C
FAF3
FB91
FBF0
FBB8
FB43
FB27
FB64
FB78
FB34
FB0B
FB55
FBA6
FB6E
FAEA
FAE4
FB72
FBAC
FB0A
FAA1
FC33
FFF2
03E0
05D5
05A7
04E1
04BA
04FE
04F4
0497
0475
04BB
0501
04F9
04E1
0504
0535
0516
04B7
0482
04A2
04D0
04C9
04A8
04A6
04B9
04AB
0479
0461
0480
04A0
0491
0481
04BD
051D
0519
0488
0414
047B
0564
054A
02F3
FEF7
FB75
FA16
FA8B
FB2D
FAF3
FA55
FA48
FADD
FB4E
FB1F
FAB1
FAA3
FAFC
FB4C
FB5E
FB64
FB84
FB94
FB75
FB56
FB6C
FB8C
FB6A
FB1C
FB08
FB55
FBB4
FBD4
FBC5
FBBD
FBAC
FB65
FB18
FB36
FBB2
FBC3
FAE6
F9FC
FACA
FE14
0280
05AC
0662
0587
04D1
04FF
057E
058B
0535
0506
0526
0532
04EB
0499
04A4
04FC
052F
04FF
04A8
0481
0492
04AD
04C2
04CF
04BC
0470
0426
043A
04A2
04D9
0499
0453
0492
051A
0527
049F
0467
0518
05AA
043D
0067
FC17
F9C3
F9EA
FAED
FB2B
FAA1
FA56
FAC4
FB5F
FB7D
FB2F
FAF7
FB07
FB1F
FB11
FAFE
FB14
FB3E
FB4D
FB45
FB4B
FB63
FB64
FB34
FAFC
FAF8
FB2A
FB54
FB4F
FB40
FB51
FB61
FB3D
FB0B
FB2A
FB8D
FB96
FB08
FAE3
FCB1
00A0
04BC
06A8
060D
04C8
04A5
0577
05DB
053E
046D
0443
0492
04AA
047A
0483
04E9
0529
04EA
048C
0490
04D6
04E1
04A1
0484
04C2
0507
0502
04DD
04EA
0516
0504
04AE
047E
04AA
04D3
049B
0451
048D
0512
049C
022B
FE5E
FB1A
F9D1
FA40
FB03
FB27
FAE4
FADF
FB31
FB64
FB41
FB15
FB32
FB7A
FB9D
FB88
FB6E
FB63
FB50
FB33
FB3A
FB69
FB6A
FB04
FA93
FAA7
FB37
FB9E
FB84
FB5B
FB98
FBE7
FB9E
FAEA
FABC
FB72
FC18
FBA9
FAC9
FB6E
FE91
02C6
0596
0600
051C
0482
04AB
0509
051B
04EC
04B4
047E
044F
0459
04BB
0530
0547
04EE
0489
0478
04AF
04DC
04D2
04AD
0497
0491
0489
0489
04A6
04CD
04BF
046D
0431
045E
04BC
04C0
0463
0451
04EE
0552
03E2
003D
FC1F
F9E4
FA26
FB57
FBBC
FB34
FAC8
FB02
FB66
FB6C
FB43
FB57
FB8C
FB70
FB00
FAC5
FB08
FB6B
FB71
FB2F
FB0D
FB2B
FB49
FB3E
FB29
FB24
FB29
FB40
FB8E
FBFF
FC1C
FB96
FAE1
FADA
FB9E
FC2F
FBA2
FA90
FAC8
FD60
015E
0494
05BA
0564
04FF
052D
056F
0531
04A6
046F
04B4
04FC
04E6
04A7
04A8
04E7
050B
04EE
04C8
04D1
04E7
04D6
04BA
04D2
0504
04EF
0480
042B
0449
049B
04AE
048B
049C
04EA
04F6
0485
0431
04A3
0554
04A8
01B1
FD8C
FA86
F9E4
FACD
FB76
FB0D
FA42
FA24
FAD7
FB86
FB7E
FAEF
FA94
FAC2
FB25
FB4D
FB35
FB1B
FB0F
FAF2
FAD4
FB04
FB8E
FBEB
FB9F
FAF7
FAC5
FB43
FBB6
FB7C
FAF6
FAF7
FB77
FB98
FB1D
FB35
FD40
00EC
0440
05A1
055A
04E0
04FE
0556
055D
0533
0543
0584
058E
0537
04CD
04A5
04B0
04B0
049F
04BA
050B
0544
0520
04C8
04B1
0503
0559
052D
0493
0440
04A5
053D
0525
046A
0423
04EE
05A6
044F
0072
FC0C
F9B1
F9FA
FB35
FB8D
FAE4
FA57
FA80
FAE4
FAE7
FAA1
FA8E
FACA
FB0B
FB24
FB36
FB4E
FB37
FADB
FA97
FAD4
FB67
FBAB
FB50
FAD3
FAD9
FB4C
FB7A
FB0D
FA9A
FAE1
FBA5
FBCF
FAEB
FA28
FB54
FECF
02E1
0560
05B7
050F
04BD
04F2
051D
04F5
04D3
0506
0557
055E
0519
04E0
04E9
0510
0519
04F5
04C5
04B5
04C9
04E5
04EC
04E8
04F6
0513
051C
0507
04F5
04FC
04F7
04C1
049F
04FD
058E
0503
024D
FE34
FB07
FA51
FB47
FBDF
FB35
FA3B
FA25
FAD8
FB4F
FB17
FABC
FAC5
FAF9
FAE8
FAB6
FAD4
FB3A
FB65
FB20
FAD4
FAE7
FB31
FB46
FB1E
FB21
FB7C
FBC7
FB84
FADE
FA95
FB08
FBA0
FB74
FA8B
FA43
FC1A
FFF6
03E3
05CA
0570
0473
045A
0514
0588
0537
04BC
04CB
0540
057B
054E
051E
052E
0543
0519
04E0
04E5
050D
04FD
04B5
04A0
04EC
0531
04FA
0471
0433
047F
04D3
04A3
0438
046F
0572
0608
0498
00F5
FCE6
FA95
FA92
FB7D
FBB8
FB0A
FA73
FAA3
FB27
FB39
FAD0
FA8C
FABB
FAFF
FAF1
FAB9
FABD
FB04
FB25
FAEF
FAB2
FAD4
FB3A
FB70
FB45
FB05
FB05
FB38
FB56
FB4B
FB4F
FB79
FB75
FAF0
FA67
FB22
FDF3
01FE
0526
05FA
0513
043C
047A
053A
0572
0506
04B4
04E3
0531
053C
0537
0572
05AC
0572
04E6
04A1
04D6
0505
04C4
0470
04A7
0544
0579
04E8
0444
045F
0507
0543
04B3
0422
047E
0576
0578
0342
FF54
FBB1
FA19
FA80
FB61
FB75
FAD9
FA82
FAD8
FB3C
FB04
FA6D
FA45
FABF
FB2F
FB03
FA8E
FA7D
FAD9
FB0D
FACE
FA87
FAB2
FB2E
FB77
FB65
FB4E
FB6B
FB83
FB5D
FB2D
FB44
FB6C
FB1A
FA60
FA4B
FC01
FF69
0306
0531
058A
0508
04CB
0506
0538
0516
04F3
0526
0583
0594
0547
0508
0525
0561
0559
051B
050C
0539
0534
04C2
044E
0461
04D4
04FB
0494
042C
0457
04E0
0510
04C1
04A4
0537
05BC
04B5
0194
FDA0
FAED
FA6F
FB3F
FBBF
FB45
FA80
FA59
FAD2
FB2E
FB08
FABE
FAC9
FB11
FB22
FAEA
FACA
FAFE
FB44
FB4E
FB41
FB6F
FBB6
FB96
FB02
FA9C
FAE9
FB8D
FBBB
FB54
FB09
FB49
FB8F
FB21
FA5A
FAB3
FD3E
0140
04B0
060F
0595
04AE
0475
04E9
0557
054F
0504
04E2
04FC
0514
0505
04F0
04F2
04F2
04D0
04AB
04B7
04E4
04E4
049F
0467
048D
04E3
04F5
04B4
048F
04BC
04D9
0483
041A
045E
0532
0548
035D
FFC6
FC54
FA98
FA8D
FB02
FB0D
FAC2
FA9D
FAB4
FAC4
FAB6
FACA
FB27
FB8C
FB92
FB3A
FAEF
FB02
FB45
FB52
FB1A
FAF5
FB27
FB7D
FB99
FB72
FB61
FB9A
FBD8
FBBD
FB5C
FB22
FB2F
FB1C
FAAC
FA83
FBC8
FEDD
02A8
055E
0615
0570
04CB
04DD
054A
0562
0506
04AB
04AE
04ED
050E
04F8
04E2
04ED
04F6
04D7
04B4
04CB
050A
0519
04D2
0478
0457
045F
0455
0448
047F
04EC
0514
04BC
0472
04DD
058D
0501
0249
FE51
FB2D
FA0D
FA55
FAB0
FA9D
FA9B
FB09
FB80
FB6C
FAE7
FA99
FADA
FB50
FB75
FB37
FAF4
FAF8
FB30
FB59
FB54
FB3D
FB3B
FB51
FB60
FB58
FB43
FB30
FB23
FB16
FB17
FB35
FB4A
FB11
FAB0
FB0C
FD21
00C0
0445
05EE
058D
0496
0470
050E
0569
050B
048F
04A2
050E
0528
04D5
04A0
04D3
0512
04F3
04A6
04A3
04E8
04F2
0489
0429
0453
04CD
04F3
04A3
046B
04B2
0510
04E2
0453
0445
050A
0583
0410
0078
FC7F
FA4E
FA66
FB5D
FBA6
FB25
FADD
FB5B
FBFC
FBDA
FB09
FA7C
FAC9
FB74
FBA2
FB2D
FAB7
FAC9
FB3A
FB86
FB7A
FB4C
FB2E
FB1F
FB1B
FB45
FBA2
FBE4
FBB4
FB3B
FB06
FB48
FB78
FB12
FAA5
FB98
FE9D
028F
054B
05C4
04EC
046A
04BF
0521
04E9
047A
0481
04E0
04F2
049B
0473
04D5
053D
0507
0473
0454
04DE
0548
04F1
0442
041A
048D
04E3
04AC
0452
0466
04C4
04D0
046D
0446
04DE
0597
0505
0262
FE7D
FB3B
FA03
FA95
FB74
FB74
FAD3
FA9C
FB21
FB92
FB39
FA89
FA83
FB4A
FBE7
FB9F
FAEB
FAC6
FB49
FBA8
FB70
FB1B
FB33
FB76
FB60
FB15
FB28
FB97
FBB7
FB3F
FAD2
FB16
FBAB
FB9C
FAE9
FAF1
FCF4
007B
03B3
0539
053E
04E7
04FD
0563
0593
0556
04F0
04BD
04C8
04D5
04C4
04B4
04C8
04E1
04C9
0481
0459
0488
04DB
04EF
04B8
0482
047C
047B
0469
0483
04F6
0569
0553
04CE
049A
0516
056A
0428
00ED
FD14
FA94
FA23
FAC3
FB0D
FAAD
FA62
FAC2
FB6F
FB98
FB19
FAA9
FAE4
FB7F
FBBD
FB85
FB6B
FBBA
FBEB
FB79
FAC1
FA99
FB28
FBAC
FB88
FB15
FB02
FB49
FB50
FAFE
FAF6
FB7A
FBBC
FAFA
F9F2
FA7E
FD88
01D5
0517
0608
0555
048D
0493
0519
055C
051B
04B8
04A7
04E3
04F9
04AA
044C
045F
04CB
04F7
049F
0440
0467
04EB
0538
0516
04CE
04A0
047C
0463
0498
0525
0577
0511
0478
04B0
05A3
05A6
0348
FF37
FBBB
FA60
FAB1
FB3F
FB4B
FB21
FB2C
FB49
FB25
FAD3
FABC
FB13
FB9D
FBF4
FBE0
FB7A
FB19
FB0A
FB35
FB43
FB15
FAF4
FB18
FB50
FB53
FB34
FB2F
FB3A
FB1A
FAE6
FB06
FB81
FBA5
FAFB
FA6D
FBAC
FF27
031F
0557
0555
0485
0455
04D4
052D
04F5
0491
048A
04DF
0525
0507
0499
0433
042D
0490
0502
0513
04C2
0478
047D
04A3
04AA
04A0
04B7
04E4
04FE
0502
0503
04EA
04A4
047A
04CE
0547
049E
01EA
FE05
FB13
FA57
FAF9
FB51
FAE0
FA82
FAEC
FBAF
FBF4
FB97
FB2C
FB1F
FB3C
FB22
FAE1
FAD4
FB1B
FB75
FB9C
FB90
FB7C
FB74
FB65
FB34
FAF1
FAD5
FB07
FB55
FB6E
FB44
FB19
FB06
FAE8
FADA
FB93
FDC0
010D
041D
05B6
05CD
0549
04E7
04B2
0476
0449
045B
0498
04CC
04F0
0512
0515
04E2
04A5
049D
04C1
04C6
0492
0465
0482
04D6
050F
0504
04D3
04AB
04A2
04BB
04DA
04B9
044C
0423
04B5
053C
0401
006D
FC3D
F9FB
FA4D
FB7D
FBBB
FB18
FACD
FB37
FB7F
FB29
FAE3
FB51
FBEE
FBD7
FB26
FABA
FAEB
FB3D
FB4D
FB54
FB91
FBC7
FB99
FB28
FAE3
FAE2
FAED
FB07
FB62
FBB7
FB74
FAE8
FB80
FE23
01C2
0456
050E
04DC
04DF
051E
0504
049E
048C
04F7
0543
0502
0490
0473
0495
0497
047E
048E
04B8
04B5
0499
04B6
04FE
04F9
0487
0438
048E
0520
0515
0471
0436
04E7
0567
0406
0091
FCC7
FAA1
FA7A
FB1E
FB55
FAFD
FAB6
FADE
FB2F
FB3E
FB12
FB03
FB36
FB75
FB82
FB62
FB45
FB42
FB4A
FB54
FB64
FB82
FB9A
FB83
FB2A
FAB4
FA78
FAC4
FB7E
FBF7
FB87
FA98
FAD0
FD7B
01BA
04F8
0590
047E
03F1
04AA
0576
0531
045E
0439
04E3
0552
04F1
0462
045A
049D
049D
0476
0497
04E3
04E4
04A3
04A4
0504
0548
0525
04F7
050E
050F
0498
0435
04A7
053B
0407
006C
FC60
FA5E
FAA6
FB6F
FB71
FB18
FB2C
FB6F
FB38
FABB
FAC9
FB6C
FBC4
FB6A
FB13
FB62
FBDB
FBBD
FB3B
FB0D
FB35
FB21
FAC6
FABF
FB34
FB70
FB04
FAA6
FB2D
FC04
FBC3
FA81
FA62
FD15
0174
04A8
0551
04A5
0475
0512
058F
0564
050B
050E
0541
052A
04C1
046B
0460
047E
04A1
04C1
04CE
04B5
048B
0489
04B4
04D7
04D6
04DD
0507
0519
04CB
0464
0492
0565
05BB
0423
0095
FCCB
FAB1
FA90
FB1F
FB36
FAE8
FADB
FB24
FB41
FB01
FAD6
FB12
FB57
FB2A
FACA
FADE
FB6F
FBC4
FB71
FAF2
FAE7
FB35
FB5C
FB44
FB37
FB3E
FB1B
FAE0
FAFB
FB65
FB6C
FAE2
FB0F
FD75
018E
04D4
0588
04A1
043B
04E9
0578
0516
0471
0478
04EF
04FA
0493
0484
0505
054E
04D9
0442
0458
04F3
055A
0559
0540
051A
04B9
045E
0491
0532
0561
04BF
0437
04B5
055C
0425
0085
FC85
FA87
FAAB
FB37
FB0F
FABA
FAF7
FB7C
FB8B
FB28
FB02
FB4F
FB88
FB4D
FAFD
FB0B
FB43
FB36
FAFB
FAFA
FB33
FB45
FB12
FAEA
FAEF
FAE0
FAA7
FAB3
FB4E
FBDD
FB7B
FA7E
FAA4
FD3D
0162
04A9
059B
04F6
046A
04A5
050F
050C
04D6
04EA
0530
0530
04D2
0482
048C
04B5
04A8
0474
0468
0499
04D4
04FC
051C
052A
050A
04E0
04FD
054F
054A
04BD
045A
04D2
0570
045F
00D8
FC93
FA3C
FA98
FBDE
FC15
FB3E
FAAD
FAF0
FB56
FB37
FAE0
FAE3
FB31
FB5A
FB52
FB68
FB97
FB84
FB2F
FB15
FB5D
FB7C
FB19
FAAD
FAC9
FB2A
FB2A
FAE0
FAF8
FB73
FB6F
FAB6
FABB
FD22
0159
04BE
0588
04A5
0426
04A7
0521
04DA
045C
0463
04C6
04E8
04C1
04C2
04FC
0509
04D3
04CC
0516
0530
04C6
045F
0491
0509
0509
049B
047F
04E0
04F8
0459
03E5
0498
059E
04BF
011D
FCAC
FA36
FA64
FB78
FBBC
FB36
FAE7
FB2F
FB91
FBA9
FB9C
FB94
FB6B
FB15
FAE1
FAF9
FB09
FAC6
FA83
FAC4
FB5D
FB9C
FB47
FAFB
FB41
FBBD
FBC7
FB7D
FB88
FBE0
FBB3
FAE8
FAFC
FD71
0198
04E3
0592
047D
03C7
044C
051D
0531
04B9
047C
049F
04B9
04AA
04B5
04E1
04E5
04B6
04B2
0501
053C
0508
04AC
04AA
04DF
04B4
042B
03F9
045E
049D
042C
03C5
0457
0533
0450
00DB
FCAE
FA7A
FACE
FBC4
FBA8
FAD1
FA8C
FB10
FB7A
FB52
FB15
FB3B
FB82
FB87
FB6B
FB76
FB7A
FB1E
FAA3
FAB2
FB50
FBAC
FB53
FAE0
FB0E
FB9B
FBCC
FBAB
FBE0
FC58
FC19
FAEB
FA6F
FC8C
00DE
04B1
05E4
0514
0463
04C6
0566
055A
04E1
04B7
04E5
04E8
049E
046C
048D
04B8
04B5
04AF
04C8
04C6
048B
047B
04E7
0563
0543
049D
0437
0464
0482
0418
03CC
0473
054C
0452
00C5
FC92
FA6D
FADA
FBF2
FBEA
FAF7
FA6A
FAB1
FB16
FB0A
FAE0
FB06
FB47
FB45
FB27
FB42
FB6E
FB45
FAE3
FAD4
FB3C
FB97
FB83
FB53
FB73
FBA2
FB5C
FADB
FAEA
FB8D
FBC0
FB0B
FAC9
FCCB
00E6
04B4
0616
0560
0487
04AE
053A
053A
04CE
04B1
0502
0537
050A
04D1
04E3
0521
0545
0546
0537
0505
04A4
0454
0462
04AF
04CF
04AE
04AA
04E1
04E8
0487
0458
04F0
0592
0485
011A
FCE9
FA67
FA5F
FB5B
FB9E
FAFF
FA7A
FA92
FAD5
FAD1
FABB
FAE8
FB29
FB18
FAC1
FA97
FAC1
FAF2
FAFA
FB0E
FB4C
FB6B
FB3B
FB12
FB50
FBB4
FBAE
FB44
FB18
FB59
FB54
FAAF
FA96
FCB5
00E5
04BE
060C
0533
0461
04D8
05CA
05F1
054C
04D1
04ED
0526
0516
0503
0538
0567
052D
04C7
04BA
050B
0541
0519
04BF
0466
041A
03FD
0450
04F4
0547
04EC
047E
04C3
0533
0426
00E7
FCF5
FA96
FA61
FAFB
FB01
FA7F
FA46
FA86
FABC
FAAB
FAB4
FB15
FB75
FB77
FB4A
FB3E
FB35
FAF2
FAB1
FAE0
FB5E
FB8B
FB36
FAF2
FB37
FBA5
FB9D
FB4F
FB71
FBF0
FBD2
FAD6
FA8A
FCC1
0120
050C
065E
0584
049F
04E5
05AA
05CE
0547
04DA
04DA
04EB
04C3
0495
04A3
04CC
04CB
04A9
0498
049F
049D
049A
04BC
04F1
04F4
04BF
049D
04A8
0495
0445
0435
04BE
0518
03C9
0075
FCBA
FAAF
FAAF
FB3C
FB0C
FA6F
FA55
FACB
FB14
FAEF
FADE
FB38
FB90
FB73
FB25
FB30
FB7F
FB87
FB3F
FB33
FB86
FB9C
FB20
FAB1
FAF6
FB84
FB85
FB19
FB32
FBF5
FC3E
FB6C
FAEA
FCD0
0106
04E4
0624
054B
047C
04B7
053D
0540
0502
0504
0513
04BE
0441
0445
04C9
0511
04C5
046D
048D
04DE
04E3
04BD
04CA
04E8
04BA
0475
04A0
0517
0502
0433
03C8
04A9
05BA
04B4
00FD
FCC0
FA8A
FA8E
FB08
FAD3
FA82
FAE4
FB9B
FBB9
FB32
FADA
FB13
FB5A
FB3B
FB0D
FB46
FBAA
FBB5
FB77
FB6B
FB96
FB7E
FB07
FAC2
FB0C
FB66
FB31
FABA
FAD3
FB70
FB8A
FAD4
FABD
FCEC
00FA
048A
05CC
0538
0487
048F
04CD
04BC
04A7
04FA
0567
0562
04F9
04AB
04A0
0487
0448
0435
0480
04D8
04ED
04EB
051F
0554
051E
04B0
04B2
051A
0502
041A
0385
0465
05CB
0546
01CC
FD54
FACB
FAE1
FBB3
FB89
FABC
FA94
FB34
FBA5
FB6A
FB0A
FB0C
FB34
FB1C
FAEB
FB01
FB3F
FB37
FAF2
FAF4
FB53
FB7F
FB23
FAC7
FB05
FB9B
FBD4
FB9C
FB75
FB7C
FB30
FA89
FAA7
FCBA
0059
039E
0514
0502
049F
0491
04AE
04C5
04EA
0516
050F
04DA
04D2
0514
0539
04E5
0469
045D
04B8
04DE
049D
0487
04FF
0575
0532
047E
0451
04E4
0558
0510
04AE
0513
05A5
0498
012D
FD06
FA8C
FA6F
FB47
FB8B
FB20
FADB
FB20
FB85
FB9C
FB7D
FB6D
FB69
FB54
FB44
FB5B
FB70
FB46
FAF8
FAE5
FB25
FB58
FB2A
FAD0
FAC8
FB2F
FB86
FB4C
FAAD
FA80
FB9D
FE2C
0170
0432
058C
0590
0517
04E9
050C
050D
04BF
0478
0488
04C0
04BC
0478
044C
045D
046D
0458
045D
04B0
0506
04F0
048E
0479
04E0
0538
050D
04C4
0503
0560
046C
016C
FD92
FAFE
FA8F
FB3F
FB96
FB44
FAF8
FB23
FB6F
FB75
FB59
FB6C
FB91
FB6E
FB0E
FAE7
FB30
FB8D
FB8E
FB47
FB2A
FB5B
FB7D
FB42
FAE5
FADD
FB2D
FB48
FADB
FA83
FB78
FE4C
0214
04F8
05CC
051A
0473
04B9
0564
0573
04C0
0417
041D
048C
04B9
048B
0476
04B6
04FB
04F9
04DB
04DB
04CE
0473
040E
0428
04B4
04F5
0490
0441
04E3
05DD
0554
0248
FE0E
FB20
FA91
FB40
FB7E
FAEB
FA5F
FA7C
FAF1
FB25
FB0E
FB02
FB15
FB0F
FAF2
FB07
FB65
FBAE
FB87
FB21
FB07
FB67
FBCE
FBB9
FB49
FB1C
FB76
FBCF
FB80
FACF
FB02
FD26
00C8
040F
056D
0506
0455
0479
0536
059D
055F
0505
0507
0530
0515
04D3
04D9
0529
053C
04CC
0446
0432
0470
0483
0468
049C
0530
0566
04B8
03DD
040A
051C
053C
02DC
FEC5
FB7D
FA9E
FB5C
FBCF
FB34
FA63
FA4F
FAD4
FB31
FB28
FB16
FB2D
FB27
FAD8
FA93
FAB6
FB1D
FB57
FB52
FB6D
FBCF
FC05
FB9A
FAD9
FA93
FB0E
FB98
FB6C
FADB
FB3C
FD7F
0107
0414
0565
0541
04DA
04EE
053A
052E
04CB
0498
04D8
052D
0525
04DD
04D5
0529
056A
0539
04D0
04A3
04B4
049F
044D
042A
0484
04F5
04EB
0491
04A4
052F
04F5
02B2
FED8
FB7D
FA44
FACB
FB5E
FB08
FA65
FA6D
FB14
FB7B
FB30
FAAA
FA80
FAA6
FABA
FAAC
FAC1
FB08
FB33
FB23
FB28
FB82
FBD7
FB9F
FB06
FAD9
FB6C
FBF1
FB6F
FA4D
FA52
FCCE
00F0
0469
05A9
052C
0491
04C5
055D
058F
0546
0505
0517
0541
053B
051D
0529
0555
0553
050C
04C0
04AA
04B0
0497
0473
0493
04FC
0533
04DC
045E
0479
0529
0535
0350
FFAC
FC1A
FA5E
FA8B
FB3A
FB37
FAA1
FA4D
FA88
FAD3
FAC8
FAA7
FADE
FB4D
FB6A
FB11
FAC1
FAE6
FB49
FB65
FB28
FAFB
FB14
FB2D
FB05
FADE
FB12
FB62
FB31
FA98
FAD0
FCFC
00AE
0402
0574
053E
04C9
0501
058F
05B6
055F
050D
050B
0515
04DF
048F
0479
04A5
04D0
04DB
04EC
051A
052B
04F0
04A5
04B9
0527
055C
04F9
0478
04AE
058B
05B1
03B1
FFBF
FBD3
F9EC
FA39
FB34
FB65
FAC3
FA49
FA84
FB0A
FB36
FB0C
FB0A
FB5A
FB96
FB70
FB20
FB0B
FB2C
FB30
FB08
FB02
FB45
FB7E
FB59
FB14
FB23
FB68
FB36
FA76
FA4F
FC27
FFEA
03BB
05B2
059D
04E0
04B7
0519
0549
050F
04E1
050B
053D
050E
04A0
046A
048F
04B4
0492
0466
0490
04FB
052E
04F4
04A4
049E
04C2
04B3
0480
04A8
0544
0567
03D5
0074
FCC2
FA94
FA61
FB0D
FB4D
FAF1
FAAB
FAE4
FB38
FB28
FAD7
FACB
FB22
FB75
FB76
FB5C
FB75
FB9F
FB7F
FB29
FB18
FB70
FBAB
FB4C
FAB1
FAAA
FB4A
FBAA
FB37
FADD
FC40
FFB3
037D
0578
053B
0449
042F
04F2
0580
0541
04B3
048A
04C8
04F0
04D2
04C0
04F4
0530
0516
04B2
0469
046C
048D
049C
04B3
04EB
0509
04C0
0444
0437
04C6
0501
0398
005A
FCC2
FAAF
FAA0
FB69
FBA8
FB2E
FACC
FB08
FB76
FB6F
FAFE
FAC2
FB01
FB4B
FB26
FAC4
FABA
FB33
FBB3
FBBC
FB65
FB1C
FB0D
FB13
FB27
FB7A
FBF3
FC07
FB67
FAD9
FBCB
FED8
02D7
05BB
066F
05A2
04BE
047A
048D
0487
0470
0486
04BD
04D4
04C3
04C5
04EA
04F5
04C3
049B
04CD
0529
0529
04AF
0447
046E
04D2
04B8
0415
03C4
0459
04FF
0415
0102
FD26
FA9D
FA3D
FB03
FB74
FB29
FACF
FAFA
FB71
FBA8
FB85
FB5F
FB60
FB4D
FAFB
FAAB
FAC5
FB3B
FB8E
FB6D
FB23
FB2A
FB82
FBBF
FBB0
FBA2
FBD1
FBE4
FB6A
FAE5
FBB8
FEB5
02C3
059D
0604
04E9
0432
04A5
056C
057F
04F6
049E
04BA
04CF
048E
0459
049C
050B
0507
0492
044C
0483
04BE
0483
042B
046B
0529
056E
04C1
03F9
042A
04EA
0472
01A4
FD8E
FA81
F9C2
FA8B
FB44
FB37
FADC
FAC8
FAF2
FB09
FB0F
FB46
FBAA
FBD7
FB87
FB03
FAD6
FB2B
FB9D
FBBD
FB8D
FB5B
FB46
FB29
FB00
FB0E
FB74
FBC4
FB76
FAE8
FB7D
FE3C
0251
0581
0649
054F
0470
04A2
053F
0552
04E9
04BC
04F4
0500
049E
0458
04A7
0518
04EC
0448
0419
04BB
055F
0528
0476
045C
04FE
054D
049E
03D1
0427
0534
04F5
0229
FE07
FB0C
FA63
FB01
FB45
FAD7
FA8A
FADF
FB61
FB70
FB21
FB00
FB3A
FB74
FB5D
FB23
FB1C
FB44
FB4D
FB25
FB19
FB4F
FB78
FB34
FABA
FAB3
FB55
FBE8
FB9B
FAD4
FB2D
FDC5
01B4
04B9
0579
04C2
045B
04EA
058E
0567
04CC
04A8
0512
053E
04C7
044F
048B
0529
0541
04AE
0445
0499
051E
04FD
045C
0431
04C8
0543
04E6
044B
0493
0586
054F
0292
FE48
FAF7
FA1A
FADE
FB73
FB25
FAAB
FAC4
FB30
FB4B
FB09
FAEC
FB24
FB46
FAFE
FAA3
FAC9
FB5B
FBB1
FB75
FB1F
FB3F
FB9C
FB88
FAF6
FAB3
FB3E
FBDD
FB75
FA53
FA61
FD19
018D
0513
05FD
052C
04AB
0539
05CF
0564
0463
0402
049B
0552
055E
0501
04F0
0536
053C
04C8
0462
048B
0501
0523
04E4
04CC
050D
0518
047A
03C8
040A
0523
0558
0307
FEA9
FAB8
F952
FA42
FB94
FBCE
FB32
FAD2
FB0A
FB46
FB16
FAC7
FAD2
FB18
FB19
FABD
FA7D
FAA5
FAE5
FAD8
FAAB
FAD9
FB53
FB81
FB2C
FAFB
FB85
FC49
FC2A
FB21
FAD7
FCF4
010B
04BE
0618
0568
0477
046A
04DE
0507
04E6
0504
0576
05AD
055C
04F5
050A
0571
0587
0521
04CD
04F8
054E
0532
04B3
0476
04BE
04F1
0481
03DF
0405
04EB
0512
030C
FF4C
FBEA
FA88
FAD6
FB4D
FB10
FA84
FA5A
FA89
FAA1
FA97
FAC3
FB28
FB44
FADC
FA72
FAA4
FB41
FB7D
FB05
FA72
FA77
FAED
FB28
FB01
FB16
FBC9
FC74
FC26
FB15
FACC
FCAF
0062
03F8
05B4
0588
04D1
04C4
055B
05BF
057A
04F3
04CB
050E
0539
0503
04BA
04C1
04FA
04FD
04C9
04C9
0523
0562
051E
04A4
048A
04C6
04B5
0436
0413
04C9
0546
03B7
FFD8
FBBA
F9BC
FA21
FB31
FB6F
FAFF
FAC7
FAF8
FB0E
FAD6
FABE
FB0B
FB5E
FB58
FB29
FB28
FB39
FB11
FADB
FB00
FB74
FBAB
FB77
FB4E
FB7B
FB7A
FAE0
FA9C
FC57
0042
044A
0624
05B4
04CF
04D4
0560
0573
0500
04BF
04F2
0514
04DD
04B5
04F5
0542
051C
04AC
0476
0492
04AB
04AC
04C6
04E3
04A6
0435
045C
054C
0598
0375
FF28
FB41
F9F1
FABF
FB86
FB2F
FA87
FA91
FB12
FB38
FAF7
FAF8
FB5B
FB7F
FB14
FAA9
FAC9
FB2C
FB45
FB25
FB32
FB5C
FB47
FB19
FB58
FBD8
FBA4
FA8E
FA39
FC8B
010E
04F6
0621
0547
0497
04EA
0550
0505
048D
04A5
04FE
04D9
045A
0455
04EF
054D
04ED
0470
0490
04FA
04F3
049A
04A7
0519
0524
049B
0472
052D
056C
033E
FEDC
FAF5
F9C4
FAAC
FB74
FB1F
FA9A
FAD6
FB68
FB74
FB0B
FAEC
FB47
FB84
FB4E
FB0C
FB1C
FB43
FB40
FB52
FBB2
FBF2
FB93
FAF9
FAF6
FB77
FB7C
FABD
FAB5
FD0E
0147
04D5
05E5
0532
04A6
04F2
054B
0514
04B5
04BA
04ED
04D4
048D
0493
04DE
04E6
048F
045C
0490
04B5
0475
0437
0476
04CD
0491
041B
0475
058D
0581
02AE
FE10
FA9B
FA06
FB1C
FBA0
FB02
FA78
FAD6
FB83
FB98
FB2D
FAF8
FB28
FB4D
FB2D
FB18
FB46
FB74
FB6A
FB5D
FB80
FB95
FB60
FB3B
FB8C
FBEE
FB97
FAC9
FB1F
FDCE
01E7
0505
05CB
0518
0495
04CA
051F
0521
0504
04FF
04E5
049C
046C
048C
04B4
0488
0444
046E
04F1
0523
04D2
0499
04DF
0515
049E
0405
0456
053F
04CD
01B7
FD4C
FA58
FA1E
FB3A
FBAF
FB27
FAA4
FAB8
FAF4
FAED
FAE4
FB23
FB63
FB45
FB0D
FB43
FBD2
FC11
FBB6
FB3D
FB11
FAFF
FAC7
FAC1
FB3F
FBB5
FB5C
FAB5
FB7E
FEAD
02DC
0588
05C1
04EC
04BB
053D
0568
04E5
0469
0488
04F8
052A
0514
0500
04F7
04CD
0493
048B
04AB
04A1
0474
048C
04F0
050C
049D
0458
04E1
0570
0449
00E5
FCF1
FAA6
FA6F
FAE4
FAD8
FA95
FACD
FB4D
FB61
FB0C
FAF1
FB3F
FB63
FB0B
FAB5
FAE8
FB5B
FB68
FB1E
FB22
FB8B
FBB4
FB59
FB2A
FB9C
FBEB
FB31
FA3D
FB32
FEE4
036A
05FD
05F2
0500
04D3
0548
0564
0507
04D8
0507
0515
04CF
04AB
04EF
0520
04C1
0431
042C
04B1
04FC
04B3
045F
0473
049A
047B
0489
0537
05A5
0423
005D
FC4C
FA4A
FA93
FB59
FB2E
FA80
FA6E
FB06
FB63
FB21
FAC9
FAE0
FB37
FB64
FB5C
FB52
FB4C
FB32
FB27
FB58
FB8C
FB60
FB05
FB21
FBAF
FBC0
FAE4
FA61
FC12
0001
03F0
05AE
0554
04B8
04FB
0583
055F
04C6
0491
04EE
0541
052A
04EB
04CB
04AD
0477
0463
0499
04C5
048D
0440
0470
04ED
04E4
043E
0416
0518
05F0
046A
0038
FBBF
F9A9
FA2A
FB43
FB5B
FAC3
FA94
FAF8
FB40
FB18
FAE0
FAE9
FB0A
FB12
FB23
FB60
FB9A
FB97
FB7C
FB8A
FBA2
FB79
FB3E
FB70
FBEA
FBCF
FAE6
FA89
FC68
0057
0416
05A6
0543
04AF
04EB
0561
0546
04D1
04B7
0502
0522
04ED
04D4
0510
053E
04F7
0477
0440
045D
0471
045D
045A
0477
046F
044E
0494
0549
0546
0340
FF79
FBE1
FA39
FA6C
FB0F
FB23
FADA
FAC1
FAE1
FAFF
FB20
FB5C
FB7A
FB36
FACB
FABB
FB19
FB71
FB7B
FB7A
FBB0
FBD2
FB8A
FB36
FB70
FBF0
FBAD
FA94
FA5B
FCBB
0119
04D2
05F9
0535
0485
04D4
0563
055E
04FC
04D3
04E0
04C8
049F
04BE
050C
0512
04C5
049D
04CD
04EA
04A5
0465
049F
04EE
0493
03E1
0413
054A
059B
031C
FE86
FAD1
F9FA
FB0E
FBBA
FB28
FA70
FA97
FB39
FB6E
FB2B
FB09
FB2D
FB3F
FB23
FB22
FB4E
FB58
FB27
FB16
FB52
FB74
FB2B
FAF2
FB68
FC0F
FBBA
FA87
FA7B
FD44
01DB
0553
0602
0502
0468
04CE
053C
04FD
0482
046B
049F
04BB
04D0
050C
0527
04D4
046C
0489
0507
052B
04C7
0494
04FE
0549
04A2
03B7
03FE
0549
0549
0249
FDAA
FA88
FA3C
FB3F
FB8A
FAF4
FAAB
FB1C
FB82
FB5B
FB23
FB54
FB89
FB40
FAD6
FAEF
FB5C
FB68
FB07
FAE8
FB46
FB75
FB10
FACF
FB70
FC38
FBCB
FA87
FAC5
FE08
02B0
05A7
05D1
04D9
04A7
0537
056C
0506
04C5
04F7
04FE
0484
0428
0477
04F8
04F6
04A8
04C0
0526
0516
047A
0436
04BA
052C
04AC
03F4
046C
05AD
0545
01BE
FCDF
F9EB
F9FD
FB41
FB9F
FB03
FAA2
FAE9
FB32
FB1D
FB1B
FB6F
FB98
FB2F
FABC
FAEF
FB89
FBC0
FB71
FB36
FB4D
FB41
FAE4
FAD1
FB6B
FBE0
FB31
FA23
FAF2
FE96
0326
05CF
05DB
0501
04DF
0550
055A
04E1
0498
04C5
04EB
04C7
04BD
0502
051F
04B8
044C
047C
04FE
0502
0482
0451
04C3
0516
04B0
044C
04EE
05DE
04EC
0130
FCA1
FA1A
FA3B
FB2F
FB41
FAA9
FA87
FB11
FB7D
FB61
FB28
FB3A
FB59
FB3C
FB21
FB4A
FB6B
FB2B
FADC
FB10
FB96
FBAB
FB33
FB07
FB99
FC01
FB44
FA42
FB3C
FF01
037A
05D8
059C
04A7
0496
051E
0530
04C2
04A0
0500
0536
04E5
0496
04C9
051D
04F8
048E
0485
04E4
0510
04CE
0491
049C
0482
0404
03D2
049E
057F
046A
00B3
FC61
FA28
FA87
FBA5
FBC7
FB14
FAAC
FAF0
FB4C
FB4D
FB27
FB14
FAF0
FAB8
FAC6
FB2F
FB6A
FB14
FAAD
FAE7
FB89
FBB9
FB5A
FB49
FBF1
FC5B
FB9B
FAB5
FBEB
FFCC
03FE
05CA
051C
0428
046F
0544
055D
04C2
0479
04D4
0520
04E3
0497
04C0
0519
0525
0506
051D
0542
0507
0494
047D
04C0
04A8
0404
03BC
0477
0512
038A
FFA9
FBC0
FA20
FAA6
FB65
FB45
FAE5
FB0F
FB7A
FB7B
FB30
FB2E
FB6A
FB47
FAC0
FA99
FB17
FB77
FB1E
FAA1
FADF
FB85
FB8B
FAE8
FABF
FB91
FC43
FBD3
FB56
FCFC
00FB
04C6
05F7
0507
043C
0499
0519
04C1
0425
044A
0504
054E
04E9
04A1
04EC
0540
051A
04DB
0508
0547
04FB
0468
0458
04C5
04CD
0431
03EB
0498
04EE
02F9
FEE2
FB42
FA3F
FB2E
FBDD
FB73
FAED
FB22
FB85
FB43
FAA5
FA8F
FB0E
FB4C
FAEB
FA92
FACC
FB38
FB42
FB21
FB58
FBC0
FBC6
FB7F
FB96
FC0A
FBEC
FAE8
FA77
FC7E
00C0
04A1
05F5
0532
046C
04AA
053A
0548
050B
051C
0560
054C
04DF
04A5
04D3
04F7
04C2
0484
0492
04A9
046E
042A
045B
04D0
04D7
0470
0478
053C
0561
032C
FEE0
FB04
F9CC
FAC8
FBB5
FB49
FA51
FA2C
FAE8
FB77
FB45
FADE
FAFD
FB7F
FBB8
FB74
FB2F
FB50
FB97
FB88
FB27
FAFC
FB4F
FBB1
FB75
FABE
FACB
FCDA
00AF
0476
064F
060B
051A
04E5
0567
05A2
051E
0471
0451
04A3
04CC
04A6
0496
04C3
04C6
045C
0403
0464
0541
0595
04EA
0425
0468
0556
0522
0284
FE64
FB13
FA06
FAA0
FB3E
FB16
FAA9
FAB1
FB23
FB70
FB5F
FB42
FB57
FB66
FB27
FAD2
FAED
FB86
FBF6
FBA8
FAE6
FA97
FB0E
FB90
FB45
FA8D
FAF7
FD9D
01B3
0509
0617
0556
047E
049D
0540
0562
04D5
0459
0483
04F9
0508
04A5
046F
04C0
0525
0504
0488
0466
04CF
0518
04BA
043D
048D
056B
052B
0281
FE46
FAEA
FA03
FADD
FB9A
FB59
FACF
FAE2
FB6C
FBA1
FB3E
FAD4
FAE2
FB2E
FB38
FB00
FAF3
FB3A
FB73
FB4A
FB05
FB2F
FBC4
FC0B
FB7C
FAB1
FB21
FDB0
0190
04C6
05E3
053B
0459
0457
04ED
052B
04C4
045D
048D
0517
0555
051F
04E9
04FF
0515
04D0
0471
047C
04E7
0501
0479
03FA
0451
0512
04A3
01F5
FDEF
FAC7
F9EF
FAD6
FBC5
FBB4
FB0A
FAB6
FAFC
FB59
FB54
FB0E
FAF6
FB25
FB42
FB13
FAD5
FAE1
FB26
FB47
FB33
FB50
FBCC
FC1C
FBA1
FACD
FB35
FDF8
0231
057E
0647
0536
043E
046F
052D
056C
050F
04C5
04ED
051F
04EC
048E
0489
04DF
0513
04E9
04B6
04D5
0509
04CE
0434
03FB
049A
054D
048D
019F
FD9B
FA96
F9C6
FA8B
FB51
FB3B
FAC2
FABF
FB3B
FB7F
FB27
FAAC
FAB9
FB3C
FB89
FB43
FADB
FADF
FB37
FB5B
FB2A
FB20
FB7D
FBC2
FB5E
FAD5
FB90
FE5B
0239
0523
05F2
0555
04D0
0513
058D
0575
04D8
046B
0498
0506
0525
04E7
04B7
04D6
0508
04FD
04D1
04DA
0511
0508
049D
045E
04D4
056B
049B
0189
FD58
FA58
F9CB
FAC2
FB67
FB03
FA6C
FA8D
FB2D
FB6E
FB17
FACF
FB16
FB8B
FB8C
FB23
FAEB
FB20
FB43
FAEF
FA88
FABB
FB69
FB9B
FAD7
FA27
FB48
FEC2
0308
05D4
063A
0543
0496
04CC
053E
0532
04CC
04AD
04FD
0534
04E4
045B
0436
048E
04D6
04AF
046F
04A3
052B
0553
04E2
0496
051E
05CB
04DD
0176
FCF5
F9E9
F998
FAE2
FBBD
FB5E
FAA4
FA9A
FB21
FB65
FB1E
FAE2
FB2D
FBAC
FBC1
FB71
FB50
FB99
FBC8
FB66
FAD6
FADE
FB77
FBA4
FAD3
FA0B
FB26
FEB5
030C
05BF
05F6
04F6
047A
04E5
055A
0527
04A0
0477
04BF
04EE
04B3
045E
0459
048B
048F
045B
0454
04A4
04DF
0490
040B
042F
0530
05DD
0495
0119
FD15
FAAA
FA72
FB30
FB6C
FAF3
FAA3
FB02
FB8F
FB8D
FB14
FAE8
FB5A
FBDA
FBC2
FB48
FB2E
FBA7
FC06
FBB2
FB15
FB16
FBC5
FC1B
FB63
FA8B
FB74
FECF
0308
05A9
05C6
04A7
0424
04B3
0556
0530
048C
0447
0498
04E9
04C4
0470
0470
04AF
04A5
0432
03E4
0436
04C8
04D0
0443
0402
049D
0532
0414
00B9
FCAA
FA2B
FA11
FB27
FBB7
FB52
FAD1
FAF5
FB7C
FBB3
FB7A
FB54
FB85
FBAC
FB5F
FAE9
FAF6
FB9F
FC24
FBE9
FB51
FB3E
FBC2
FBED
FB33
FAA0
FC06
FFCC
040D
0650
0601
04C5
0466
04FC
0559
04E0
0438
0438
04B1
04CD
0459
0410
047E
052B
0536
048E
0409
0435
049B
0476
03ED
03F1
04D0
0556
03D4
0017
FBF1
F9A1
F9C2
FAFB
FB9C
FB3B
FAB0
FAC6
FB54
FBAE
FB91
FB59
FB5E
FB7B
FB6A
FB3E
FB49
FB86
FB8F
FB3D
FB0F
FB8B
FC55
FC67
FB77
FAD2
FC3A
FFE9
0400
063A
0619
050B
04A3
0503
0542
04E2
0461
0465
04CB
04EE
049B
0451
047F
04DF
04DB
046E
042F
047E
04E5
04B8
0416
03DA
0469
04C8
0374
001C
FC4E
FA0E
F9EF
FAC7
FB33
FAFC
FAE1
FB49
FBB4
FB8A
FAFE
FAC6
FB1F
FB83
FB76
FB31
FB45
FBBA
FBFC
FBB4
FB50
FB63
FBC6
FBBC
FB23
FB10
FCD1
005C
0407
0600
05F3
0515
04B0
04E9
050D
04B3
0441
044F
04CD
0527
0505
04B1
0491
049A
0475
0425
0415
0474
04CB
0498
041F
0434
04F3
051F
0347
FF88
FBC9
F9F7
FA38
FB18
FB4E
FAED
FACC
FB32
FB98
FB83
FB2C
FB15
FB4F
FB78
FB61
FB57
FBA2
FC06
FC06
FB97
FB44
FB78
FBDC
FBB8
FB06
FADE
FC85
FFFB
03AD
05C6
05D1
04F0
048B
04F2
056A
0550
04D1
047C
047C
0481
045F
0455
0491
04CA
0497
0415
03DA
042C
0495
048C
0443
0473
052C
0548
0371
FFC2
FC05
FA21
FA5E
FB5E
FBAA
FB14
FA7C
FA91
FB1A
FB76
FB7B
FB7E
FBB4
FBDA
FBA7
FB50
FB4B
FBAA
FBF4
FBD0
FB86
FB87
FBAB
FB56
FA96
FAA3
FCC1
009E
043A
05C2
0547
0464
045C
04F5
053E
04F5
04B4
04E8
052F
04F9
0462
040D
043C
047B
0458
0415
0445
04DA
0514
048A
03EC
0438
0545
0578
035F
FF6E
FBC8
FA3E
FAAD
FB81
FB8F
FB15
FAF4
FB59
FBA4
FB59
FAD2
FABC
FB35
FBBA
FBE1
FBCC
FBC4
FBB5
FB5D
FAE5
FADC
FB73
FBFF
FBB1
FAC5
FAAD
FCB4
007C
041D
05D5
058D
049E
044B
04A7
04F4
04C3
0467
045F
04A6
04D3
04B8
0495
04A1
04B2
0486
0447
045F
04D4
0517
04C5
0457
049B
0566
0546
02EC
FEE4
FB5B
FA15
FAC8
FBBA
FBBD
FB29
FAEB
FB3A
FB8C
FB8D
FB82
FBAC
FBC3
FB68
FADC
FACB
FB5C
FBE0
FBAA
FB02
FACB
FB48
FBB2
FB43
FA73
FACB
FD4D
013C
049A
05E9
055F
0469
0431
04AF
0516
04E7
0470
0444
047B
04AA
048C
045D
047B
04D0
04F9
04D7
04BA
04D5
04E2
0496
044A
04A3
0569
0535
02C8
FEB4
FB28
F9E2
FA8E
FB77
FB7C
FB02
FAF5
FB6E
FBC3
FB94
FB46
FB55
FB9B
FB9D
FB48
FB0E
FB36
FB6C
FB41
FAE4
FAF1
FB88
FBEA
FB61
FA6B
FAA0
FD21
013E
04DA
0647
05B1
04A4
0460
04D7
0536
0508
049B
0466
0476
048A
0488
0497
04C2
04D3
04AB
0483
04A2
04E8
04EA
0495
0472
04F1
0588
04E4
0240
FE72
FB5F
FA42
FAAB
FB3C
FB2F
FADD
FAEA
FB51
FB88
FB56
FB1D
FB42
FB95
FBA1
FB58
FB21
FB31
FB3D
FB03
FAD5
FB34
FBF3
FC29
FB58
FA66
FB00
FDE4
01EC
0503
05F8
0555
0480
0459
04B6
04F9
04E4
04BD
04CD
04F9
04F1
04A8
046F
0486
04CC
04EF
04E1
04DF
04F9
04E5
0482
044C
04CB
057F
04DB
01E7
FDAA
FA80
F9DA
FAEE
FBE1
FBD0
FB4E
FB21
FB3A
FB29
FAFD
FB17
FB68
FB71
FB19
FAEE
FB4C
FBB2
FB73
FAD1
FAB7
FB51
FBA7
FB13
FAA9
FC3F
000F
0406
05E1
0586
04BE
04DE
0577
0570
04B6
042E
0456
04B6
04BB
048F
04A6
04EE
04EE
049D
047B
04BF
04EF
04A8
045F
04B6
052D
0445
0147
FD78
FAF2
FA75
FAE3
FAF3
FAAD
FAD7
FB77
FBB9
FB3B
FAB4
FAED
FB9D
FBD7
FB66
FB06
FB33
FB76
FB41
FAEA
FB1F
FBA1
FB7A
FAA6
FAC5
FD5A
01A3
0508
05D5
04E9
044E
04C9
056B
0546
04A7
0461
0498
04D0
04D2
04DE
04FD
04CE
0441
03F8
046A
050E
0500
046A
0471
056C
05D9
03D5
FF95
FB90
F9FE
FAA4
FB8C
FB7A
FAEE
FADD
FB42
FB6B
FB30
FB15
FB5C
FB8C
FB3D
FAD0
FAE9
FB6E
FBA8
FB5B
FB28
FB79
FBB9
FB2D
FA7A
FB6A
FEC8
0306
05A0
05B2
04A7
0448
04CA
0527
04DE
048B
04C1
0527
0513
049B
0468
04AB
04E0
04B0
0480
04B7
04FD
04BA
0435
0457
051B
04EF
0263
FE35
FAE4
FA1E
FB1D
FBDC
FB79
FAC5
FABA
FB33
FB6C
FB2E
FAEC
FAF0
FB08
FB0D
FB2E
FB81
FBB0
FB75
FB24
FB43
FBA8
FB8A
FACC
FAAE
FC9B
0056
03E8
058D
055D
04CF
04E0
0540
0538
04C9
048A
04BA
04FC
04F8
04DC
04F5
0525
0514
04C0
0485
0488
047A
0435
0427
04B7
0542
0454
0146
FD64
FAD4
FA76
FB28
FB5B
FACF
FA6F
FAC1
FB3B
FB37
FAF0
FB08
FB72
FB7D
FAF3
FA84
FAC6
FB5D
FB96
FB76
FB8F
FBDA
FBA2
FAE1
FB06
FD7B
0193
04D1
058F
04AE
042D
04B7
0552
0533
04D7
04FE
0562
0533
047E
0435
04B8
0541
050D
0483
0478
04D3
04C4
043F
043B
0513
0561
0362
FF62
FBC5
FA7C
FB0B
FB94
FB41
FACB
FAF6
FB68
FB65
FB02
FAE7
FB37
FB64
FB24
FAEE
FB32
FB92
FB71
FAFE
FB02
FB9B
FBDF
FB37
FA9B
FBCA
FF2D
0315
055B
057C
04BB
0467
049D
04C8
04B9
04C5
0504
0513
04BA
045F
047C
04F1
052C
0500
04D5
04EB
04E9
0479
0411
046A
052D
04CA
0228
FE32
FB25
FA51
FAF9
FB87
FB5E
FB15
FB32
FB72
FB63
FB27
FB24
FB55
FB5D
FB39
FB42
FB81
FB79
FAEB
FA6C
FAAC
FB5C
FB76
FAD0
FACD
FCDE
00A2
040C
0582
054E
04D7
04DA
04FA
04C2
046F
0479
04CA
04E2
049D
045C
0471
04B0
04D6
04F5
0534
055A
0510
048B
048F
0557
05CB
045C
00D6
FCF7
FAD6
FADD
FBA1
FBB8
FB1D
FABC
FAF9
FB4C
FB39
FB10
FB57
FBE0
FBF8
FB74
FAEE
FAE9
FB1C
FB06
FACD
FAF3
FB52
FB2D
FA80
FAB5
FD33
015E
04CB
05BC
04DD
0420
0469
04F6
04EF
049A
04AA
0507
0500
0478
0422
046C
04DA
04D7
04A6
04E1
055B
0551
04B3
047E
053C
05BE
0428
0057
FC67
FA84
FAB9
FB5A
FB41
FAD7
FAEC
FB62
FB83
FB36
FB1A
FB7E
FBDE
FBB5
FB44
FB21
FB46
FB2F
FAD2
FAC9
FB4B
FB91
FAEC
FA2A
FB21
FE77
0282
04E7
050F
0478
04A1
0561
059A
04FF
0468
0480
04E3
04DD
0477
044B
048F
04DB
04E6
04E9
0511
050F
04AA
046B
04FB
05D6
054E
0266
FE4F
FB60
FABB
FB5C
FBAA
FB40
FADE
FAFC
FB31
FB10
FAE1
FB21
FBA7
FBD2
FB77
FB13
FB02
FB09
FADD
FAC5
FB23
FB98
FB52
FA60
FA3A
FC50
003B
03DD
057B
054A
04BD
04B7
04F0
04EA
04C6
04E1
0511
04E4
046B
0445
04B4
0525
04FE
048A
0492
0526
056D
04EF
046C
04D0
0587
04B8
017B
FD4B
FAA7
FA73
FB4B
FB7A
FAE4
FA9B
FB17
FBA7
FB95
FB29
FB19
FB6E
FB98
FB5B
FB23
FB3A
FB4A
FB05
FAC3
FB04
FB75
FB3B
FA74
FAAF
FD45
016C
04B4
058F
04D5
0468
04E8
0561
0508
0465
0466
04F8
0532
04BF
044D
0475
04E1
04F0
04BF
04DD
0537
051E
047C
0446
050C
0596
03F3
FFFD
FC02
FA58
FAED
FBC6
FB9C
FB03
FAF9
FB58
FB52
FAEB
FAF3
FB93
FBEA
FB64
FABA
FADB
FB75
FB74
FAC1
FA86
FB54
FC07
FB5B
FA2F
FAF5
FEA6
0330
05A7
056C
0457
0422
04AA
04EC
04BA
04B1
04FB
0509
049C
044C
0499
050F
04F7
0484
048D
052F
057D
04E0
042C
0491
05AB
0576
029C
FE43
FB09
FA50
FB1E
FBAB
FB69
FB16
FB45
FB99
FB81
FB22
FB10
FB5E
FB8D
FB56
FB1C
FB3B
FB6D
FB37
FACD
FAD8
FB58
FB74
FACC
FA89
FC50
001F
03DF
0583
051B
0465
0484
0501
04FF
0496
047A
04BF
04D6
048E
0467
04B5
050A
04E4
0491
04BC
0542
054B
04A8
0459
050F
05C5
049B
0126
FD32
FAE4
FAA4
FB34
FB6F
FB49
FB34
FB3A
FB26
FB18
FB52
FBA8
FBA1
FB32
FAEA
FB21
FB73
FB47
FABC
FA98
FB2A
FBB8
FB66
FA95
FADF
FD5D
0147
0480
0599
0507
0454
046B
04EB
0512
04D0
04AE
04DB
04F4
04B4
046C
047A
04BA
04CD
04C4
04FB
0557
053E
0496
043C
04D4
0557
03DC
000D
FC09
FA3D
FAC1
FBA5
FB89
FAFC
FB18
FBB4
FBC4
FB1B
FAB4
FB23
FBBB
FBA7
FB32
FB25
FB75
FB68
FAE9
FACA
FB58
FBA4
FAE4
FA24
FB71
FF37
0357
0568
053E
0496
04A2
04F7
04D6
047A
0499
0518
052B
0496
0418
0457
04EA
0503
049F
0470
04B9
04EC
04AA
0484
051D
05DA
0518
020B
FDF4
FB0D
FA62
FB08
FB81
FB53
FB0D
FB20
FB51
FB4A
FB35
FB60
FBA3
FB88
FB0C
FAC1
FB04
FB6D
FB67
FB14
FB11
FB66
FB5A
FAB7
FAAD
FCB6
009A
043A
05AC
052B
0473
0492
0502
04EE
0484
047F
04E9
050F
04A8
0452
0497
0512
050B
049E
048E
050A
054E
04D7
0457
04B6
055E
0479
012F
FD0B
FA84
FA60
FB35
FB68
FAF3
FAD0
FB43
FB8E
FB38
FACF
FAFE
FB87
FBA4
FB3F
FB00
FB32
FB4A
FAE3
FA8A
FAF7
FBC0
FBB7
FAD1
FACD
FD4E
019A
0511
05FC
052A
048F
04E1
054F
051F
04AB
049D
04E6
04FC
04C5
04A3
04B8
04BD
04A2
04CD
0555
058F
04EE
0419
0444
0564
05B5
0392
FF79
FBBE
FA2B
FA71
FB0E
FB25
FB00
FB12
FB3B
FB2C
FAFE
FB09
FB4B
FB6A
FB3F
FB0F
FB1A
FB2C
FAF5
FAA9
FAD3
FB72
FBB4
FB0C
FA5E
FB6E
FEE5
0338
05F8
0632
0520
0480
04BA
0506
04ED
04D3
050B
0531
04E2
047C
049D
0522
054F
04F1
04B2
0502
054F
04F8
0483
04F1
05D5
0532
01E4
FD70
FA89
FA27
FAEA
FB2F
FADB
FAC0
FB0F
FB3D
FB15
FB04
FB34
FB32
FAD5
FAAC
FB14
FB7C
FB40
FAC1
FACE
FB3A
FB19
FA83
FB23
FE3E
029F
0593
05E8
0508
04CE
0555
0586
050F
04AC
04C9
04F5
04C5
0486
04A9
0507
052A
0510
050D
0516
04DB
0495
04DC
0558
0479
014D
FD1A
FA4B
F9E6
FACB
FB5D
FB32
FADD
FABF
FAB2
FAA5
FAD0
FB30
FB67
FB52
FB43
FB52
FB24
FAAF
FA95
FB2D
FBAD
FB3E
FAA1
FBC2
FF57
038E
05DF
05C1
04DE
04BB
051D
0522
04CB
04C7
0533
057E
0559
0503
04BE
0487
0474
04B4
0519
050F
0483
0448
04F2
0575
03E7
0001
FBEF
FA11
FA76
FB4E
FB55
FAE0
FAB9
FAE9
FAFE
FAE1
FAD9
FAF6
FAFF
FAF9
FB23
FB65
FB5F
FB1F
FB30
FB96
FB88
FACA
FAAA
FCB8
00A2
0436
05AD
0557
04C3
04C9
050A
0514
0515
053F
0549
0500
04BE
04CF
04EC
04CA
04AF
04EA
0512
049E
0404
0455
056D
056A
02B9
FE5B
FB17
FA67
FB1E
FB64
FAF9
FABF
FAF7
FB05
FAB9
FA9D
FB01
FB6D
FB6A
FB2F
FB26
FB2F
FAFE
FAE6
FB65
FBF3
FB75
FA3F
FA7B
FDA1
023D
0555
05B7
04DF
04A2
0513
0538
04DC
04C4
053A
058D
0538
04AC
047D
0489
0484
04A5
050E
0530
04A0
041D
04BB
05EB
0577
0217
FD64
FA54
FA03
FAE6
FB34
FAE7
FAE8
FB45
FB50
FAF6
FACC
FB04
FB2E
FB14
FB1A
FB71
FBA5
FB55
FAFC
FB35
FB8F
FB17
FA3D
FAF6
FE4E
02AC
0568
05B7
0508
04D7
051B
0516
04BE
04A6
04EF
051B
04E3
04A5
04B1
04D6
04DB
04DF
04E2
0496
0417
0438
054B
0603
0486
00BC
FCC7
FACF
FAD5
FB3D
FB13
FAD3
FB16
FB76
FB57
FAF0
FAE1
FB29
FB4F
FB3F
FB41
FB50
FB22
FAE1
FB1E
FBCB
FBE6
FAE8
FA25
FBAE
FFA8
03B4
0581
0532
0492
04A0
04DD
04B3
0470
0496
04FA
0515
04D8
04A4
049A
048A
0486
04D2
0537
0512
046E
044C
0512
0568
0389
FF9F
FBE8
FA55
FAAD
FB50
FB56
FB2E
FB68
FBC1
FBB5
FB55
FB12
FB18
FB49
FB90
FBC0
FB8B
FAFF
FAC0
FB36
FBBE
FB5B
FA5B
FA86
FD2B
0153
0497
05B4
057A
0536
0516
04B1
043D
044D
04C8
04FF
04BD
0483
049A
049F
044D
041F
0496
0536
051F
048F
04B2
058E
0549
0269
FE0D
FAE6
FA32
FABF
FAF1
FAB5
FAE6
FB93
FBDA
FB5A
FACD
FAE6
FB62
FBA2
FB9E
FB9A
FB83
FB38
FB12
FB5F
FB95
FAF9
FA1A
FACC
FE13
0281
0576
05E2
051B
04CE
051C
0528
04B6
0462
048D
04E8
0511
04FC
04C3
0478
0450
0488
04F1
04F8
0483
045D
0525
05E5
04BA
012D
FD1C
FABD
FA5E
FAB7
FAE2
FB0B
FB69
FB96
FB47
FAF0
FB17
FB75
FB60
FAF4
FAF5
FB79
FBB0
FB47
FB09
FB75
FBB2
FAEB
FA32
FBA4
FF9A
03BE
0596
0538
04A6
04FA
0568
050F
0472
0474
04D9
04D2
046A
045A
04C8
050F
04DC
04A0
04AA
04A1
0450
045C
053D
05C7
0402
FFCE
FBA5
F9F5
FA86
FB4A
FB22
FAB4
FAD2
FB38
FB42
FB0E
FB2C
FBA0
FBD5
FB92
FB3E
FB2D
FB34
FB41
FB91
FBF0
FBA0
FAA3
FA7E
FCC2
00E9
0495
0606
05A4
04FE
04DE
04F7
04FF
0522
055D
053C
04B0
045C
0498
04DB
04AF
0481
04CE
0513
0489
03AF
03E3
0527
0561
02B2
FE20
FAB7
FA0A
FAC9
FB13
FACE
FAE4
FB4B
FB2A
FA81
FA48
FADC
FB68
FB3A
FACE
FAEB
FB4E
FB36
FADF
FB39
FC18
FC18
FB03
FAF3
FDD6
0289
05DF
0646
0530
04B6
0516
053C
04DE
04CE
055F
05BF
0559
04CD
04DE
0544
054E
0510
0509
0515
04C0
045B
04AF
0560
04AC
0174
FD07
FA0B
F9A2
FA87
FB0C
FAF4
FAE0
FAF1
FAD7
FAAE
FAC9
FAFB
FADA
FA92
FAA8
FB0C
FB15
FAAB
FAA4
FB68
FBE9
FB0C
F9DF
FAF3
FF08
03AB
0607
05FA
0572
057D
057F
0500
04B5
0537
05CF
057B
04A6
0496
0567
05D9
0558
04D9
0515
0541
049A
0416
04F7
0634
0513
00C0
FBEA
F9C3
FA60
FB2E
FAAD
F9F7
FA63
FB4E
FB50
FA8C
FA45
FAD0
FB3A
FAF3
FA8B
FA98
FAD5
FADB
FAF4
FB6F
FBAF
FAFB
FA3A
FB90
FF97
040F
0637
05D4
04E1
04DD
0574
05B7
058A
0562
0561
0548
0517
050D
052C
0535
052C
0548
054E
04C6
0415
045F
05B4
0625
03CA
FF4B
FB63
F9F6
FA5D
FADD
FACE
FAB5
FAC9
FA9B
FA25
FA19
FAB6
FB36
FB05
FAAD
FAD4
FB1A
FADD
FA8D
FB14
FC09
FBE1
FA58
F9AB
FC2E
011F
052E
0648
0593
052E
0562
0538
04AC
04C7
05BD
065F
05D6
04D7
0493
050C
055F
0534
04FF
04E5
047A
03FC
0475
05E6
0644
03A0
FED7
FAF2
F9CE
FA75
FAE9
FAA9
FA9A
FB20
FB73
FAF8
FA3C
FA1B
FA94
FB10
FB46
FB43
FB04
FAB6
FAEC
FBCC
FC5E
FB91
FA04
F9F5
FCD1
0148
0496
0581
053C
0548
059C
0569
04C1
047B
04DF
0564
0592
0579
053D
04DD
048E
04B9
053D
053E
045C
03A9
046C
05E9
059A
0246
FDD9
FB46
FB2E
FBB0
FB39
FA4B
FA34
FB0A
FBBF
FBB1
FB3C
FADA
FA8A
FA5E
FAB1
FB68
FBB1
FB2D
FAB1
FB10
FBB4
FB6F
FA9C
FB45
FE95
02F2
0581
0554
0428
03F8
04C4
0541
04E6
0457
043C
0487
04E8
0536
0553
0524
04D1
04BD
04FA
051F
04ED
04D3
0534
054D
03A3
FFFA
FC1B
FA1F
FA50
FB41
FBB2
FB9C
FB8C
FBA9
FBB8
FB9F
FB79
FB48
FB04
FAD8
FAFA
FB39
FB29
FADB
FACE
FB07
FAD9
FA2E
FA57
FCC0
00F2
04A2
0609
0591
04E9
04E4
04F3
0485
0400
040A
048A
04EB
04F4
04D4
04A3
0471
047D
04E8
0549
051C
04B4
0505
0616
063B
03B0
FEFD
FAE4
F98F
FA73
FB72
FB6D
FAFD
FB03
FB76
FBBE
FB9A
FB41
FAF6
FADE
FB0C
FB68
FB8F
FB41
FAE3
FB09
FB6A
FB18
FA18
FA16
FCA9
0126
04F9
0641
057D
0481
0450
048E
04A5
0499
04AC
04C8
04CC
04E1
0525
054B
0517
04D8
04F4
052F
0501
048F
04A2
0548
0524
02C4
FEA2
FB08
F9C7
FA80
FB88
FBE7
FBD2
FBB6
FB8F
FB49
FB1A
FB30
FB4E
FB1D
FAB6
FA88
FABD
FB0B
FB20
FAFB
FAB9
FA7A
FAAA
FC05
FEC9
021F
04A1
059B
0574
0500
04AB
046E
0441
0444
047A
04B5
04C9
04C0
04B7
04BE
04E2
051B
0524
04CC
047A
04EB
060C
0671
0497
00B8
FCD7
FACC
FA8F
FACB
FAB4
FAAB
FB1E
FBA8
FBB2
FB64
FB50
FB8C
FBAE
FB87
FB5B
FB4A
FB1A
FACA
FACF
FB54
FB9B
FAE4
F9F9
FAD7
FE5E
02E0
05C3
0635
0595
0561
0590
054A
047C
03FC
0445
04D6
04F8
04A5
044D
0423
041B
0451
04E4
057C
058D
0529
051B
05C8
063C
04E9
0170
FD52
FA99
F9FC
FA90
FB14
FB26
FB1F
FB41
FB62
FB4D
FB25
FB39
FB94
FBE4
FBDE
FB8D
FB29
FAC2
FA55
FA0B
FA1F
FA76
FAA0
FA95
FB38
FDA7
01AE
0561
06BC
05AD
040E
0399
044C
0504
051E
04EB
04CD
04A2
043F
0403
045B
050A
0569
055E
056D
05BF
05C5
0532
04BB
050E
055B
03CE
FFE0
FB8C
F974
FA1F
FBA4
FC16
FB73
FAF0
FB16
FB5F
FB5F
FB5D
FBA6
FBE3
FBA1
FB14
FACE
FADE
FAC9
FA74
FA73
FB14
FB9E
FB3A
FA80
FB38
FE4B
0267
0537
05C2
051F
04CD
050E
052A
04CA
0464
0460
0478
044E
041C
045D
04EE
0525
04D1
0494
04EF
0566
0529
0465
0430
04E3
051A
0327
FF4B
FBCA
FA87
FB11
FB89
FAFF
FA41
FA5D
FB31
FBCA
FBC7
FB97
FB8C
FB6A
FB0F
FAE8
FB48
FBB1
FB69
FAAD
FA88
FB4C
FBEB
FB6D
FAAE
FBBD
FF43
0356
056C
051B
0440
0488
05A0
061A
0574
048F
0456
04A3
04CE
04A9
048B
049C
04AE
04B5
04E5
0528
0502
0456
03EF
0496
05A0
0524
0213
FDC5
FACB
FA4E
FB20
FB76
FAF5
FA8A
FAC0
FB0C
FADB
FA8A
FAC6
FB6A
FBAA
FB3C
FAC4
FAD2
FB21
FB31
FB34
FBA9
FC39
FBDF
FAA0
FA48
FC9F
0110
04E4
0619
054D
048E
04CD
054B
0537
04E3
04FB
054F
0532
04B2
049D
0532
05A4
053D
0478
0454
04D3
04FC
046D
0418
04C9
057F
0433
0064
FC11
F9C3
F9F4
FAFD
FB43
FAD1
FA99
FAEE
FB42
FB2C
FAED
FAE1
FAF1
FAE5
FAE2
FB26
FB75
FB57
FAE7
FAE0
FB88
FC02
FB65
FA5D
FAEB
FE28
02A2
05AC
061C
0533
04CB
053B
058A
052E
04BD
04E1
0554
0563
04FD
04B2
04C0
04CD
04B1
04C7
0536
0559
04A9
03D4
0424
057B
05CE
0346
FEA9
FAD5
F9BD
FA9C
FB63
FB35
FACF
FADD
FB00
FAAE
FA45
FA82
FB4E
FBC1
FB67
FAD7
FAC2
FB04
FB14
FB09
FB69
FC04
FBE2
FAB8
F9F8
FB95
FFB3
041B
065A
060F
04DA
0456
04AF
052A
0556
0556
0547
050C
04AE
0489
04CD
0523
051A
04D0
04B8
04DC
04BA
0430
03FA
04C1
05B8
04FE
01B2
FD4D
FA5E
F9FD
FAF1
FB6C
FB06
FA9F
FAD1
FB2E
FB26
FAE1
FADA
FB10
FB23
FB0C
FB28
FB79
FB7D
FB0C
FAD0
FB5E
FC1A
FBD7
FAB4
FA9A
FD24
017E
0508
0613
055F
04BE
04E9
053E
0529
04F6
0518
0555
053E
04F4
04F0
0527
050B
0480
042E
0494
0531
051F
0470
042C
04C9
0528
03AE
003B
FC7F
FA49
F9EC
FA6B
FAD6
FB01
FB1B
FB19
FADD
FA93
FA8D
FACA
FAFB
FAFF
FB11
FB50
FB6B
FB16
FAAD
FAE1
FBAE
FC1A
FB69
FA76
FB2A
FE61
02A5
0581
05F5
0530
04E1
055C
05C5
058E
0525
051B
054A
0533
04D9
04B4
04E3
04FD
04CD
04B2
04EE
0513
04A8
042A
048E
05A0
058E
02D5
FE5C
FAD9
F9FD
FAD3
FB45
FAA6
FA06
FA4D
FAFD
FB1A
FAA5
FA75
FAE8
FB65
FB5D
FB15
FB1B
FB5B
FB5C
FB22
FB36
FBA4
FBA8
FADE
FA5C
FBD9
FF9D
03C9
061D
0624
054C
04FE
0547
056F
053F
0525
0555
056D
051B
04B0
04A4
04DF
04E4
049D
0480
04C7
04FB
04B2
045C
04B2
0554
04AA
01AB
FD71
FA63
F9C9
FAA7
FB2F
FAD5
FA73
FAB4
FB2D
FB27
FAB7
FA86
FAD0
FB2E
FB52
FB66
FB8A
FB6E
FAE9
FA89
FAF1
FBBD
FBCF
FAFE
FAE7
FD3F
0182
0523
0630
0549
0487
04E5
0584
0557
04A9
0480
0508
0573
0535
04BD
04AC
04EA
04F9
04D8
04ED
0532
0519
048B
044C
04DC
053A
03A5
FFDB
FBD8
F9EF
FA5A
FB4F
FB52
FABA
FAA6
FB39
FB8A
FB20
FAA1
FACE
FB67
FB97
FB2D
FAC7
FACA
FAE8
FACF
FAD0
FB44
FBB6
FB6C
FACF
FB88
FE96
02C2
0593
05EA
04F9
048E
0500
0550
04EC
046F
0493
051E
0553
0511
04E1
0500
050F
04D6
04BE
0522
0589
053F
0484
0460
0503
04F5
02A1
FE80
FAFA
F9DE
FA9B
FB49
FB0A
FAA3
FAED
FB8C
FB9B
FB10
FAB7
FAF6
FB4A
FB27
FAD5
FAE2
FB32
FB2B
FAC8
FAB3
FB2E
FB76
FAF9
FAAB
FC56
0044
045C
0632
059C
0495
04B7
058D
05BA
0504
0474
04B7
0539
0529
04AA
0474
04AB
04CD
04A9
04B7
0535
058E
0532
049D
04C1
0556
04A2
017F
FD1D
FA0E
F998
FA9C
FB3E
FAFD
FAAA
FAD9
FB1C
FAEE
FA94
FAAB
FB30
FB94
FB90
FB69
FB54
FB1C
FAB0
FA8D
FB12
FBB4
FB80
FA9E
FAB4
FD29
014E
04D0
0619
05B1
052E
053E
0557
0502
04A9
04DA
0557
0567
04EC
0486
04A1
04E9
04E9
04D2
0514
057E
0568
04CD
0489
050B
053B
037C
FFCE
FC2B
FA79
FA8E
FAD8
FA84
FA4A
FAE5
FBBB
FBAB
FABF
FA2F
FAB2
FB96
FBCB
FB53
FAFB
FB06
FAF3
FA91
FA7E
FB13
FB83
FAF3
FA27
FB29
FED1
0357
0604
0606
04FB
04AF
052C
055E
04E3
0470
0495
04FD
051B
0501
0509
0515
04C6
044C
0460
052D
05D0
0580
04C4
04CE
0592
0556
02AA
FE67
FB09
FA13
FAA9
FB01
FA92
FA4E
FAE7
FBBB
FBC7
FB14
FA90
FAC7
FB48
FB79
FB67
FB6D
FB70
FB18
FA97
FA99
FB2B
FB64
FAB4
FA41
FBF6
0012
0455
0639
0598
0481
048C
053F
0553
04B8
047E
050D
0580
050D
0442
042C
04C4
0511
04AC
0455
04AD
0534
0522
04CB
0521
05D7
0518
01B7
FD1A
FA05
F9AF
FAC3
FB5A
FB20
FAFA
FB4D
FB7B
FB17
FAAB
FADF
FB70
FBA6
FB6A
FB42
FB53
FB2D
FAB5
FA9A
FB4C
FBF6
FB60
F9F1
F9D8
FCB4
0170
052A
0634
0575
04D6
0505
0547
0509
04B7
04DB
0530
050D
0478
0424
046A
04CE
04D2
04AD
04E1
0549
0546
04CD
04AF
0557
05B3
0410
003D
FC2F
FA23
FA5A
FB31
FB3F
FABE
FAB0
FB39
FB86
FB20
FAA3
FACF
FB71
FBB7
FB68
FB21
FB4A
FB71
FB0B
FA6B
FA5A
FAE8
FB4B
FB3A
FBBF
FE17
01DC
050F
0624
058B
04DA
04E6
0531
0510
04AA
0489
04BB
04D8
04BE
04B6
04E2
04FC
04DD
04D6
0528
057A
0554
04FD
052B
05B3
0529
0270
FE6B
FB65
FAA5
FB36
FB59
FAAA
FA29
FA83
FB22
FB34
FAE9
FB05
FB99
FBE4
FB7F
FAFC
FAFD
FB3F
FB1D
FAB8
FAD2
FB7A
FBA6
FAB3
F9CB
FAFB
FEBE
031D
05A2
05CF
0528
051E
059D
05BF
0549
04DB
04E8
051A
04F1
048D
046D
04AC
04D6
04A2
0464
0494
0515
054F
0506
04C8
053E
0616
05F9
03D1
0012
FC7D
FA98
FA69
FACA
FAD0
FA96
FAB6
FB40
FB9F
FB68
FAEF
FAD1
FB23
FB68
FB4A
FB09
FB0E
FB53
FB6A
FB2A
FAEC
FB03
FB31
FAF9
FA72
FA8D
FC45
FF8F
032B
0599
063F
05AF
04ED
0492
0499
04BE
04E6
050C
0513
04D9
047C
045B
04A4
0509
0519
04D6
04B3
04E9
0510
04B9
0439
0469
055C
05BE
03F9
0012
FBFB
F9D3
F9FD
FB1A
FBB2
FB85
FB32
FB1B
FB0E
FAD9
FABB
FAFF
FB72
FB98
FB4F
FB02
FB0E
FB45
FB3D
FAF8
FAF3
FB66
FBC9
FB6F
FAA3
FAC4
FCFE
00D6
045A
05D8
055A
0455
040C
047D
04E1
04DC
04C9
0503
054B
0535
04D4
04AE
04F1
0528
04DA
044F
043F
04D3
0558
0527
048B
0460
04BF
0485
0280
FEF5
FBA7
FA32
FA94
FB79
FBC0
FB69
FB17
FB16
FB21
FAFF
FAE3
FB0C
FB4E
FB40
FAE1
FAB1
FB0A
FB91
FBA1
FB27
FAD1
FB25
FBBB
FBBA
FB1F
FB2D
FD31
00E4
0465
05F3
0588
0497
045E
04D3
0529
0504
04C8
04D3
04F1
04CB
0482
048D
0503
055F
0538
04D2
04BA
04EF
04DC
0448
03E4
0474
057B
0551
02D1
FECA
FB6D
FA34
FAA5
FB32
FB03
FA92
FAA4
FB28
FB69
FB19
FAB9
FAE0
FB66
FB9B
FB36
FAB9
FABD
FB2B
FB66
FB31
FB02
FB44
FB9B
FB56
FAA0
FAD1
FD1B
0101
0480
05F4
0599
04F3
04FF
0559
0538
04AF
0486
0507
0585
0550
04AD
0473
04D6
0528
04DA
0458
046E
0514
056C
04FF
0484
04E0
05B0
0550
02B2
FEB7
FB76
FA33
FA71
FAEB
FB08
FB0D
FB3A
FB4D
FB05
FAA8
FAB4
FB23
FB66
FB27
FAC6
FAD4
FB45
FB7A
FB1E
FAAF
FADA
FB81
FBB8
FAF4
FA04
FA86
FD4D
0160
04BB
0609
059E
04D1
049A
04E7
0520
050C
04EE
04FD
050C
04D9
048A
0490
050C
0588
0583
0511
04BC
04C5
04D6
049E
046B
04C8
0570
051B
02B7
FED1
FB59
F9E2
FA3E
FB00
FB23
FAD7
FACB
FB20
FB60
FB49
FB2A
FB57
FB98
FB75
FAEC
FA89
FAAE
FB14
FB2E
FAF6
FAEA
FB46
FB8A
FB28
FA84
FAF5
FD6E
0147
04A1
0613
05D1
0527
0505
0541
0543
04F1
04B1
04BC
04CA
049A
0463
0488
04EC
050A
04B5
0478
04DB
0586
0591
04C8
0422
0492
058C
053A
0273
FE2D
FABF
F9A6
FA5C
FB40
FB59
FAF1
FABD
FAE5
FB12
FB0E
FB0F
FB4A
FB9A
FBAA
FB6E
FB33
FB32
FB3B
FB06
FAAB
FA9A
FAFD
FB5B
FB2C
FAC8
FB70
FE0C
01EF
0527
0646
05A2
04BF
049F
04FD
051A
04DF
04CD
0513
0536
04CD
0432
0418
049D
0523
0528
04E6
04E5
052D
0540
04EB
04AA
04EE
0535
0448
018D
FDE9
FB13
FA0F
FA6D
FB02
FB20
FAFE
FB09
FB3B
FB3F
FB0C
FB03
FB5F
FBCB
FBBE
FB32
FAB6
FABC
FB06
FB0B
FAC5
FABA
FB26
FB7B
FB26
FAA2
FB59
FE26
0222
0549
064B
0599
04A6
0464
04B2
04FB
04FF
04E6
04D7
04C4
049D
0482
04A2
04F7
053E
0542
0512
04E4
04D1
04C3
04B1
04D0
0545
0591
049A
01B1
FDA8
FA7F
F9A7
FA9F
FB9B
FB7A
FACD
FABF
FB71
FBE7
FB7E
FACA
FAB3
FB33
FB7B
FB2C
FAD1
FAF7
FB57
FB52
FAFB
FB02
FB8A
FBC1
FB10
FA56
FB46
FE74
026D
0511
0599
0508
04C3
0528
0590
0568
04D9
047A
0498
04F5
0523
04F8
04AC
048B
04A4
04C6
04CC
04C3
04BE
04AA
047C
046F
04C8
0529
046F
01C7
FDE7
FAD3
F9FF
FADE
FBA4
FB4E
FA83
FA5F
FAE7
FB32
FAD7
FA87
FB03
FBF0
FC49
FBBA
FB04
FAEF
FB54
FB8B
FB6F
FB74
FBBE
FBB5
FAF6
FA5A
FB70
FEB8
02C1
0562
05C1
04EC
047A
04E0
055F
0540
04BC
0484
04C7
0504
04D5
0479
046F
04B6
04D2
0484
0428
042F
0475
047C
0443
0469
052F
05A6
0459
00FC
FD10
FA9F
FA51
FB0E
FB67
FB09
FAA5
FAC5
FB26
FB47
FB29
FB39
FB9D
FBF3
FBD5
FB6A
FB37
FB76
FBD0
FBDF
FBB2
FBA4
FBB7
FB76
FAAE
FA30
FB5F
FEB6
02E5
05BB
0623
0515
045E
04B9
0558
0541
049E
045F
04E3
0570
053E
047B
03F9
0415
045A
0452
042B
044E
049A
048F
0430
0432
04EC
0573
0442
00FC
FD14
FA8B
FA16
FAC0
FB37
FB1F
FAFF
FB3B
FB8D
FB7E
FB16
FACA
FAE3
FB2E
FB55
FB50
FB60
FB9C
FBC9
FBB8
FB97
FBB3
FBE9
FBA8
FACF
FA50
FB96
FEFD
0313
05BA
0617
0536
04AA
04E9
0538
04FA
048B
0496
0509
052C
04BA
044F
048F
052C
0548
04AE
041D
0442
04C2
04C4
0442
042F
050A
05BE
0487
0100
FCE1
FA6F
FA50
FB36
FB8C
FB0C
FA8C
FAAC
FB1D
FB45
FB15
FAF5
FB10
FB18
FAD9
FAA8
FAF9
FBA7
FC00
FBA5
FB17
FB13
FB8A
FBA4
FAFE
FA8D
FBDD
FF42
032E
0586
059C
049B
0414
0478
0510
0534
0502
04F4
051A
0521
04F4
04E6
0531
0580
055A
04D2
047D
04A7
04E5
04B4
044F
047C
0553
05A2
03F8
004D
FC62
FA34
FA35
FB30
FBC0
FB97
FB48
FB3F
FB4F
FB35
FB0F
FB20
FB4C
FB34
FACB
FA85
FABC
FB29
FB3C
FAE9
FACA
FB47
FBDB
FB9E
FA93
FA19
FBBA
FF77
0385
05D9
05F1
0502
0484
04CF
052F
050A
0494
045F
048A
04B3
049F
0495
04E5
055D
0578
0516
04AD
04A7
04CF
04B9
0488
04D7
05A9
05D5
0401
0045
FC69
FA58
FA5E
FB2B
FB6A
FAFC
FAA2
FAD3
FB47
FB80
FB65
FB3A
FB2F
FB31
FB21
FB03
FAEE
FAE7
FAEF
FB17
FB6C
FBBE
FBA7
FAF4
FA21
FA46
FC4C
FFF7
03C1
05EF
0600
0502
046C
04B2
0524
050D
049C
047C
04D8
052E
051E
04EF
050F
054F
052A
049C
0446
048D
0501
04FE
04B0
04E0
05A4
05B8
03B2
FFC2
FBCD
F9B8
F9C7
FABF
FB55
FB3F
FAFB
FAFD
FB40
FB7F
FB8B
FB63
FB1D
FAD5
FA9F
FA91
FAB8
FB0C
FB59
FB6B
FB4A
FB31
FB39
FB26
FADA
FAE8
FC59
FF8B
035D
05F7
067B
05BB
0520
0523
053A
04EF
048C
0495
04FE
0544
0529
04EB
04C8
04B2
049F
04C7
053B
0585
0521
0455
0413
04D1
05B7
0547
02DF
FF67
FC6B
FAD8
FA8A
FAC8
FAF3
FAD3
FA9A
FA9F
FAF5
FB4F
FB55
FB0F
FAD4
FAD5
FAE4
FACD
FAAC
FAC2
FB09
FB45
FB6C
FBA4
FBC6
FB61
FA92
FA83
FC76
0035
03E7
05C3
05B8
051F
0507
0543
0534
04D3
049E
04CA
0510
0527
0518
0503
04ED
04E0
04FD
0542
055C
0511
04A3
0480
049C
048E
045E
049F
0555
0547
0320
FF34
FB9A
FA22
FA98
FB64
FB7D
FB31
FB1A
FB22
FAF4
FAB9
FAD9
FB33
FB3E
FADF
FAA1
FAE0
FB38
FB1B
FAAD
FA90
FAF6
FB6A
FB91
FB98
FBA2
FB62
FADB
FB0F
FD26
00D1
0429
0588
052A
0495
04B2
050D
04F2
0484
045C
0498
04D4
04DF
04E7
0504
050E
04FC
0504
0539
0551
0515
04D4
04EB
0513
04BD
0422
0432
0509
051D
02CF
FEA3
FB17
FA0F
FAF5
FBC7
FB88
FAF2
FAEF
FB58
FB7B
FB40
FB19
FB30
FB45
FB38
FB3A
FB54
FB40
FAE3
FA9B
FAB6
FAF3
FAEF
FADB
FB36
FBCB
FBC2
FB17
FB46
FDBD
01D3
0523
0603
051F
0450
046E
04DB
04E6
04C0
04DD
051B
050E
04BE
0490
049F
04AF
04AB
04C8
0507
051D
04F1
04DA
0509
0513
0492
040A
0462
0541
04DA
01F0
FDAD
FA9E
FA02
FAC9
FB43
FB12
FAF3
FB35
FB54
FB02
FAB4
FAD8
FB1C
FB0A
FAE0
FB1F
FB9C
FBA5
FB1A
FAB9
FB08
FB92
FBA5
FB62
FB64
FB89
FB16
FA4E
FAEB
FE22
02B6
05E5
064C
0521
046D
04CB
0554
054D
04F9
04DC
04EC
04ED
04F7
0528
053D
04F3
0493
049C
04EF
04F5
048F
044E
048B
04C5
0479
0428
04AD
057C
04A9
013D
FCD5
FA21
FA04
FAFD
FB59
FB01
FADD
FB23
FB35
FAD4
FA93
FAD5
FB27
FB06
FAC0
FAE6
FB53
FB62
FB00
FACA
FB0A
FB4D
FB37
FB31
FBB1
FC30
FBCE
FB01
FBA8
FECB
02F4
0596
05CA
04E8
048D
04E6
052D
051D
0521
055D
0565
050B
04BF
04D2
04F0
04BC
048C
04E1
057A
059C
052B
04CD
04CE
04A0
03E4
0361
040B
0523
047A
0113
FCBA
FA36
FA4A
FB50
FB8D
FAFF
FA9C
FAB6
FAD1
FAB2
FABA
FB17
FB5C
FB37
FAF9
FB05
FB24
FAF7
FAB7
FAE3
FB57
FB73
FB2B
FB41
FBFF
FC69
FB92
FA76
FB62
FF21
0397
05F1
05AB
04A4
0482
0511
0546
04F1
04BC
04F2
0520
0500
04E6
050E
0522
04D8
0492
04BF
0511
04EB
046C
044C
04AB
04C4
0433
03D5
048F
0579
0469
00AC
FC4F
FA06
FA42
FB36
FB52
FADA
FAD6
FB5F
FBB0
FB66
FAF0
FAC1
FAC7
FAD5
FB0B
FB69
FB88
FB30
FAD8
FB04
FB6B
FB64
FB04
FB1B
FBD0
FC13
FB26
FA45
FBAA
FFB6
040D
060E
059E
04BA
04C3
053C
0524
0490
0453
04A4
04F6
04EF
04D7
04EA
04E3
049A
0470
04B6
0508
04E2
0482
0492
0500
0500
0468
0436
0511
05B6
040C
FFE8
FBC3
FA20
FAD7
FBBF
FB80
FAC1
FAA6
FB28
FB73
FB44
FB17
FB34
FB46
FB1B
FB03
FB34
FB54
FB1A
FAE7
FB2F
FB9A
FB78
FAE9
FAD0
FB69
FBBD
FB1A
FAA4
FC52
004A
043A
05D6
054A
0481
049D
050B
04FC
04A9
04BA
0516
0515
049F
0456
0493
04E2
04D8
04B5
04D9
0509
04E4
04A4
04CB
0526
04FD
0453
042D
0500
056C
0386
FF6F
FB9A
FA27
FAAB
FB3F
FB08
FAC7
FB26
FBA0
FB75
FAE3
FAC0
FB2F
FB7D
FB51
FB1A
FB37
FB4C
FAFA
FA9E
FAC3
FB33
FB50
FB24
FB4E
FBCA
FBB2
FACA
FA92
FCD4
0125
04DD
05F7
052F
049F
050D
0577
0506
044D
043D
04C0
050E
04ED
04DC
0512
0524
04DE
04B8
0509
0556
0510
0489
0478
04C9
04BD
0442
0443
0512
053F
0305
FEC5
FB15
F9EC
FAA3
FB3E
FAFD
FAB9
FB14
FB88
FB69
FB01
FAFE
FB47
FB2F
FAA3
FA5D
FAC2
FB3D
FB37
FAF6
FB09
FB55
FB63
FB52
FB9F
FC0D
FBB6
FAA9
FAA8
FD54
01CD
053B
05E8
04F6
0484
0504
054F
04CE
0452
04A6
0551
0566
04EC
04B9
0513
055E
0532
04F6
050B
051B
04C9
0478
04A6
04EB
0483
03C0
03E9
0529
0588
02FC
FE3C
FA6A
F9A3
FADA
FBA0
FB23
FA81
FAAC
FB31
FB49
FB07
FAFB
FB2E
FB32
FB05
FB12
FB58
FB47
FAC1
FA74
FAD1
FB46
FB29
FAE1
FB3C
FBEE
FBCA
FACC
FAE3
FDC6
0268
05C0
062D
0514
04AC
0543
058F
04FB
0467
049C
0529
0535
04D1
04AA
04E3
0501
04E8
050C
0580
0599
0504
0478
04A8
0516
04DC
0444
0479
0568
050F
01D8
FD12
F9F0
F9ED
FB56
FBC0
FAE6
FA43
FA9B
FB24
FB0E
FAAD
FAB2
FB06
FB13
FAD2
FAC0
FAF7
FB02
FACF
FAEA
FB75
FBBB
FB48
FAD9
FB43
FBEE
FB85
FA4D
FA91
FDF5
02F2
062E
0630
04BF
044D
051B
05BE
0581
0517
052B
056A
054C
0505
0511
054F
0540
04F2
04E9
0526
050D
047B
042F
049A
0505
04B3
043F
04C8
05CC
0522
019F
FD04
FA4A
FA48
FB24
FB0E
FA5E
FA59
FAFC
FB28
FA84
FA00
FA53
FAF8
FB25
FB03
FB38
FBA4
FB86
FAD0
FA6C
FAD7
FB62
FB52
FB12
FB54
FBAE
FB2A
FA46
FB10
FEA7
0351
060F
05EA
04BA
048D
0553
05BA
055C
0509
054A
05AA
0598
0539
04F5
04C7
047C
044A
0488
04FB
050B
04C4
04D1
0549
0558
049C
041E
04E7
05FA
04ED
00E8
FC20
F99A
F9EB
FB11
FB45
FAD0
FAC7
FB29
FB27
FAAF
FA83
FAEC
FB49
FB20
FAE2
FB23
FB93
FB79
FAF0
FAC7
FB3A
FB8D
FB4F
FB12
FB5C
FB8A
FAE3
FA4A
FBBF
FFBD
0411
0614
0591
049F
04C8
0576
056A
04BD
0479
04E3
0530
04E3
047D
0493
04EF
0504
04D8
04DA
0508
04F0
048E
046B
04B0
04CA
0471
045F
0522
05A4
03F9
FFE1
FBA0
F9C0
FA64
FB82
FB86
FADC
FAB5
FB3A
FBA0
FB7F
FB32
FB12
FB0C
FB09
FB2D
FB75
FB86
FB2F
FAD7
FAF0
FB3D
FB2F
FAF1
FB3F
FC0D
FC32
FB2B
FA78
FC3A
006E
0486
0621
057D
04A5
04B5
04FA
04A5
0430
047B
053F
0573
04D7
0442
045F
04D4
04FA
04D8
04DF
050A
04EC
048B
0467
049F
04A3
043E
0423
04CC
052D
0385
FFA8
FBAF
F9E9
FA7A
FB8E
FBAB
FB14
FAD1
FB2E
FB9B
FBA9
FB70
FB28
FAE8
FACE
FAFD
FB54
FB7E
FB66
FB59
FB87
FB9D
FB4E
FAFD
FB46
FBE1
FBC7
FAD1
FA92
FCB9
00D3
0473
05C0
053C
04B2
04EB
0530
04DB
0463
0486
0513
0540
04DB
047B
048B
04BE
04AD
0476
0477
04AD
04BB
0483
0447
043A
044B
0488
0522
05BC
0529
028F
FEB1
FB88
FA66
FAC7
FB36
FB03
FAA5
FAA7
FAE7
FAFF
FB02
FB3D
FBA1
FBC7
FB92
FB59
FB6D
FBB0
FBD1
FBA8
FB49
FADF
FAB5
FB1A
FBEF
FC62
FBBA
FA8C
FAA3
FD29
0129
0463
059A
0588
0587
05D4
05AF
04D8
041F
0447
04F7
053F
04D8
0456
0437
044D
0440
0425
044E
04AC
04DE
04C3
04AE
04D3
04E7
0496
042F
0459
0522
059C
04A4
0201
FE9C
FBCC
FA5D
FA40
FACC
FB4B
FB61
FB29
FAFB
FB07
FB35
FB59
FB6C
FB80
FB97
FBA0
FB9A
FB93
FB8F
FB85
FB77
FB70
FB5D
FB14
FAAF
FA9C
FB20
FBC0
FBA8
FAE7
FAE0
FCFD
00E6
0478
05D7
0536
0457
0470
0515
0544
04D6
047E
04A0
04D1
049C
043A
0435
0492
04D2
04B5
0485
0486
0489
044E
0424
0489
054F
059C
050B
0462
04A5
0589
0568
0309
FF27
FBD5
FA73
FA99
FB06
FB16
FB13
FB55
FBA4
FB9E
FB4F
FB1E
FB33
FB4E
FB3B
FB2A
FB62
FBC4
FBE1
FB88
FB11
FAF3
FB2D
FB53
FB29
FAF8
FB14
FB4A
FB19
FA97
FAD1
FCDB
0074
03DF
056E
0516
0447
0445
04EF
0555
050D
0495
047D
04AB
04B5
0494
049D
04D4
04D3
0474
0431
047D
050A
0528
04C6
0490
04E6
0534
04CA
0419
0449
0571
05E4
03E3
FFCF
FC0B
FA8B
FB03
FBB5
FB90
FAFA
FAB8
FAD5
FAE9
FAEE
FB38
FBB9
FBE3
FB70
FADE
FAD4
FB40
FB78
FB2D
FAD9
FB07
FB82
FBA0
FB3D
FAF8
FB46
FBAC
FB4E
FA4C
FA1B
FC25
001A
03EA
05AB
0551
046A
044A
04D6
0522
04D4
047F
04AF
051C
051C
04A3
044B
0471
04B7
04AC
0484
04BF
0549
0571
04EE
0469
049E
0549
0575
04E6
047F
04E1
0521
0395
FFFA
FC28
FA4E
FABD
FBDA
FC1A
FB77
FAE6
FAEE
FB3F
FB6C
FB70
FB6D
FB50
FB07
FAD6
FB14
FB96
FBC3
FB54
FAC3
FAB4
FB19
FB48
FAF2
FA9C
FAE5
FB8B
FBA7
FAFC
FAAF
FC41
FFCA
038A
0579
052C
0406
039E
043E
050F
0554
052A
050C
0513
04FE
04C5
04B1
04E1
0506
04D4
0485
048B
04E8
0519
04D2
0476
0489
04EA
04F8
0498
0477
0506
056D
0425
00C7
FCDD
FA88
FA77
FB74
FBEB
FB79
FADE
FABD
FAEB
FAEF
FAB5
FA90
FAAC
FAE2
FB0B
FB35
FB6A
FB83
FB59
FB1F
FB2D
FB7B
FB99
FB49
FAF0
FB12
FB7D
FB61
FA82
FA06
FB89
FF42
0366
05BC
05B5
04AF
044B
04CB
0556
0550
0506
0501
0537
053E
0504
04E7
051B
054B
0519
04AB
046D
0475
0474
044A
0450
04C3
053C
0525
04A0
048C
0548
05C9
046F
00E8
FCD9
FA65
FA2B
FAF6
FB46
FAD5
FA66
FA86
FAEA
FB0E
FAF1
FAF6
FB31
FB48
FB07
FABE
FAD7
FB39
FB6A
FB45
FB2C
FB6C
FBB1
FB79
FAEE
FACB
FB51
FBBD
FB4C
FA9E
FB6F
FE9D
02D4
05AA
060B
0520
04B0
052C
05A4
0562
04D2
04BA
051B
0550
0511
04CB
04E1
0515
04F9
04A8
049C
04E5
0503
04AA
0443
0457
04BE
04D8
0490
0499
0551
05C2
0466
00F6
FD12
FABD
FA77
FB0D
FB30
FAC5
FA83
FABC
FB00
FAE7
FAB1
FAD8
FB52
FB8F
FB4A
FAEB
FAF1
FB43
FB5B
FB15
FAEC
FB44
FBC0
FBB6
FB2A
FAD9
FB31
FB97
FB41
FAA5
FB65
FE76
02A0
057A
05D6
04D7
0460
04F2
058C
0556
04BD
04A3
0508
0526
04B2
0450
0498
052B
0540
04CA
0487
04D9
0530
04E9
044F
0432
04B6
0510
04C2
0465
04C2
0560
04AE
01DC
FE0B
FB3E
FA5A
FA91
FAB1
FA7B
FA79
FAE3
FB53
FB65
FB45
FB48
FB65
FB52
FB14
FB0B
FB5F
FBA6
FB6E
FAE7
FABD
FB33
FBBE
FBB6
FB3A
FB07
FB68
FBAE
FB1C
FA38
FAB5
FDA0
01EA
052A
05F9
0531
04B1
0536
05D8
0596
04B7
0447
0497
04F1
04BF
0467
048F
0511
052C
04B4
045D
04B2
0530
04FD
0433
03CC
0442
04E5
04ED
04AE
0505
05B6
0533
0267
FE49
FB19
FA22
FAA9
FB28
FAFF
FAA8
FAAA
FAF4
FB36
FB62
FB8C
FB99
FB65
FB19
FB0E
FB50
FB7F
FB53
FB13
FB3D
FBCB
FC1E
FBC6
FB17
FAD3
FB35
FB97
FB3D
FA80
FACC
FD41
0144
04C6
061B
057E
0496
0495
0526
0542
04B2
0440
047D
04FA
04FF
0499
0478
04D8
0525
04D4
042E
03E7
0423
0468
0477
04A0
0506
052C
04AF
0428
048F
05A7
05B2
0334
FEE5
FB32
F9D8
FA67
FB36
FB58
FB28
FB37
FB6F
FB6B
FB2B
FB08
FB24
FB3E
FB2A
FB1B
FB4E
FBA6
FBD1
FBC0
FBAE
FBBD
FBBC
FB73
FB07
FAE2
FB28
FB73
FB3C
FAB1
FAE4
FCE5
0087
0426
05FB
05B6
04A9
0450
04D4
053F
04F6
0476
0481
04FE
052B
04BB
043E
0451
04C5
04F7
04B6
0465
0454
0459
044E
0466
04C8
0515
04E2
047E
04AC
055A
0531
02F1
FF23
FBE1
FAB7
FB25
FB8A
FB1A
FA79
FA82
FB13
FB67
FB36
FAFF
FB35
FBA2
FBC0
FB7A
FB3E
FB59
FB9F
FBB8
FB96
FB6D
FB5B
FB49
FB2E
FB33
FB74
FBAB
FB68
FACA
FAD3
FC9C
0017
03BA
05BA
05A8
04B9
0462
04DF
054C
0507
0475
045C
04C9
0517
04E6
0498
04A5
04E5
04D1
045F
041D
0463
04D2
04EB
04BC
04AA
04B3
047D
041F
0447
0523
0584
03D1
0001
FC16
FA2E
FA71
FB45
FB58
FAE6
FADC
FB62
FBC5
FB99
FB3F
FB39
FB68
FB5A
FB0C
FAEC
FB26
FB63
FB4E
FB17
FB22
FB69
FB86
FB55
FB38
FB7C
FBC5
FB75
FAB3
FAAF
FC8F
001F
03B9
05A8
05A1
04CF
047C
04DA
0534
050F
04B6
04A1
04BA
048A
040D
03E2
0474
054C
0595
052D
04C1
04CB
04EF
04AB
0437
0435
04AA
04E4
0492
0460
04EC
0563
040D
0068
FC38
F9DF
F9FA
FB17
FB99
FB54
FB0C
FB1C
FB2B
FB05
FB04
FB72
FBEB
FBDF
FB62
FB08
FB0D
FB11
FACD
FA99
FAED
FB93
FBD0
FB65
FAF4
FB25
FBA6
FB8A
FAB8
FA7E
FC51
000E
03D5
05BF
0591
04A9
045B
04BD
050F
04EA
04A7
04B7
04FA
0504
04C2
0492
04A8
04C1
0490
0443
044F
04BE
0515
04FC
04BC
04D3
052B
053C
04E5
04BD
0528
0557
03DB
005C
FC65
FA12
FA08
FB0D
FB99
FB68
FB37
FB6D
FB95
FB42
FAC5
FABE
FB2C
FB75
FB50
FB29
FB67
FBC2
FBAA
FB36
FB0E
FB67
FBA0
FB32
FA93
FAA8
FB5D
FB9C
FAD9
FA40
FB9E
FF38
0338
057F
05A8
04F9
04AC
04D4
04E7
04BD
04AD
04E6
051F
0501
049D
0454
045D
049D
04D9
04F2
04E5
04BD
0493
0485
049D
04BD
04BD
049B
0494
04EE
057C
0575
03F5
00E5
FD67
FB12
FA9B
FB42
FBB0
FB55
FAB4
FA7C
FAB0
FAE5
FAFE
FB3B
FBA6
FBD7
FB85
FB09
FAF9
FB57
FB98
FB6B
FB2C
FB41
FB79
FB5D
FB08
FB17
FBA5
FBE4
FB2E
FA4D
FB01
FE09
020A
04D2
0582
0515
04E6
0539
056E
0531
04E3
04E2
04FB
04C7
0458
0422
045C
04BF
04EE
04DF
04BF
04AA
0494
0473
045C
0464
0495
04E7
0532
0532
04D5
0485
04C4
0551
0500
02D7
FF4D
FC11
FA7E
FA73
FAD7
FAED
FAD5
FAE1
FB0C
FB2F
FB5D
FB9F
FBB6
FB68
FAFB
FAF0
FB52
FB9D
FB79
FB2C
FB25
FB49
FB32
FAED
FAF4
FB58
FB8C
FB49
FB15
FB6A
FBC6
FB5B
FA99
FB39
FE3F
0267
0545
05CB
051C
04CC
0518
053B
04E8
049E
04C0
0509
0514
04E6
04BD
04A1
047B
0461
047B
04AB
04B1
04A5
04DD
053F
0535
0499
0419
0447
04AC
047D
03FC
044D
0594
060B
03C3
FF33
FB1F
F9B7
FA86
FB80
FB80
FAFB
FAB8
FAC1
FACE
FAE5
FB2F
FB74
FB5C
FB0A
FAFE
FB58
FBA3
FB89
FB4F
FB4C
FB57
FB26
FAF0
FB21
FB98
FBBC
FB69
FB3D
FB98
FBD5
FB33
FA5F
FB3C
FEA8
0313
05EE
063B
0534
0485
049D
04E3
04EF
04EF
050A
050B
04D2
049F
04AC
04C5
04A9
047F
048F
04C0
04BA
0482
0481
04D2
04FC
04AB
044B
0477
04F5
04F8
046A
043C
04DF
0510
0315
FF0D
FB3F
F9C0
FA50
FB14
FAF0
FA7C
FAA0
FB38
FB85
FB5E
FB3E
FB61
FB7A
FB55
FB2B
FB3B
FB65
FB6F
FB6A
FB7B
FB7A
FB2D
FAD4
FAEE
FB60
FB7B
FB11
FAE3
FB78
FC0C
FB90
FA91
FB21
FE66
02DC
05C6
061F
0555
0518
056E
0569
04DD
0486
04C3
0518
0512
04E2
04D4
04B6
0444
03D5
0406
04C0
0535
04FF
04A3
04AA
04D1
049B
0442
045E
04D2
04E3
0472
0450
04E5
050C
0327
FF56
FBB8
FA2D
FA70
FAE6
FABC
FA78
FAB1
FB24
FB3D
FAFE
FAE3
FB1E
FB67
FB7D
FB6E
FB52
FB23
FAFA
FB19
FB72
FB8E
FB32
FAD6
FB0A
FB94
FBB7
FB55
FB2A
FBAB
FC24
FBB4
FAF0
FBAA
FEC5
02CC
055B
05A2
04E8
04B8
053A
059A
0568
0504
04DC
04E1
04DE
04E3
050C
0523
04E5
047E
0459
048A
04B9
04B3
04B2
04F2
053B
052A
04C7
0472
0449
040C
03CD
040D
04D2
04EF
02F9
FF1D
FB68
F9D6
FA58
FB39
FB3C
FAC2
FAB9
FB31
FB72
FB2E
FAD9
FAE6
FB26
FB2C
FAF9
FAE8
FB1B
FB57
FB6C
FB67
FB58
FB31
FB0A
FB21
FB72
FB9F
FB78
FB59
FB9A
FBD9
FB81
FAFC
FBC3
FEB6
02AA
055B
05C8
050E
04BF
0517
0544
04ED
0497
04AF
04EE
04EE
04D5
0500
054B
053B
04C0
045A
045A
047D
047C
0487
04D1
0511
04EB
049A
049B
04D2
04A7
041D
0417
04FB
057A
03AD
FF84
FB5D
F9A2
FA4D
FB61
FB68
FAC2
FA86
FAF4
FB6C
FB75
FB3B
FB11
FB04
FB04
FB2A
FB7A
FBB0
FB8D
FB31
FAEA
FAD0
FAD1
FAF7
FB4C
FB92
FB7A
FB24
FB1D
FB88
FBBB
FB21
FA79
FB75
FEC1
02E2
0582
05C2
04D8
0465
04D0
0556
055D
0512
04DD
04C9
04AC
0491
04A4
04D0
04D4
04A6
0488
04AA
04EE
051C
052A
0529
0512
04E1
04B9
04BD
04C5
048B
043E
0476
053C
056A
0392
FFBE
FBDB
F9F8
FA44
FB25
FB2F
FA8E
FA4C
FAC5
FB57
FB5E
FAFE
FAC8
FAF7
FB51
FB8A
FB8D
FB5D
FB0E
FAD6
FAEB
FB34
FB55
FB2E
FB05
FB0F
FB1F
FB09
FB0A
FB61
FBAC
FB4E
FA9B
FB23
FE0E
026A
05C1
0697
05C2
0503
04FA
04FC
0498
044B
0499
052C
0552
0504
04D8
050B
052C
04E4
048D
049E
04F6
050C
04B9
0453
042D
0455
04B8
0531
0568
0513
0488
0491
0549
055C
0334
FF09
FB24
F9A2
FA56
FB5E
FB70
FAE8
FABB
FB1C
FB7E
FB7F
FB42
FAFC
FAB9
FA95
FAC8
FB3D
FB7C
FB4F
FB19
FB46
FB9A
FB8B
FB20
FAED
FB35
FB83
FB60
FB0A
FB05
FB2C
FAF2
FAA3
FB96
FEA1
02A5
056D
05EA
0519
0496
04D6
0525
04F2
048F
0482
04C2
04E9
04DB
04D7
04FA
0511
04F0
04B8
04A1
04B3
04CB
04D7
04D9
04D2
04C9
04D9
0503
0504
04A2
042F
045E
0532
056D
0399
FFCB
FBF9
FA2A
FA80
FB61
FB76
FAF0
FAC1
FB31
FBA0
FB89
FB1A
FAC9
FABC
FADE
FB2C
FB9F
FBE2
FB96
FAEB
FA8A
FAC7
FB34
FB42
FAF9
FAC9
FAE0
FB11
FB45
FB86
FB9F
FB39
FAB3
FB62
FE3C
0253
0551
05DC
04E5
0448
049F
0512
04EE
0497
04AC
0508
0512
04BA
0487
04B0
04D3
04B3
04A7
04F2
0538
050E
04B4
04B9
050F
0528
04E1
04C0
050D
054C
0505
04AC
04E6
0518
03A4
000F
FC1F
FA18
FA48
FB14
FB2E
FADD
FAF6
FB6C
FB87
FB20
FAD7
FB09
FB50
FB46
FB2D
FB61
FB9D
FB64
FADE
FAAB
FB02
FB68
FB72
FB3D
FB0D
FADC
FAA1
FAB7
FB58
FBE9
FB86
FA97
FAF3
FDD1
0204
0503
0599
04E6
049D
050B
0549
04E4
0471
048E
04FD
052A
0508
04EF
04EA
04C3
048B
049D
04FA
0524
04D5
0479
049C
051B
0553
050F
04C6
04CF
04DF
04AF
0499
04F5
050B
0378
FFF3
FC21
FA1A
FA50
FB51
FBAC
FB5A
FB2A
FB5E
FB7F
FB42
FAF9
FAFA
FB1F
FB1A
FB00
FB1D
FB69
FB81
FB43
FAF9
FAE5
FAEA
FADF
FAE1
FB06
FB10
FAD2
FAAA
FB10
FBBB
FBD8
FB66
FBCE
FE60
025E
0559
05D0
04BF
0426
049A
0515
04C9
0437
0436
04B4
04F9
04D2
04BB
04E9
04F9
04B3
048C
04E5
0554
053C
04BD
0484
04C5
0505
04F6
04E0
0504
0510
04B4
0464
04B0
04E9
0371
FFDE
FC05
FA2D
FA90
FB6D
FB5F
FAB9
FA86
FAEC
FB3E
FB28
FB13
FB44
FB6E
FB4F
FB35
FB67
FB8F
FB4A
FAE8
FB09
FB9A
FBE5
FB91
FB1D
FB0C
FB2B
FB0F
FAEC
FB3A
FBA9
FB5D
FA88
FAE4
FDC6
021F
054C
05DD
04E4
0450
04C0
055F
056F
0529
050B
050E
04F3
04DB
0508
053F
0507
0469
03F9
041E
0494
04DD
04D0
049C
0463
0432
0437
0491
04F7
04E8
0477
0467
0515
0584
042A
00C3
FCEE
FAAC
FA74
FB10
FB36
FAC5
FA72
FAA9
FB21
FB63
FB46
FAF5
FAAE
FAA9
FAF8
FB6C
FBAA
FB89
FB43
FB31
FB5D
FB8A
FB94
FB93
FB8C
FB57
FAF8
FAD6
FB33
FB9C
FB5B
FAAF
FB01
FD7D
0171
04B8
05D3
0548
04A9
04B7
04F9
04E0
04A0
04B8
0516
053E
050D
04E5
0508
052B
04F8
0498
046E
0489
049F
048D
0481
0498
04B7
04C4
04D6
0504
052B
052B
052E
054F
0502
035A
0033
FCC5
FAA2
FA40
FAC7
FB2C
FB1D
FAE5
FAC9
FAD6
FB04
FB42
FB5B
FB29
FAE1
FAEB
FB46
FB72
FB26
FABE
FABD
FB15
FB53
FB55
FB61
FB90
FB87
FB19
FABC
FAEF
FB5A
FB2F
FA8D
FAE2
FD5F
0152
049B
05D3
0577
04FA
0518
0567
054E
04DE
049B
04C0
0506
0519
04F9
04E4
0501
0525
0506
049A
0443
046F
0503
0561
0521
0496
0463
04B0
0507
04FE
04BD
04AB
04D8
0500
04FE
04D6
0437
027F
FF96
FC82
FA9C
FA42
FAA3
FADB
FADD
FB18
FB89
FBAC
FB42
FAC2
FABA
FB10
FB38
FB03
FAD4
FB06
FB6C
FB91
FB51
FAF9
FAD8
FAE6
FAF1
FAF6
FB25
FB81
FBB9
FB89
FB28
FB0D
FB55
FB84
FB3C
FB10
FC47
FF65
0330
0597
05BF
04CC
0476
051C
05AA
0540
045A
0408
047C
04E5
04B1
0455
048B
0538
0590
053C
04CA
04DD
054D
0571
050A
0488
0456
0454
0431
0409
0439
04B6
04F6
04B7
0481
04E5
0568
049B
01B7
FDC7
FAE5
FA37
FAEF
FB6D
FB07
FA70
FA81
FB24
FB9B
FB8B
FB4B
FB48
FB68
FB51
FAFD
FACB
FAEF
FB23
FB05
FAA2
FA77
FAD4
FB78
FBDF
FBD9
FBA4
FB84
FB74
FB52
FB38
FB5B
FB8F
FB56
FAB8
FAD7
FCFD
00F3
04AE
0628
056A
0457
0472
0553
059F
04FC
045F
0486
04F4
04DB
0464
0465
050A
0584
0534
048D
0469
04D9
0525
04E9
0491
0498
04CA
04B0
0465
0471
04E0
0516
04B0
042E
045F
0530
0561
03AC
002D
FC82
FA76
FA7C
FB75
FBDE
FB46
FA87
FA92
FB42
FBA4
FB49
FAD0
FAEC
FB61
FB71
FB06
FAD3
FB3A
FBA4
FB61
FABB
FA9D
FB31
FB9A
FB44
FACB
FB0F
FBD3
FC14
FB85
FAF9
FB12
FB3D
FAB4
FA1D
FB34
FEA4
02C6
0538
0551
0484
0466
0507
056D
051B
0497
0491
04F9
0539
050C
04C5
04C3
04F3
04F7
04AE
045B
0455
049D
04E3
04E7
04BA
0493
0481
0475
0483
04D5
0546
0560
04F0
047F
04C0
0572
0529
02BD
FED0
FB82
FA5C
FAE1
FB6C
FB1F
FA91
FA98
FB12
FB3A
FAE0
FAA5
FAFC
FB79
FB70
FAFD
FAE2
FB68
FBE5
FBA4
FAE7
FA94
FAFF
FB84
FB79
FB14
FB05
FB5C
FB6F
FAE4
FA51
FA70
FB01
FB18
FA95
FAB9
FCD1
007E
03D7
0550
0524
04B8
04EF
0575
0593
0534
04DA
04D7
04F7
04EF
04CC
04D4
0512
0541
0520
04CA
0492
049E
04C2
04C8
04BF
04D8
050D
0523
050A
050A
055B
05AF
057D
04D3
047E
04F6
055C
0418
00BA
FCD1
FA72
FA2C
FAC4
FAEB
FA9B
FA98
FB10
FB63
FB26
FAC5
FACD
FB1A
FB18
FABB
FA99
FB0E
FBAB
FBCA
FB5D
FAF2
FAE7
FAFF
FAE1
FAAA
FAC4
FB32
FB70
FB20
FA9C
FA92
FB1E
FB8A
FB3C
FABE
FB7D
FE4A
022C
051E
05FB
056C
04E3
04FE
053F
0523
04E9
050E
056A
055B
04C5
0454
048F
051B
0539
04D0
047A
049F
04ED
04EE
04B8
04C1
0519
0548
0500
049A
0499
04E9
04FD
04A5
0469
04CA
0558
04D7
0273
FECA
FB97
FA3A
FA95
FB61
FB8B
FB0E
FA96
FA88
FAB5
FAD1
FAED
FB34
FB78
FB62
FB07
FAED
FB48
FB9E
FB64
FACE
FA97
FAF8
FB59
FB2C
FABC
FAC4
FB4D
FB9C
FB43
FAD7
FB19
FBC6
FBDC
FB1B
FABD
FC3F
FF9C
0323
051F
055B
04EF
04DB
0522
0540
0504
04BC
04B1
04C8
04C2
049F
04A0
04DD
0518
050B
04D6
04D4
051E
0559
052F
04CD
04AC
04F0
0533
0512
04BE
04AF
04EB
04F0
0486
043B
049E
0524
0455
0171
FD95
FAE2
FA68
FB45
FBDC
FB97
FB1D
FB18
FB56
FB47
FAED
FAC7
FB02
FB2E
FAEF
FA96
FAAE
FB25
FB5A
FAFE
FA8B
FA9A
FB0C
FB3D
FAF6
FAB5
FAEF
FB5E
FB74
FB35
FB37
FBB0
FC07
FBA7
FB0F
FB98
FE01
0171
042C
0531
04F5
049C
04BB
0507
0501
04A7
0472
04AB
051A
0553
054A
0546
0566
0567
0512
04AF
04C1
054A
05A6
0556
04B8
0497
0511
056D
0521
048F
0468
04A2
0497
0426
040A
04A1
04E4
033E
FF96
FBD1
FA00
FA58
FB52
FB97
FB33
FAF0
FB1A
FB4C
FB35
FB02
FAFF
FB1A
FB09
FACA
FAA7
FACB
FB04
FB0C
FAE1
FABE
FACF
FAFA
FB09
FAF0
FAE2
FB01
FB29
FB23
FB07
FB31
FBA6
FBE4
FB84
FB29
FC3C
FF5B
0340
05B4
05D0
04D0
047E
0526
059E
051A
0449
044D
0526
05BD
0565
04B0
0488
04EC
051F
04CD
0476
049D
0502
0513
04CC
04BA
0524
0597
0586
050F
04C4
04CF
04C1
045B
0417
0480
051A
047B
01CC
FDF9
FB0B
FA37
FAD7
FB63
FB24
FAA5
FAA0
FAFD
FB22
FAE4
FABB
FAFD
FB56
FB49
FAF0
FAE5
FB5C
FBCD
FBA7
FB1A
FAD7
FB21
FB7B
FB68
FB16
FB07
FB3E
FB39
FAD0
FA9D
FB25
FBEA
FBDF
FAF5
FAB6
FCC2
00D2
04A2
0627
0579
0468
045B
0511
0572
0520
04BF
04E5
055A
057F
0532
04DD
04CD
04DA
04C4
049F
04AB
04DC
04E7
04B2
047F
048E
04BC
04C2
04A8
04C1
0518
053E
04D9
044C
0462
052F
058D
040C
0095
FCC4
FA85
FA51
FB02
FB40
FAD8
FA88
FACB
FB3E
FB45
FAE2
FA9C
FABB
FAF4
FAF3
FADD
FB08
FB66
FB93
FB60
FB20
FB25
FB4D
FB39
FAE8
FAC5
FB07
FB5A
FB5C
FB37
FB69
FBEB
FC07
FB48
FA77
FB25
FE15
0224
0524
05D7
04F8
0446
04AC
0598
05FC
059A
051F
0515
053D
0510
049D
0477
04D5
053A
051D
04AC
0481
04C3
04F9
04CB
0484
049E
0500
0527
04EE
04C2
04DE
04D5
0447
03B6
0407
0508
051A
02D5
FED6
FB66
FA39
FAE5
FBB2
FB9E
FB12
FAD7
FAF9
FAF7
FAAD
FA85
FAC4
FB18
FB0C
FAB9
FAAC
FB16
FB82
FB73
FB12
FAF6
FB48
FB8E
FB58
FAE5
FACE
FB29
FB69
FB32
FAF0
FB3C
FBD6
FBD6
FB14
FAE1
FCC2
0086
041F
05A6
0537
0478
048D
050F
0510
0488
0440
049E
0528
054E
0531
0541
0571
0549
04B8
0458
0499
0514
050B
047B
0422
0476
04FF
0502
048B
0451
04A5
04F3
04A6
0420
044F
054A
05CC
0463
0105
FD37
FAAA
F9E6
FA38
FAB5
FAF4
FB0D
FB25
FB3F
FB4F
FB56
FB55
FB49
FB32
FB18
FB07
FB01
FB0C
FB31
FB71
FBAD
FBB5
FB78
FB22
FAFE
FB21
FB57
FB59
FB32
FB3A
FBA1
FC09
FBCF
FAE2
FA33
FB12
FDE2
0190
0468
0589
0578
054D
0585
05C3
0594
0517
04CB
04D4
04D7
048D
0437
044F
04DC
0551
053D
04CD
0486
048D
0486
0439
03FF
0456
0517
057D
050B
0433
03D3
042E
04B3
04D6
04AE
0482
0405
027C
FFCE
FCF9
FB35
FABC
FAC7
FAA9
FA7E
FAB0
FB1D
FB41
FAF6
FAB0
FAC7
FAF9
FAE1
FAAE
FAE2
FB7A
FBC3
FB53
FABE
FADF
FBA9
FC24
FBC3
FB24
FB2F
FBBE
FBD5
FB1F
FA92
FB1B
FC2B
FC4A
FB28
FA70
FC09
FFD2
039D
0578
0572
0500
0512
055E
054A
04EF
04D4
0514
0548
0537
0528
055E
05A2
058C
0529
04E5
04E8
04DA
0478
0414
042B
04AC
04F8
04C0
0470
0490
04F4
04F3
046B
0404
044F
04EF
051E
04CC
04AE
0506
04D2
02CC
FF1A
FB82
F9B6
F9C2
FA5E
FA93
FA8E
FAD4
FB4B
FB5B
FADE
FA65
FA74
FADF
FB16
FAE5
FA9E
FA9D
FADC
FB21
FB55
FB7C
FB8A
FB6F
FB46
FB40
FB59
FB56
FB22
FAF7
FB0F
FB42
FB46
FB2A
FB58
FBD8
FC0B
FB6E
FAAE
FB5C
FE4B
0268
0582
0653
0585
04B8
04D1
0573
05D2
05A4
052E
04C8
049C
04BA
0519
0580
059F
0568
0520
0500
04E5
0493
042C
041A
047F
04FA
051C
04F7
04E8
04F8
04D6
046A
0425
045F
04B1
046E
03BD
03A3
049A
0570
0437
0084
FC37
F9B6
F9A2
FA9A
FB1A
FAF7
FAEC
FB46
FB8F
FB5E
FAEC
FA9E
FA77
FA4F
FA48
FAAB
FB4B
FB9A
FB63
FB19
FB2F
FB65
FB28
FA8D
FA59
FAF2
FBB7
FBCD
FB4C
FB13
FB7C
FBE2
FBB2
FB62
FBC2
FC89
FC74
FB2A
FA57
FC14
0058
049D
0669
05B6
0488
0470
0528
058A
0536
04C4
04B8
04EE
0518
053B
0570
057D
0520
0499
0473
04C4
04FE
04BD
046B
04AE
0566
05B5
0527
0451
0407
0445
0459
0409
03EB
0462
04DA
0495
03F0
040E
050A
0534
02CD
FE5D
FA8B
F96F
FA82
FB93
FB5B
FA84
FA4D
FAE0
FB75
FB89
FB61
FB50
FB36
FAE7
FAA7
FAD3
FB42
FB62
FB06
FAA7
FAB5
FAFE
FB0E
FAEA
FB03
FB77
FBD4
FBBD
FB7C
FB87
FBBB
FB97
FB21
FB09
FB9B
FC0C
FB75
FA6E
FAEB
FE15
029F
05D1
0645
0519
0466
04E5
0596
055E
0469
03BE
03F1
04A6
053C
0576
0576
055C
053C
0533
054C
0552
050B
04A0
048D
0505
0596
05A1
0512
046B
0414
0402
040F
0457
04E3
0531
04AD
03AA
035B
0455
055B
045C
00CE
FC99
FA46
FA70
FB7D
FBB7
FB0B
FA8F
FAD2
FB4E
FB59
FB04
FABF
FA9E
FA67
FA2B
FA48
FACB
FB38
FB2B
FAE5
FAE8
FB35
FB56
FB1D
FAEA
FB0D
FB42
FB21
FAD6
FAF0
FB7D
FBD7
FB97
FB40
FB7F
FC01
FBC1
FAB0
FA69
FC99
00D1
049A
05EB
051F
0429
0444
04EE
051D
04C4
04A9
052E
05D5
0600
05B3
0555
050D
04C4
0497
04D3
0565
05B4
0555
04AA
0476
04DF
053D
0506
0481
0452
048E
04B7
048E
046E
04A4
04D9
0498
0437
0480
0554
0530
02B9
FE97
FB25
FA1A
FAE6
FBA3
FB4F
FA8C
FA57
FAB8
FB05
FAF6
FAE0
FAFB
FB04
FAC6
FA93
FAD3
FB5B
FB95
FB4D
FAF5
FAF2
FB15
FAF7
FAA9
FA97
FADF
FB23
FB25
FB25
FB69
FBB0
FB8E
FB31
FB40
FBCF
FBFB
FB19
FA11
FAD1
FE25
0282
056D
05EA
052D
04E7
0572
05E3
058E
04DD
049E
04F4
0555
0550
0507
04D6
04D9
04E5
04D8
04B6
0497
0494
04C8
052E
057D
055B
04D3
046D
0491
0503
0525
04D2
0495
04D9
0533
04EF
042E
03F7
04BF
0555
03E4
0029
FC1C
FA0E
FA58
FB59
FB82
FAE0
FA7C
FAC3
FB23
FB10
FAC3
FAB9
FAEC
FAFC
FAD9
FAD9
FB20
FB55
FB30
FAF3
FB0E
FB72
FB99
FB47
FAD3
FAAA
FAC5
FAE6
FB10
FB64
FBAE
FB82
FAFF
FAEA
FBAA
FC80
FC4F
FB48
FB2B
FD66
013C
045C
0548
04B3
0457
04DF
0580
0567
04D8
04AA
050F
0565
0534
04C9
04B8
050B
0547
051D
04C3
0493
049F
04B8
04BF
04B8
049E
0469
0442
0470
04E7
0535
0503
0495
0471
0499
0480
03EE
0392
042A
0529
04D6
0224
FE29
FB38
FA8B
FB36
FB90
FB1D
FAAE
FAE4
FB50
FB39
FAB5
FA80
FAE5
FB5E
FB62
FB15
FAF5
FB18
FB2D
FB15
FB0F
FB45
FB81
FB82
FB60
FB54
FB4B
FB15
FAE7
FB3B
FC05
FC74
FBED
FAFF
FAC9
FB79
FBF2
FB5F
FAA7
FBB1
FF14
031F
057E
058C
04A0
0442
04A9
0518
051D
04F5
04ED
04E9
04BA
048F
04AF
0500
0514
04C7
0477
047F
04BC
04CB
049C
0484
04B8
04FD
04FD
04BF
048E
0488
0489
048A
04B8
050A
0508
046B
03C9
0425
057A
0627
0466
005D
FC4C
FA5E
FA9D
FB57
FB4A
FAD1
FADC
FB70
FBB2
FB3A
FA9B
FA8E
FAFE
FB4C
FB3D
FB2D
FB59
FB85
FB70
FB4C
FB6B
FBAC
FBAB
FB5D
FB22
FB24
FB15
FABB
FA7A
FACD
FB6A
FB7F
FAE0
FA79
FB0E
FC00
FBFA
FAEC
FA98
FCAF
00AA
0426
055C
04C9
0433
0487
053B
057C
054A
052F
0553
055C
0510
04B2
049C
04C5
04E1
04C9
0495
045A
041C
0401
0446
04E5
056F
057E
0531
04FD
050A
0506
04C3
049B
04F1
0569
0532
043D
03AD
047E
05DF
059A
0274
FDD3
FA80
F9E4
FAE7
FB93
FB43
FACE
FAEC
FB47
FB3D
FAE4
FAD1
FB22
FB5A
FB2E
FAFF
FB3A
FBA2
FBA3
FB2F
FAD0
FAE3
FB23
FB29
FB09
FB10
FB35
FB32
FB11
FB2A
FB7B
FB83
FB0C
FAC3
FB67
FC77
FC7F
FB13
F9EC
FB4E
FF60
03BC
05E4
05A3
04B4
047A
04C6
04D6
04A5
04C1
0535
0557
04C8
0415
03FE
0486
04FE
0500
04D9
04F4
0537
0538
04EE
04B9
04CF
04ED
04BE
0455
040A
0401
041F
0460
04E1
0576
0594
04F2
0431
0452
0551
05AA
03C3
FFCA
FBCD
F9CC
F9F1
FAD6
FB45
FB3B
FB41
FB73
FB78
FB3D
FB1E
FB4C
FB7D
FB6B
FB4F
FB82
FBD6
FBC0
FB2E
FAC5
FB0D
FBA4
FBB8
FB22
FAA1
FADC
FB91
FC04
FBF0
FBA6
FB6C
FB31
FAFC
FB21
FBB3
FC09
FB76
FA77
FAAD
FD30
0125
046D
05A5
0540
04A6
04A3
04F8
051D
04F8
04C8
04B7
04BF
04DC
050D
0529
0503
04A6
0461
0461
0480
047E
045F
0463
049B
04CB
04C0
04A3
04C1
0512
0532
04ED
0493
048C
04BE
04AB
0437
03F6
0463
04E8
041F
015B
FDAC
FB03
FA5A
FAEE
FB5F
FB34
FAFB
FB33
FB98
FBA1
FB4A
FB03
FB03
FB13
FB0B
FB1C
FB72
FBC6
FBB5
FB51
FB0E
FB23
FB45
FB29
FAFB
FB0C
FB47
FB50
FB24
FB2E
FB91
FBCC
FB71
FAE5
FAE9
FB75
FBA6
FB14
FACC
FC50
FFAF
0335
0528
0579
055D
059B
05D7
058A
04ED
04A7
04D3
04F0
04AF
0460
0463
048C
046C
0408
03E1
0445
04DF
0538
0546
0556
0580
0585
053C
04DA
04A0
0485
045E
0440
0462
049E
0476
03D7
0385
0446
059D
05CC
0386
FF71
FBB1
F9EB
F9F4
FA81
FAB5
FAAF
FACA
FAFA
FB0B
FB18
FB58
FBA3
FB8D
FB16
FAD4
FB2E
FBC4
FBE0
FB6E
FB14
FB43
FBA6
FBAC
FB55
FB19
FB25
FB29
FAEF
FABD
FAE0
FB28
FB32
FB1D
FB61
FBFA
FC34
FB9B
FAB9
FA72
FAD0
FB19
FB1B
FBCB
FE19
0185
0459
0578
0558
0521
0548
056F
054B
0506
04CD
047F
0419
0401
047F
0529
053F
04AE
043E
0488
052E
0564
0507
04B1
04C5
04F8
04E6
04BC
04E3
053F
053B
04AA
0425
044B
04EE
055D
0547
04F7
04B4
046C
0420
043B
04F6
0586
048A
018D
FDD5
FB44
FA94
FAEA
FB1B
FAEE
FADE
FB27
FB6F
FB66
FB34
FB1C
FB11
FAE8
FAD4
FB30
FBD8
FC13
FB77
FA8C
FA43
FAC8
FB55
FB30
FA95
FA46
FA8D
FAFD
FB2E
FB3E
FB78
FBC2
FBC6
FB7F
FB42
FB38
FB39
FB3A
FB74
FBDD
FBDD
FB18
FA72
FB89
FED8
02C6
0513
052C
047D
047F
051F
055A
04EB
048F
04D2
054B
0557
0510
0501
0535
052C
04C6
049D
051B
05BE
05B3
04FE
0470
0491
0501
0525
0500
04F8
051F
051B
04D5
04A5
04C0
04DB
04B1
0489
04BA
04F7
04AC
0410
0428
0541
05EE
044F
005F
FC5E
FA8E
FAF2
FBC1
FBAF
FB12
FADD
FB2B
FB57
FB12
FAC3
FACD
FAFD
FAF6
FACB
FACF
FAFA
FAED
FA9A
FA74
FAD8
FB7D
FBC7
FB86
FB1E
FAF5
FB03
FB14
FB21
FB3E
FB51
FB2F
FAF8
FB04
FB5C
FB97
FB73
FB49
FB8A
FBE8
FB8E
FA7B
FA22
FC13
000E
03E6
05A0
0555
04AD
04C6
0538
0528
04A2
0466
04BB
0520
0527
050C
052F
0560
0528
04A0
0474
04F3
058D
0593
0515
04B4
04B9
04D7
04C4
04A4
04AC
04B6
0489
0454
0473
04CD
04DE
0489
0459
04AB
0503
04C8
045C
04B6
05BB
05B6
032C
FEE9
FB7D
FA8B
FB43
FBC5
FB64
FAED
FB07
FB48
FB0C
FA8C
FA7C
FAEC
FB3A
FB0C
FACC
FAE8
FB1D
FAED
FA7A
FA66
FADE
FB57
FB5A
FB25
FB3A
FB94
FBBE
FB8F
FB5B
FB5A
FB4C
FB06
FAE6
FB49
FBCD
FBB2
FB04
FAB3
FB40
FBD0
FB43
FA1A
FA66
FD72
01FB
054C
060B
0546
04CF
052F
05A1
058A
0537
0527
0540
0523
04E1
04DB
050B
04FF
048E
043A
047C
050D
053B
04E0
0490
04C0
0524
052E
04DB
04A6
04C2
04E6
04D6
04CA
0502
053F
0525
04E5
050D
0597
05C5
052F
048F
04C8
054A
0446
00DE
FC9C
FA12
FA1E
FB36
FB7C
FAC9
FA44
FA88
FB07
FB27
FB26
FB79
FBDA
FBA7
FAF5
FA95
FAE8
FB4D
FB1E
FAAD
FACA
FB77
FBD8
FB6D
FACA
FABE
FB3D
FB90
FB76
FB5D
FB8B
FB9B
FB38
FAC1
FAC1
FB0B
FB0A
FAC7
FAF4
FBAC
FBF3
FB1B
FA46
FB87
FF4F
037A
058B
054B
0499
04E0
05A6
05C0
051C
04A7
04CF
0503
04C0
0468
049A
0525
054B
04DC
0476
049D
0507
0521
04E6
04CF
0506
052D
04F3
0490
046B
048D
04B2
04C6
04E4
04F7
04B9
0438
0400
0468
0500
0518
04C3
04D4
057E
0585
0366
FF54
FB81
F9FE
FAAC
FBAC
FB9F
FAEE
FAC2
FB50
FBBD
FB7B
FB03
FB06
FB68
FB74
FAF3
FA75
FA7F
FAE0
FB19
FB1D
FB3E
FB92
FBC1
FB96
FB4E
FB3D
FB52
FB47
FB24
FB2C
FB65
FB7F
FB5E
FB4C
FB74
FB88
FB46
FB05
FB49
FBC6
FB95
FAA8
FA86
FCCB
00FD
04A0
05C4
04F9
0443
04A5
0558
0551
04AF
0453
048D
04E5
04FB
04FE
052A
0546
0510
04BD
04B2
04E1
04DE
0489
0445
045F
04A7
04C5
04BD
04CD
04EE
04DC
049E
0499
04EE
0525
04D4
0450
043F
0499
04AB
0432
03F4
04B8
05D0
0565
027A
FE47
FB26
FA52
FAFE
FBA0
FB8E
FB2D
FAFE
FAFF
FAF9
FAF9
FB26
FB62
FB5A
FB01
FAAE
FAB6
FB00
FB3B
FB49
FB50
FB6B
FB80
FB78
FB70
FB85
FB9C
FB7B
FB25
FAE1
FADD
FB01
FB2C
FB6D
FBC8
FBEF
FB90
FAF0
FAC3
FB37
FB8C
FB17
FA8F
FB97
FECA
02A2
04DC
04DE
0423
0443
0532
05C8
057F
04F2
04CC
04E8
04D2
049B
04AD
050D
0539
04F7
04A9
04B2
04DE
04C7
0485
048D
04EB
0526
04F2
049E
049B
04D1
04D2
0494
047E
04C0
0504
0508
050C
0546
054E
04A1
03B8
03CF
0531
0639
04C5
00B6
FC66
FA58
FAC7
FBDF
FC00
FB35
FA81
FA6C
FAB3
FAFC
FB44
FB93
FBB4
FB84
FB41
FB3C
FB63
FB60
FB2A
FB17
FB54
FB8F
FB68
FB02
FAD6
FB06
FB32
FB10
FAD7
FADF
FB12
FB1B
FAFD
FB17
FB7E
FBBD
FB7A
FB18
FB35
FBA1
FB81
FAB5
FA93
FC98
0075
040A
057E
0505
0448
0462
04FA
053C
0509
04D5
04D2
04C6
049D
0496
04D0
0501
04E4
04A8
04AB
04E2
04EE
04C2
04CE
0549
05BB
058A
04DE
047F
04CB
0542
053C
04CB
0483
049F
04C5
04B1
049A
04BA
04C8
0472
0419
047A
0562
0559
0314
FF2B
FBC8
FA87
FAFB
FB8E
FB5C
FAD4
FAAC
FAE7
FB15
FB1F
FB42
FB83
FB91
FB56
FB30
FB63
FB9F
FB75
FB01
FACB
FAF4
FB02
FAA5
FA4C
FA98
FB5F
FBCC
FB7B
FB01
FB0D
FB82
FBBC
FB8D
FB59
FB5B
FB48
FAF3
FACB
FB2F
FBA1
FB4E
FA85
FAEC
FDAD
01CF
04FD
05DC
0528
047B
048C
04EE
0520
0523
051A
04E7
0482
0446
0482
04F7
051B
04E0
04BC
04EE
0523
0500
04B5
04B9
0508
051B
04B4
0449
0461
04D6
050F
04E2
04B9
04E4
051C
04FD
04AD
04A0
04D7
04D3
0469
0430
04B3
054E
047F
0195
FDBC
FB06
FA66
FB00
FB65
FB16
FAA2
FA9C
FAEC
FB2D
FB44
FB55
FB5E
FB3D
FB0B
FB0D
FB48
FB6B
FB50
FB45
FB8E
FBDC
FBA7
FB03
FAAD
FB0E
FB93
FB6E
FABD
FA66
FACB
FB4E
FB4E
FB1B
FB56
FBD2
FBC2
FB11
FAAE
FB2A
FBB6
FB40
FA66
FB32
FE93
02DC
0571
058D
04AD
046D
04E6
0545
0540
0538
0550
0527
04A4
044E
0486
04E4
04D5
0483
048B
04F2
0513
04A7
044B
04A5
055F
0590
050C
04A0
04E5
0561
0547
04B4
047E
04F0
0556
050F
0484
0483
0508
053A
04BC
044B
0496
04E4
0398
003D
FC77
FA72
FAA9
FBA7
FBE0
FB45
FAC9
FAF1
FB51
FB6A
FB5D
FB7D
FBA2
FB60
FAC6
FA68
FA9A
FB03
FB30
FB34
FB60
FB9C
FB83
FB17
FAEC
FB53
FBC5
FB8E
FAD3
FA6C
FAB4
FB17
FB01
FABC
FAE3
FB5B
FB82
FB3C
FB29
FB8C
FBB5
FB23
FAD4
FC7D
0041
0404
058E
04F4
0426
0473
0548
0575
04EA
048F
04D4
0535
0525
04D3
04BA
04D3
04C8
04A2
04C2
052E
056F
053A
04DD
04C8
04EB
04E0
0495
046F
04A7
04ED
04E6
04B9
04CD
0523
0551
0529
04F6
04F6
04F1
04A9
0478
04EA
059E
0521
0265
FE4B
FB1B
FA49
FB11
FB9B
FB18
FA5D
FA71
FB28
FB86
FB24
FAA4
FAB1
FB23
FB5A
FB2E
FB09
FB32
FB68
FB61
FB3D
FB3D
FB4D
FB2A
FAE0
FAC9
FAFE
FB30
FB21
FB11
FB53
FBB6
FBB9
FB58
FB1F
FB56
FB87
FB31
FA9C
FA7C
FAE3
FB2D
FB0B
FB03
FB88
FC03
FB90
FAA8
FB2F
FE48
02A4
05AA
062D
0556
04E7
0538
056B
0507
049F
04D4
055F
0586
051D
04A3
047F
0499
04C1
04FC
0548
055A
04FA
0473
0455
04B9
0516
04F5
048B
0462
0495
04C0
04AB
049F
04E7
0545
053F
04DC
04A5
04E1
052B
050D
04B3
04A6
04EC
04F2
047F
043A
04B1
051F
03E7
0091
FCBA
FA91
FA98
FB61
FB72
FAD6
FA86
FAD6
FB28
FB02
FABE
FADA
FB2F
FB46
FB20
FB2D
FB82
FBAB
FB65
FB17
FB3F
FBAE
FBCA
FB77
FB40
FB7E
FBC9
FB9D
FB25
FAF9
FB35
FB62
FB3A
FB0F
FB3C
FB86
FB7C
FB33
FB2F
FB8D
FBC2
FB78
FB26
FB5E
FBC7
FB7C
FA8F
FA7E
FCB3
00B1
0452
05E1
059A
04FB
04F5
053F
053E
04EE
04BA
04C6
04CD
04AB
049E
04D9
0523
0519
04BA
046D
0477
04A3
04A0
047C
0485
04C3
04DF
04A9
0461
0468
04B7
04F7
04F5
04D7
04BE
048E
0438
0401
0431
049B
04C7
04A7
04A4
04E8
04F8
0478
03FA
0458
053A
04EC
0232
FE02
FAC8
F9E9
FA96
FB33
FB3C
FB4A
FBA9
FBD0
FB4E
FA99
FA71
FADD
FB33
FB1D
FAFA
FB31
FB8C
FB95
FB51
FB30
FB59
FB84
FB76
FB54
FB5B
FB7D
FB88
FB75
FB6A
FB63
FB38
FAF7
FAF8
FB64
FBDE
FBF5
FBB8
FB95
FBB1
FBAE
FB54
FB06
FB48
FBDC
FBE2
FB0B
FA71
FBAF
FF13
0305
0575
05CF
0538
0507
0568
059F
0545
04D2
04D7
0529
0528
04B1
0453
0482
04FE
0535
0501
04BF
04B7
04C8
04B3
0480
0460
0462
0466
046B
0489
04B6
04C6
04B8
04C6
0503
0529
04FF
04B8
04AB
04C4
049F
0440
042E
04AB
051E
04CF
0416
0417
0507
055D
0361
FF61
FBAB
FA34
FABB
FB84
FB70
FADD
FAA3
FAD3
FAE7
FAAA
FA77
FA9F
FB00
FB4B
FB68
FB78
FB93
FBB6
FBD7
FBE7
FBCA
FB72
FB0C
FAE4
FB0F
FB44
FB36
FAF2
FAC9
FAE3
FB13
FB2A
FB38
FB66
FB9C
FB97
FB52
FB28
FB5E
FBB4
FBA3
FB25
FAE2
FB4F
FBEB
FBC9
FB03
FB18
FD68
0162
04CB
05F5
0562
04DD
0546
05D6
0592
04AF
042E
046F
04DE
04EA
04BC
04C2
04F4
04F3
04BC
04AF
04EC
0516
04ED
04BA
04D7
0513
04FE
04A2
0487
04F1
057D
05A9
057D
0557
054B
0516
04B4
0489
04C3
04F6
04B6
044A
0453
04D0
050D
04B2
045F
04C7
0554
046B
0148
FD3F
FA9C
FA5E
FB6A
FBFD
FB89
FADF
FAD4
FB49
FB91
FB6F
FB3E
FB4F
FB74
FB5C
FB18
FAFE
FB22
FB3E
FB26
FB0A
FB22
FB48
FB23
FAB4
FA64
FA83
FAE4
FB22
FB1F
FB10
FB15
FB17
FB09
FB11
FB3E
FB61
FB57
FB48
FB5E
FB78
FB5C
FB39
FB78
FBFB
FBF3
FAFF
FA37
FB66
FEF0
0303
0550
0550
046D
041C
046C
049A
0468
0453
04AA
050C
0505
04B6
0490
04A7
04B2
0499
049C
04DF
052A
0537
0516
0508
051F
052F
0524
0520
0537
0546
052E
0518
0534
0559
0530
04B4
044F
044D
0478
0473
0459
049C
0537
057D
04FC
0453
0499
05BF
061C
0410
0007
FC4F
FAC9
FB2A
FBBC
FB7A
FAE7
FAE3
FB56
FB82
FB38
FB0E
FB69
FBDB
FBC6
FB42
FAE9
FAF2
FAFF
FAC9
FA93
FAB4
FB01
FB18
FAFE
FB19
FB77
FBA4
FB52
FADC
FABD
FADE
FAC8
FA7A
FA76
FAEF
FB64
FB52
FAFB
FAFF
FB55
FB51
FAC6
FA77
FAF0
FB76
FAEC
F9B5
F9DF
FCD9
017D
04FD
05CC
04EF
0465
04D4
054F
0510
0482
0474
04E7
0525
04DF
048F
04B5
0526
0556
0523
04E9
04E5
04F0
04D7
04BF
04DE
050F
04FA
04A1
0468
0488
04C0
04BE
04A7
04DA
0557
05B0
05A6
0581
058F
05A1
055E
04F1
04E1
0533
053F
04B9
045E
04FA
05DF
0529
01EB
FDA4
FAE7
FAB0
FB99
FBC7
FAF9
FA44
FA57
FABE
FACF
FAA2
FAC0
FB3D
FBA0
FB94
FB50
FB2B
FB2E
FB32
FB35
FB4C
FB5A
FB2D
FAD3
FAA0
FABC
FAF3
FB09
FB10
FB3A
FB71
FB64
FB03
FAA8
FA9E
FAC2
FABC
FA92
FA9B
FAE6
FB0A
FAC9
FA99
FB0C
FBD9
FBF9
FB13
FA6F
FBD9
FF89
0396
05D0
05DA
0521
04EE
0529
0512
0493
044E
049E
051A
0541
0520
0514
0529
0523
0500
0507
053D
0540
04D7
0460
0450
0493
04BB
04B5
04DF
0557
05A7
0569
04EF
04E0
054D
0596
055E
050E
051E
054E
0511
0488
046E
04F5
054B
04C1
03EE
040B
0514
054F
0329
FF34
FBBE
FA74
FADC
FB5A
FB1E
FAA8
FAAB
FB0F
FB40
FB15
FAEB
FAFF
FB1A
FAFE
FAD1
FAE1
FB1F
FB34
FB05
FADD
FAF7
FB29
FB2F
FB1C
FB36
FB7C
FB8B
FB35
FAD5
FADC
FB30
FB5A
FB38
FB28
FB59
FB77
FB34
FAE3
FB09
FB8A
FBBA
FB65
FB2E
FB92
FBEC
FB47
FA19
FA59
FD4F
01CD
052B
0603
054A
04C9
0513
0576
055F
0519
0518
053B
051E
04D3
04C5
0509
0543
0533
0508
0500
0503
04D8
0497
0492
04D8
0510
04F5
04B0
0493
04A2
04A1
0482
047E
04B4
04EE
04F1
04D4
04D3
04E4
04BD
0457
0421
047B
0514
053A
04D7
04A6
052D
059D
0462
00F6
FCD5
FA3B
F9F7
FADB
FB46
FADF
FA75
FAA1
FB0E
FB2C
FAFE
FAEA
FB00
FAF7
FABD
FAA7
FAE6
FB34
FB37
FB08
FB05
FB3B
FB50
FB1A
FAE2
FAF7
FB34
FB44
FB22
FB0E
FB1C
FB1C
FB06
FB12
FB5A
FB94
FB79
FB40
FB58
FBB4
FBC0
FB45
FADA
FB17
FB9D
FB7B
FAA6
FA80
FC78
0049
03FF
05CB
05A2
04E1
04B5
0521
057C
0573
0542
0532
053E
0538
0517
04FD
04F4
04E8
04D1
04CF
04F7
0523
051E
04EC
04CD
04E6
0514
051C
04EF
04AA
046B
044A
0460
04B0
0503
050F
04D2
049F
04B1
04CB
0497
0443
0458
04E3
0538
04DF
0468
04B8
058B
0542
02A0
FE73
FB06
F9E2
FA79
FB2B
FB23
FACD
FACD
FB1A
FB41
FB1A
FAE4
FAD7
FAE9
FAF9
FB08
FB20
FB28
FAFF
FAB5
FA89
FAA2
FAE5
FB1D
FB32
FB31
FB32
FB42
FB60
FB80
FB87
FB60
FB1D
FAF9
FB29
FB8A
FBB9
FB81
FB30
FB36
FB8B
FBB0
FB67
FB11
FB1C
FB4F
FB16
FAB3
FB7B
FE69
028C
058F
0616
0513
047E
0516
05EB
05E6
0525
0491
0494
04CC
04CC
04B2
04C8
0501
051D
051B
052E
0556
0558
051A
04D7
04CD
04FD
0534
0548
0532
04FC
04B8
048A
0492
04C3
04E0
04BE
0478
044C
0452
046A
0472
046E
047F
04B7
04F6
04FD
04BE
047F
048D
04C5
04B5
0451
0432
04C0
053B
0420
00E0
FCEA
FA77
FA49
FB15
FB40
FA9E
FA20
FA4D
FAB0
FAC1
FAA4
FACA
FB29
FB56
FB2B
FAFB
FAFD
FAFA
FAB6
FA67
FA6D
FAC9
FB21
FB3C
FB2B
FB11
FAFE
FB00
FB26
FB65
FB96
FBA1
FB96
FB8D
FB7E
FB4F
FB0F
FAEE
FAFC
FB17
FB26
FB35
FB45
FB40
FB2E
FB42
FB82
FBB2
FBB3
FBB9
FBD8
FBB1
FB00
FA88
FBC1
FF2B
033F
05B4
05D2
0500
04DA
0570
05CA
0589
053A
054A
056A
0537
04E6
04E2
051D
051B
04BE
0473
0489
04BC
04B0
0481
048B
04D3
050A
0502
04DA
04B5
049D
04A4
04DB
0529
054D
0523
04CB
0480
0458
0447
0457
0492
04CD
04CE
04A6
04A4
04CF
04D4
049E
0483
04A9
04B2
0461
043A
04C1
0541
040E
0088
FC5A
F9FB
FA10
FAF8
FB07
FA57
FA04
FA5E
FABC
FAB9
FABB
FB15
FB75
FB6B
FB20
FB11
FB46
FB4E
FAFD
FABC
FAE2
FB30
FB38
FAFE
FAD3
FACF
FAD4
FADF
FB0A
FB40
FB4E
FB33
FB23
FB38
FB50
FB4C
FB42
FB50
FB64
FB58
FB3E
FB42
FB50
FB2D
FAF2
FAFC
FB46
FB60
FB31
FB40
FBC4
FC03
FB5D
FAB9
FBFC
FFB3
03ED
0618
05C1
04BE
04AC
053C
054E
04C9
0482
04CF
0526
051E
0506
053A
057E
0561
04FE
04D9
0513
053D
0508
04BC
04B7
04DF
04E3
04C4
04BB
04C9
04C2
04AB
04AB
04BB
04B3
048E
047E
049A
04BA
04B5
049B
0495
049B
048F
0485
04A8
04D2
04B5
046D
046E
04B8
04BA
044F
043E
0502
057F
03DB
FFE2
FBC6
F9F5
FA84
FB6D
FB33
FA5E
FA28
FAA6
FB08
FAF9
FAEA
FB19
FB2B
FADC
FA80
FA87
FAD7
FB04
FAF8
FAFF
FB33
FB45
FB07
FAC3
FACB
FB03
FB23
FB2D
FB4B
FB6B
FB60
FB3C
FB3D
FB69
FB88
FB7A
FB62
FB64
FB6D
FB60
FB4D
FB56
FB62
FB45
FB1F
FB36
FB72
FB73
FB47
FB68
FBCF
FBB1
FAC9
FA6C
FC67
00A6
04C1
065B
058F
0470
0470
0511
053D
04EC
04D4
0520
0547
0506
04C0
04D0
0507
0512
04FD
050A
0538
0542
0518
04F2
04F5
04F5
04D3
04B7
04C6
04D8
04BD
0491
0487
048D
0474
044E
0456
0494
04CD
04D6
04C3
04AE
048B
0450
0426
043D
0473
0489
048C
04B1
04CA
0473
03EC
0419
051B
0572
0367
FF41
FB65
F9EE
FA99
FB7D
FB72
FAFB
FAF7
FB4A
FB55
FB0C
FAEF
FB1D
FB30
FAEF
FAA9
FAAF
FAE4
FAFD
FAF5
FB00
FB25
FB2F
FB08
FADE
FADD
FAEE
FAFA
FB13
FB45
FB63
FB4F
FB33
FB41
FB61
FB5A
FB34
FB26
FB40
FB56
FB52
FB57
FB84
FBB5
FBB5
FB94
FB82
FB74
FB47
FB32
FB8C
FC0A
FBD8
FAED
FAB6
FCB9
009C
042F
059F
0531
048B
04AB
0527
0547
0515
0503
051D
051A
04FA
0502
0534
0542
050C
04D1
04CA
04D9
04C5
0498
0493
04C9
050A
0524
0520
0512
04F7
04D2
04C5
04D5
04DC
04C9
04C0
04D8
04E1
04AE
046A
045F
0484
048C
0464
0452
0483
04B9
04AF
0496
04C2
0501
04D2
0459
0467
051B
0518
02E4
FEE6
FB5D
FA15
FAB4
FB7B
FB61
FAD2
FA9A
FACB
FAFC
FB0C
FB24
FB40
FB34
FB10
FB11
FB35
FB36
FAFF
FAD2
FAEE
FB2E
FB40
FB16
FAF1
FAFA
FB0F
FB01
FADD
FAD2
FAEB
FB14
FB39
FB49
FB36
FB17
FB1E
FB4B
FB61
FB49
FB3D
FB70
FBAA
FB91
FB3B
FB24
FB76
FBB3
FB74
FB1E
FB55
FBCC
FB84
FA82
FA79
FCF9
014C
04E6
0605
0546
047F
0497
050C
052C
0503
04F6
0506
0500
04F2
0505
051B
04FE
04D0
04DE
0518
051B
04C3
046D
0472
04AE
04BA
0487
0472
04AE
04F4
04EF
04B0
0485
0488
0499
04A2
04A7
04AA
04AE
04C0
04D7
04D0
04AB
04A4
04E2
0525
0505
0494
045A
0492
04B2
043B
03B7
0428
054A
0539
028A
FE3E
FAF1
FA20
FAF0
FB96
FB61
FAE9
FACD
FAED
FAF2
FAE6
FAF8
FB12
FB0E
FB0F
FB3E
FB6C
FB5B
FB2D
FB3A
FB78
FB84
FB3A
FAF5
FB0D
FB59
FB6F
FB44
FB31
FB60
FB8A
FB73
FB44
FB3A
FB43
FB32
FB19
FB21
FB3E
FB4B
FB55
FB75
FB8C
FB70
FB44
FB60
FBBB
FBD8
FB81
FB41
FB9D
FC0F
FB9E
FAA0
FAF9
FDF4
0256
0575
0604
0520
0495
04E2
0546
0538
0503
0508
0519
04F0
04B8
04BC
04DC
04D0
04AA
04B0
04D3
04CC
0498
048F
04D2
0513
0501
04B8
0495
04AD
04C2
04B7
04BB
04E9
050A
04EB
04AE
048C
0481
0477
0477
0488
0481
0451
0436
0467
04AD
04A5
0461
0463
04C6
04EB
0467
03EC
046C
055C
04C1
018F
FD42
FA70
FA0A
FACE
FB30
FAFD
FAE3
FB1E
FB46
FB24
FB07
FB1F
FB24
FAE8
FAC4
FB03
FB5A
FB59
FB20
FB1D
FB4B
FB3E
FADD
FA97
FABD
FB0B
FB17
FAF4
FB0F
FB75
FBB4
FB8C
FB4C
FB50
FB71
FB5D
FB21
FB0C
FB33
FB6C
FBA0
FBD0
FBE1
FBB7
FB75
FB5C
FB6D
FB5C
FB22
FB27
FB99
FBD5
FB36
FA6D
FB47
FE8E
02C2
0582
05F6
0542
04D4
04F7
0523
0518
0511
052E
053E
0527
051D
0536
0533
04F0
04B1
04BA
04DE
04D8
04C6
04E9
0525
051E
04CB
048B
0498
04B5
049E
0480
04AE
050A
051A
04BB
0464
046D
049C
0498
047C
048D
04B5
04AF
048A
0491
04C6
04DB
04BA
04A8
04C4
04B5
044F
0424
04CE
0599
04BE
0173
FD35
FA65
F9DD
FA82
FAEC
FAD8
FACD
FB09
FB41
FB3B
FB1D
FB0F
FAFA
FAD0
FAC4
FAF3
FB25
FB18
FAEE
FAF1
FB22
FB4B
FB5B
FB6B
FB78
FB65
FB37
FB29
FB54
FB87
FB89
FB6B
FB60
FB5F
FB2B
FACF
FAAC
FAED
FB43
FB5F
FB5C
FB78
FB9D
FB95
FB73
FB73
FB82
FB5B
FB0F
FB1B
FB96
FBC8
FB1D
FA6A
FB71
FECF
02EA
056F
05AC
04DD
0477
04BE
0519
0528
0517
051F
052B
0514
04EA
04C7
04A8
0486
0485
04BC
0503
0517
04F6
04CD
04B2
0498
047D
0476
048A
04A9
04C4
04DC
04ED
04E8
04CF
04C6
04EC
051F
051A
04D0
0483
0467
0475
0493
04BD
04D9
04B9
046D
0460
04BF
0511
04BC
040A
0402
04FD
05AD
0440
0091
FCA1
FA93
FAA1
FB63
FBAC
FB87
FB7C
FB97
FB82
FB2D
FAED
FAF1
FB0E
FB19
FB2A
FB59
FB7C
FB65
FB36
FB3B
FB71
FB87
FB57
FB11
FAF5
FAFF
FB04
FAFB
FB05
FB30
FB56
FB57
FB48
FB4F
FB61
FB51
FB1F
FB09
FB37
FB7C
FB8D
FB6C
FB71
FBC8
FC03
FB84
FA81
FA55
FC55
003E
0410
05D8
0574
046C
0427
04A9
050D
04E2
048D
0483
04B0
04BF
04AA
049D
0499
0477
044C
045B
04A9
04E2
04C7
048B
0484
04B4
04CE
04BC
04BB
04E5
04F2
04AC
045B
046D
04D6
0516
04E6
048D
0467
0464
044A
0438
0488
051D
0555
04E5
0477
04D8
059F
0532
0274
FE49
FAEC
F9D4
FA7E
FB4D
FB52
FAE6
FABF
FAFE
FB42
FB53
FB58
FB6E
FB72
FB4A
FB23
FB35
FB69
FB75
FB49
FB25
FB36
FB52
FB3E
FB0B
FAFD
FB1B
FB2D
FB21
FB34
FB8D
FBE5
FBD8
FB72
FB25
FB31
FB59
FB53
FB33
FB34
FB42
FB16
FAD1
FAF0
FB80
FBBF
FB19
FA51
FB1A
FE3A
0260
0547
05E0
051C
0486
04A6
04E7
04C7
047D
047C
04B7
04CD
04A1
047F
04A5
04ED
050F
0502
04F4
04F2
04DA
049B
045B
0441
0445
044A
0450
0463
0470
0455
0428
0432
0492
0502
052A
0506
04D9
04BF
0491
044A
0438
048F
04F4
04E4
0489
04A3
0564
05A6
03EB
0036
FC64
FA74
FAA2
FB7D
FBB0
FB3B
FAEB
FB16
FB5B
FB5A
FB30
FB25
FB34
FB2C
FB0B
FB03
FB27
FB4E
FB53
FB43
FB37
FB28
FB11
FB0D
FB36
FB61
FB50
FB11
FB02
FB50
FBA7
FB9B
FB40
FB19
FB66
FBCB
FBD7
FB9E
FB85
FB92
FB64
FAE8
FAAE
FB26
FBC7
FB96
FAA8
FA8E
FCBF
00BB
0442
058E
04F1
041C
041C
0496
04C1
0490
047E
04B5
04DF
04C8
04A9
04C1
04E7
04CF
0483
045D
047E
04AB
04B7
04BA
04D4
04E0
04B3
0481
04A4
0509
052E
04C8
043A
0413
0458
0487
045A
0423
0439
0470
046A
0441
0469
04E9
0522
04B7
0447
04AC
058F
0549
02A3
FE77
FB15
FA00
FAA7
FB6A
FB79
FB49
FB77
FBD7
FBE4
FB96
FB62
FB79
FB87
FB41
FADF
FACB
FB08
FB39
FB33
FB27
FB38
FB35
FAF7
FABD
FADE
FB44
FB7C
FB59
FB2E
FB4D
FB8D
FB98
FB78
FB84
FBC0
FBC4
FB61
FB04
FB1F
FB79
FB80
FB35
FB2C
FB95
FBBD
FB10
FA5E
FB5F
FEBA
02F0
05B1
061A
0539
0488
046F
0471
0446
0438
048B
04F5
0504
04BD
048B
04A4
04D4
04DE
04D6
04E2
04E7
04AE
044C
0427
047C
0507
054A
051B
04C1
0487
0475
0476
0499
04EC
053C
053C
04F4
04C2
04D8
04F1
04BF
0470
0470
04BA
04CA
0475
0450
04CA
050B
0388
FFFC
FC33
FA5C
FABD
FBA8
FB9D
FAD2
FA6C
FAC8
FB32
FB21
FAED
FB10
FB55
FB39
FAD6
FAC4
FB31
FB94
FB74
FB11
FAFD
FB49
FB7F
FB58
FB18
FB13
FB33
FB2F
FB04
FAEC
FAF5
FAF4
FAE2
FAEE
FB28
FB50
FB2D
FAEB
FAE9
FB34
FB77
FB7D
FB81
FBBB
FBD9
FB58
FA85
FAB6
FD13
011B
04BF
0632
0588
0468
0433
04CF
0540
0517
04CC
04D6
04FC
04D0
0471
0462
04BC
0501
04CF
046D
0460
04AA
04D5
04B2
0495
04C3
0500
04F7
04C2
04BD
04F0
0510
04F9
04E0
04F0
04FE
04DE
04B8
04C9
04E9
04BE
0469
0470
04E9
052D
04CC
0461
04C3
057A
04CF
01C1
FD85
FA84
F9EB
FABD
FB50
FB26
FAEC
FB20
FB71
FB6C
FB24
FAFB
FB05
FB08
FAEF
FAEC
FB25
FB6D
FB87
FB77
FB6C
FB6E
FB54
FB13
FAE2
FAED
FB18
FB28
FB11
FB01
FB1D
FB54
FB83
FBA7
FBC7
FBC1
FB6D
FAED
FAB8
FB08
FB7E
FB93
FB57
FB5C
FBC8
FBE9
FB33
FA7F
FB91
FF0A
033E
05AC
0594
0484
044F
0505
0576
0511
0485
0494
0501
0524
04F9
0508
0567
057E
04F7
045E
045E
04D7
0524
0515
0511
0549
0552
04D0
0428
0405
0477
04E4
04EC
04D0
04D9
04D0
046F
0405
041F
04A8
04EC
049C
0445
0472
04CC
0495
03F2
03EF
04E8
0576
03BF
FFC3
FBBB
F9EB
FA6D
FB7B
FBA2
FB0D
FAB9
FAF3
FB2A
FAF5
FAA4
FAAD
FAEF
FAEC
FA94
FA61
FAA9
FB24
FB59
FB3E
FB29
FB3B
FB3D
FB0A
FADE
FAFB
FB3C
FB45
FB11
FAFA
FB29
FB5A
FB4D
FB2D
FB41
FB72
FB74
FB55
FB70
FBCE
FBE9
FB72
FAEC
FB0F
FBA2
FBAF
FB11
FB31
FD81
0179
04D4
05EB
0551
04C8
051A
0593
0567
04DB
04B3
050A
0550
0534
0505
050E
051F
04EC
0498
0484
04C3
0501
0509
0503
0515
0511
04C0
045A
0451
04B4
050F
050B
04D5
04C4
04D2
04B6
0474
0468
04B7
04FC
04CE
0464
044F
049D
04BF
0471
044C
04E5
0592
04B0
018B
FD85
FAE3
FA7F
FB20
FB28
FA65
F9D8
FA25
FAD4
FB29
FB1F
FB2A
FB5C
FB56
FAF9
FAB0
FAD5
FB31
FB59
FB49
FB57
FB90
FB94
FB33
FACA
FACB
FB16
FB33
FB04
FAEE
FB2D
FB7B
FB7B
FB4C
FB56
FBA7
FBD7
FBAF
FB72
FB63
FB50
FAFF
FABC
FB0A
FBAE
FBB6
FAD4
FA50
FBF1
FFD7
03F6
0610
05E3
050A
04E7
0552
055F
04DA
046E
0494
04FB
051B
04FA
04F6
0515
0502
04A5
045F
0487
04ED
0527
0521
051E
0532
051A
04B5
0451
0455
04AA
04DF
04BD
0480
046C
0474
046F
046F
0499
04C8
04B5
046F
0465
04B4
04D8
0465
03DB
0427
0529
0548
030B
FEFC
FB6B
FA1E
FAAC
FB53
FB17
FA82
FA7A
FAF7
FB4B
FB2F
FB0C
FB3E
FB86
FB81
FB40
FB21
FB37
FB38
FAFE
FAC9
FAD5
FAFF
FB01
FAEA
FB0E
FB7A
FBC9
FBA5
FB3A
FAF3
FAF6
FB12
FB27
FB4A
FB7C
FB89
FB61
FB4E
FB96
FBFF
FC06
FBA4
FB69
FBA1
FBBC
FB1B
FA51
FAFF
FE00
0220
0512
05BA
0514
04C1
0532
059C
055D
04D1
04A6
04E9
051A
04FE
04DF
04FA
051F
0500
04B5
0496
04B1
04C4
04B4
04BA
0506
055B
0555
04F2
049D
04A4
04E2
050B
050A
04F4
04C7
0475
0426
0422
046C
04AE
04AC
04A1
04D4
050E
04D8
0454
0449
050A
058A
042D
00AC
FCB7
FA67
FA32
FACC
FAE3
FA7E
FA69
FAE2
FB4D
FB2B
FAC2
FAA2
FAD7
FAF6
FACE
FAAB
FAD7
FB28
FB4C
FB44
FB48
FB64
FB58
FB10
FAD4
FAF5
FB60
FBB1
FBB0
FB7C
FB48
FB21
FB0D
FB1F
FB52
FB6B
FB40
FB02
FB09
FB50
FB76
FB54
FB4F
FBBB
FC23
FBB3
FA93
FA4E
FC64
006D
0438
05E9
05AA
0510
0528
0591
0584
0508
04CE
051D
0577
055B
04F4
04C4
04EC
0514
04F7
04B8
0499
049B
049B
049F
04CA
050E
052A
04FC
04AF
0487
0491
04AF
04CF
04EC
04F4
04D9
04BF
04DD
0518
0502
0470
03E7
040D
04B8
0500
046D
03CB
0433
055E
0571
02F3
FEA4
FAEF
F98B
FA08
FAC6
FADC
FAA7
FABF
FB02
FAF5
FA97
FA68
FAB1
FB23
FB4D
FB30
FB1B
FB35
FB59
FB5E
FB4A
FB30
FB0A
FAD7
FAB5
FAC1
FAE7
FB02
FB0E
FB1E
FB26
FB07
FAD9
FAEC
FB59
FBB9
FB9E
FB3C
FB37
FBAE
FBD9
FB25
FA5A
FB30
FE57
0260
0506
0570
04CC
04AA
0540
059E
0540
04B7
04C5
054D
058E
0535
04B4
049B
04DE
050A
04EA
04B3
04A4
04BA
04D2
04DE
04E4
04E3
04E4
04FD
0531
054B
0518
04B8
0487
04A9
04D9
04D4
04B5
04BA
04C4
0484
0424
044D
0528
059C
0423
0097
FCBD
FAA5
FAA3
FB49
FB41
FAA8
FA75
FAF2
FB68
FB3C
FAC1
FAAF
FB1B
FB6F
FB48
FAF4
FAF4
FB4A
FB89
FB72
FB36
FB1A
FB2A
FB49
FB66
FB7B
FB73
FB44
FB0A
FAEB
FADE
FAC2
FAA1
FABA
FB16
FB64
FB61
FB47
FB77
FBC0
FB72
FA7C
FA15
FBBF
FF80
0380
05C1
05F8
0575
055F
059D
0581
0503
04C1
04FB
0533
04E7
0455
042B
0492
0503
0506
04C3
04AC
04D3
04E6
04AF
0462
044C
0475
04AA
04C3
04B7
0489
0453
0446
047C
04C3
04CC
0499
048F
04DB
051B
04DC
0467
047D
0525
051D
030E
FF42
FBB3
FA25
FA7B
FB2A
FB1D
FAA1
FA7F
FACD
FAFC
FACD
FAA2
FAD2
FB1B
FB11
FACC
FACD
FB41
FBB8
FBB9
FB56
FB06
FB0B
FB45
FB78
FB92
FB95
FB76
FB40
FB1F
FB30
FB4E
FB4C
FB42
FB68
FBB2
FBC6
FB8E
FB70
FBB5
FBEC
FB64
FA6C
FA91
FD16
0148
04D9
0612
0560
0483
048D
051D
055B
052D
050D
0530
0549
0528
050A
0530
0567
054E
04E8
049F
04B0
04E4
04EE
04D3
04C9
04D7
04CE
04A5
0483
047C
046B
043E
0423
0449
0484
0484
044F
0445
0481
04A0
045A
041B
0473
04FD
0452
0197
FDC6
FAFD
FA64
FB25
FBA0
FB36
FA97
FA81
FADA
FB14
FB04
FAEE
FAED
FACD
FA82
FA66
FABB
FB36
FB53
FAFF
FAAC
FAAF
FAE6
FB05
FB08
FB22
FB51
FB61
FB48
FB40
FB69
FB8F
FB78
FB45
FB3E
FB62
FB74
FB78
FBB8
FC2B
FC2C
FB58
FA8C
FB74
FEBB
02F8
05DE
066B
0594
04E2
04D7
04F6
04DD
04CA
04F3
050E
04C2
044E
044B
04CF
0546
0534
04D2
04B0
04F4
0545
055F
0569
0594
05BD
059F
053F
04E1
04A9
0485
046D
047F
04B5
04CF
04A5
0477
0492
04C3
0494
041C
041B
04E0
055B
03EE
0054
FC4E
FA03
F9F0
FABF
FB11
FAD3
FAB6
FAF0
FB0E
FAD1
FAA4
FAEA
FB5C
FB68
FB0D
FADC
FB2C
FB99
FB95
FB20
FAB9
FAB0
FAD9
FAEF
FAEA
FAE2
FADC
FAD6
FAEF
FB38
FB72
FB4E
FAE7
FABA
FB02
FB62
FB70
FB58
FB86
FBCF
FB80
FA8E
FA4D
FC44
0044
0432
0609
05C3
04F8
04DD
053D
0550
0503
04E7
052F
0567
052F
04D1
04C2
04F4
04EF
0493
0449
0469
04C0
04E9
04D8
04D2
04F8
051E
0525
0526
052E
0516
04CD
049B
04CF
0534
0543
04DC
047D
048D
04C6
04A9
0467
04AE
0560
051E
02AC
FEA6
FB3F
FA1E
FAD1
FBA3
FB9B
FB27
FAFE
FB15
FAF9
FAAE
FAAB
FB0C
FB52
FB1B
FAB1
FAA1
FAF5
FB3A
FB2F
FB17
FB37
FB6E
FB76
FB5B
FB62
FB87
FB7C
FB2A
FAE7
FAF9
FB2F
FB2F
FB03
FAFC
FB20
FB16
FACD
FAC5
FB4E
FBD8
FB90
FACA
FB1C
FDA6
0185
0482
055D
04E1
04A0
0514
0582
0552
04E0
04C7
04F8
04F9
04BA
04B4
051C
0580
0566
04F3
04AB
04B3
04B3
0479
0443
045B
04A3
04CF
04E1
0510
054A
0533
04B8
044E
0461
04C5
0502
04FE
0503
0511
04C4
0415
03D0
049B
05A5
050A
01E5
FDA4
FAC7
FA5A
FB35
FBA7
FB48
FADE
FAE9
FB0A
FAD5
FA90
FAB6
FB29
FB53
FB03
FAB3
FAD1
FB37
FB76
FB79
FB7F
FB95
FB84
FB3C
FB05
FB0B
FB0E
FACD
FA84
FAAD
FB3E
FB9B
FB62
FAF1
FADD
FB1C
FB37
FB1F
FB4E
FBDF
FC1E
FB88
FAF7
FC0D
FF37
02DA
04DB
04D6
043F
0470
053D
059A
0538
04C5
04D9
0534
054A
050D
04D7
04C6
04A0
0458
043F
0482
04DA
04F2
04E5
0504
0541
0539
04DA
049A
04D4
0532
051F
04A4
0467
04BF
0537
053B
04E0
049F
0482
0430
03C2
03F1
04E5
055B
03AC
FFDA
FBFC
FA37
FA9E
FB7E
FB7A
FAD7
FA92
FAEC
FB4D
FB45
FB11
FB04
FB0C
FAF7
FAF4
FB42
FBA9
FBA2
FB1C
FAAB
FACC
FB43
FB7E
FB5E
FB47
FB65
FB69
FB1A
FAD3
FB03
FB84
FBBF
FB83
FB3A
FB37
FB37
FAEC
FAA9
FAFE
FBAC
FBC1
FB07
FAD8
FCCE
00B6
0469
05FA
058E
04CA
04C7
0531
054E
0525
0535
0583
0592
0530
04D0
04D1
04F3
04C1
0455
043A
049A
04FC
04F1
04AE
04A7
04E0
04F9
04D1
04B4
04CC
04D3
0486
042B
0441
04C6
0531
0537
0520
052B
050A
0470
03DB
0422
050B
04EE
026E
FE50
FB01
FA26
FB0A
FBC6
FB73
FABB
FA7E
FAA6
FA9F
FA5F
FA68
FAE7
FB5F
FB5E
FB1B
FB11
FB44
FB58
FB2B
FB0B
FB28
FB45
FB20
FAEF
FB18
FB94
FBE1
FBAD
FB40
FB08
FB10
FB1C
FB1C
FB2C
FB38
FB08
FAC4
FAF5
FBB9
FC43
FBBC
FAB8
FB1B
FE10
0268
058D
0613
04FD
0442
04A9
0564
058F
0545
0526
0552
055C
050C
04AE
0494
04A9
04B2
04B9
04E6
0519
04FD
048D
0436
0454
04B9
04F4
04DD
04AE
04A0
04AA
04B8
04DD
051B
053F
051B
04DF
04D8
04EC
04B6
0440
0438
04FB
0595
045A
00CE
FC91
FA03
F9F8
FB23
FBBB
FB46
FA95
FA63
FA98
FAC2
FACF
FAF5
FB30
FB3B
FB09
FAEA
FB19
FB68
FB85
FB68
FB4E
FB54
FB59
FB43
FB27
FB1C
FB14
FAFF
FAFB
FB2D
FB72
FB7C
FB3A
FAF6
FAE8
FAEF
FAE3
FAF7
FB74
FC0D
FBFF
FB2A
FABD
FC3E
FFCB
03AA
05E4
0610
0559
04EF
04F6
04EF
04BB
04B3
04F9
052C
04FA
049F
0491
04DA
0508
04CB
0456
0412
042C
047B
04C9
04F9
04FD
04E1
04D4
04F8
0527
0507
0490
0437
046E
0503
0553
0518
04B8
04A4
04B7
0486
0432
0454
04E6
04C0
02B3
FF1B
FBD5
FA71
FAB2
FB20
FAD7
FA49
FA4D
FAE6
FB5B
FB40
FAE6
FACF
FB0C
FB4D
FB5F
FB58
FB54
FB4C
FB39
FB2C
FB2E
FB35
FB46
FB7C
FBC9
FBD6
FB68
FACF
FAA6
FB10
FB76
FB4B
FACF
FAC7
FB67
FBFC
FBE2
FB66
FB4D
FBA3
FBAA
FB2E
FB57
FD8E
0192
0546
06AC
05D4
0489
0445
04EE
0582
0575
0519
04EA
04F5
0503
04F9
04E5
04D5
04D3
04F3
0529
0533
04D7
044A
0415
046E
04F2
051D
04F1
04DB
04FD
04F9
0497
0444
0487
0528
0555
04C4
0438
047A
0504
0443
016C
FDA1
FAE4
FA11
FA48
FA4C
F9FC
FA19
FAF0
FBCC
FBD5
FB1D
FA77
FA77
FAE3
FB28
FB0B
FAC9
FAB4
FAE6
FB3E
FB80
FB7A
FB2F
FAED
FB0C
FB82
FBDE
FBCD
FB80
FB64
FB7E
FB66
FAF4
FAA6
FAFB
FBA2
FBB8
FB0A
FABF
FC46
FFAF
035E
0593
05F6
0584
053D
0546
054A
0530
0530
055A
057A
0569
054A
0546
0547
051F
04D5
04A8
04AF
04BF
04B1
049A
04A5
04CA
04DE
04D7
04D4
04D7
04BD
0487
0483
04EB
0569
0559
04A7
0421
048B
0575
054D
02F7
FF19
FBA3
FA04
FA08
FA7F
FAAA
FAB6
FB03
FB68
FB6B
FAFC
FA8F
FA80
FAA6
FAA3
FA74
FA62
FA8E
FAC3
FAD0
FAD5
FB0E
FB6D
FBA5
FB92
FB64
FB4A
FB38
FB1C
FB14
FB3E
FB69
FB48
FAFA
FB01
FB81
FBCF
FB42
FA68
FAE7
FDC6
0200
0549
063F
0598
04FC
0526
057B
053C
0498
044B
049F
0525
0566
0567
0563
0563
0547
0521
052D
0566
057D
053F
04E4
04C6
04E7
0502
04F7
04EB
04F9
04FA
04CD
04A7
04C7
04FD
04DE
047F
048E
0558
05E6
04AA
013E
FD1E
FA62
F9CF
FA70
FAF1
FAF0
FADC
FB06
FB40
FB58
FB67
FB8B
FB92
FB39
FAA3
FA45
FA60
FAB4
FAE2
FAE1
FAF0
FB25
FB4A
FB32
FAF6
FAD7
FAF3
FB36
FB7F
FBA8
FB81
FAFE
FA76
FA7B
FB2E
FBDC
FBA0
FAA1
FA59
FC42
0020
03EF
05C0
057C
04A8
0493
0520
0567
0510
04A6
04AC
04F1
04FA
04C3
04B1
04F1
053A
0544
0524
0511
0505
04E1
04C5
04F7
0566
0596
053F
04B2
0470
048B
04B4
04C6
04F1
053C
054A
04E7
0498
0504
05CF
0578
02E4
FED1
FB60
FA19
FA98
FB55
FB55
FADB
FA9C
FACC
FB1A
FB4A
FB6E
FB90
FB85
FB33
FAD1
FAB0
FAD6
FAFE
FB00
FAFC
FB1E
FB5A
FB85
FB94
FB99
FB8D
FB5A
FB16
FB00
FB2A
FB3D
FAEC
FA78
FA74
FAEB
FB28
FAA6
FA1A
FB06
FE16
0221
0524
061B
05B1
0531
0521
0528
04F1
04AC
04AD
04E3
04FC
04DF
04CA
04E9
051D
0528
0504
04DD
04C3
04A3
047B
0472
04A7
04F8
0528
051F
04F0
04A8
044D
040C
0434
04CD
0558
054D
04D4
04BE
0561
05C1
0460
00FF
FD3A
FB0D
FAE4
FB75
FB6F
FAD9
FA96
FAF7
FB65
FB4D
FAE5
FAB1
FAC2
FAC9
FABF
FAF8
FB84
FBE5
FBAC
FB1E
FADE
FB16
FB56
FB48
FB29
FB4F
FB8F
FB80
FB2A
FAFE
FB29
FB49
FB15
FAEF
FB52
FBE8
FBCB
FAE9
FAA0
FC6F
001B
03A7
054E
0520
0481
0469
04A4
04A9
048E
04C1
0531
054F
04E5
0475
0493
051E
0578
055B
0519
0508
050D
04ED
04C1
04D2
0510
0517
04C5
0484
04B5
0520
0537
04E8
04AD
04CE
04F0
04AD
045E
04AC
0561
0524
02D9
FF17
FBCF
FA6E
FAA7
FB28
FB2A
FAF5
FB0C
FB62
FB8D
FB63
FB20
FAF2
FACB
FA97
FA78
FA8D
FABD
FAD7
FAE0
FB07
FB4D
FB74
FB55
FB20
FB1A
FB39
FB3B
FB15
FB07
FB31
FB4B
FB0F
FABE
FADF
FB6B
FB9F
FB00
FA5E
FB48
FE61
026B
0555
0621
0586
04DF
04D1
051D
055D
0580
0590
0576
0521
04C9
04B8
04EC
0520
052B
0521
0518
04FD
04CC
04B6
04E6
0523
050B
04A8
0484
04F5
058B
058B
04E6
045B
0474
04D2
04C3
045E
047A
0553
05B9
0419
005E
FC5C
FA19
F9F3
FAA6
FAF1
FAC3
FAC3
FB25
FB6F
FB35
FAB1
FA63
FA75
FAB0
FAEB
FB36
FB91
FBBD
FB89
FB23
FAEB
FAFE
FB22
FB2A
FB2D
FB4A
FB61
FB43
FB0F
FB17
FB5C
FB72
FB17
FAB0
FAD0
FB59
FB88
FB1A
FB15
FCDD
0076
0420
05EF
05AE
04D7
04C6
0566
05BD
055F
04D8
04CA
0517
0533
04F7
04C8
04F3
0541
054F
0517
04E1
04DD
04E6
04D3
04A9
0487
0474
046D
0486
04C8
0507
050B
04E2
04D1
04E6
04D3
046B
041F
0484
0544
04FE
0297
FEA9
FB41
F9F1
FA71
FB30
FB1F
FA92
FA66
FAD5
FB57
FB71
FB41
FB21
FB21
FB0F
FAD7
FA9F
FA86
FA81
FA89
FAB1
FAFE
FB44
FB5B
FB5C
FB7A
FBA7
FBA5
FB73
FB6E
FBC5
FC0A
FBBC
FB19
FAFD
FBAF
FC45
FBD1
FAF7
FBA4
FED4
0313
05C7
05E5
04CF
046A
0500
0570
0507
0461
045F
04EA
053F
0519
04F6
053D
05A0
059F
0546
04FC
04E0
04B6
0475
0470
04C7
0515
04EF
048A
046B
049C
0496
0427
03E6
045C
0511
0509
043C
03CF
0475
0509
038F
FFB7
FBA4
F9D3
FA7D
FBAA
FBA5
FAB7
FA43
FACA
FB79
FB7F
FB19
FB01
FB5A
FB9D
FB77
FB2C
FB12
FB11
FAE9
FAAF
FABC
FB22
FB91
FBC1
FBBF
FBAD
FB80
FB35
FB0C
FB3D
FB89
FB78
FB11
FAF5
FB80
FC0E
FBB4
FAB7
FABD
FD1D
012D
04A9
05EB
055D
04A5
04BC
0538
0542
04C1
044A
0443
0479
04A1
04CA
052D
05A9
05CF
056E
04CE
045B
043A
0446
0460
0484
04A3
049F
0485
048E
04CE
0501
04EB
04BC
04D3
051B
050F
0491
0456
04FB
05C6
04F8
01BC
FD6F
FA7B
F9FA
FADF
FB80
FB61
FB2A
FB55
FB91
FB71
FB18
FAE5
FAE2
FAD3
FAC5
FAFE
FB6D
FB8E
FB27
FAB2
FACB
FB4F
FB8F
FB47
FAF3
FB15
FB75
FB87
FB3B
FB0F
FB3C
FB60
FB26
FAF0
FB4A
FBEC
FBD9
FAD4
FA30
FBA7
FF58
0359
0582
0571
048D
044A
04D1
0562
057F
0558
053D
0522
04E1
049F
04A7
04FA
0545
0540
04FA
04A4
045E
0448
0492
0532
05A7
0560
0480
03E3
0427
04ED
054C
04FA
0498
04B6
0503
04CF
0433
0416
04D1
0542
03CD
0042
FC69
FA53
FA63
FB35
FB58
FABA
FA51
FAB2
FB68
FBAE
FB63
FB0F
FB13
FB47
FB53
FB29
FAF9
FAE0
FADA
FAEE
FB2D
FB78
FB89
FB4B
FB12
FB31
FB7F
FB8E
FB50
FB2E
FB5E
FB89
FB57
FB03
FAFB
FB1D
FAE4
FA7D
FB25
FDCD
01A0
048A
055A
04DF
049D
04F7
052D
04D4
0482
04D9
057A
0587
04DB
0446
0476
051F
0577
0536
04C4
0499
04CE
0538
059A
05AC
0542
0495
042A
0449
049F
04AA
0473
048C
0538
05DF
05BE
04FC
0498
0515
0582
0446
00FD
FD30
FAFC
FB01
FBED
FC16
FB3B
FA70
FA8A
FB1C
FB31
FA97
FA13
FA4A
FAF0
FB46
FB12
FACA
FAD3
FB0A
FB22
FB21
FB43
FB79
FB72
FB1C
FAD7
FAF1
FB3B
FB4E
FB1E
FB07
FB2B
FB2E
FAC5
FA74
FB52
FDD5
011D
03A5
04AA
04B0
04A9
04E7
050F
04E0
04AC
04DA
054B
0581
0551
050C
04F4
04E3
04AD
048B
04D3
0554
0574
04FC
0476
0480
04E7
04EE
045F
03EC
043C
04F6
0536
04BF
0459
04BB
057D
054C
033E
FFD6
FCA6
FAFA
FADE
FB52
FB64
FB02
FACC
FB24
FBA3
FB9E
FB0A
FA85
FA86
FADB
FB21
FB50
FB8C
FBAA
FB5D
FAD2
FAA9
FB1A
FB91
FB6C
FAF4
FAF1
FB72
FBA1
FB12
FA9C
FB31
FC4E
FC6B
FB1A
FA09
FB57
FF1F
0336
055E
0551
0475
041D
046E
04D8
04F9
04E3
04CD
04D3
04E6
04EB
04D3
04AD
0497
04AE
04EE
052C
0533
04EF
0490
045F
0478
04AA
04AF
048F
04A4
0514
056F
0522
0459
0410
04CE
05A3
04CE
01AA
FDA0
FAED
FA7C
FB44
FBB0
FB4D
FAD9
FAFE
FB77
FB97
FB39
FADD
FAE9
FB2E
FB43
FB1A
FB04
FB25
FB40
FB18
FAD6
FAC8
FAE1
FAD5
FAAA
FACC
FB64
FBDC
FB8F
FABD
FA6F
FB1C
FBE9
FBAF
FAB0
FAB3
FD18
0128
04A3
05F2
0577
04BF
04CB
0554
0588
051D
0492
0478
04C7
0505
04E9
04A4
0486
048F
0484
0469
0490
0515
0580
054F
04BD
0483
04DD
0536
0518
04E1
0518
0567
0501
0403
03B9
04C8
05B9
043E
0011
FBB2
F9CE
FA77
FB94
FB90
FAC9
FA5F
FA8C
FAA8
FA67
FA42
FAAD
FB68
FBE3
FBF9
FBE1
FBB5
FB68
FB1C
FB16
FB56
FB78
FB31
FAB4
FA87
FAEA
FB81
FBAA
FB33
FAA0
FAA0
FB2F
FB85
FB15
FA97
FBA7
FEFC
032E
05CC
05D9
04B1
044F
050E
05B4
055B
049F
049A
055A
05E2
0590
04DE
048E
049E
047D
040C
03D3
0429
04AE
04CC
0489
0469
049D
04C0
047D
042D
046C
051A
055D
04C1
0408
0443
0530
0511
028D
FE6F
FB08
F9E7
FA78
FB13
FAF0
FA9B
FAC3
FB34
FB4D
FB03
FAE0
FB32
FBA2
FBB5
FB66
FB14
FB06
FB30
FB5F
FB81
FBA0
FBBC
FBC7
FBB9
FB9E
FB82
FB5B
FB23
FAF2
FB08
FB8C
FC22
FC0D
FB29
FAA7
FC2E
FFEF
03EE
05DA
056E
0485
04CE
05EF
0662
05A0
04A8
0471
04B8
04C0
048A
0494
04D4
04B6
0428
03E9
0472
0529
051A
044F
03CA
041C
04A8
049B
041E
0400
0475
04CC
0482
0410
0455
054F
05CE
047F
014D
FD9A
FB1D
FA71
FACA
FAFA
FAA4
FA5B
FAA9
FB37
FB43
FABD
FA70
FAF0
FBBD
FBE1
FB38
FA9D
FACA
FB78
FBD5
FB8C
FB15
FAF9
FB3B
FB91
FBDD
FC24
FC3E
FBF3
FB74
FB48
FB98
FBC8
FB3D
FA6B
FAC9
FD58
0149
0480
0587
04E1
0433
0471
0529
0580
054E
0500
04D5
04A8
047B
0497
0506
0542
04DB
043E
044E
0529
05DF
059B
04AD
0414
0434
0494
04B9
04C1
04E4
04E6
0466
03B1
03B9
04E0
0628
05DD
033B
FF3F
FBE1
FA7D
FAD9
FB91
FB87
FAEC
FAB5
FB3A
FBBB
FB6F
FAAC
FA77
FB21
FBCE
FBAC
FB16
FB0A
FBB1
FC21
FBB7
FAFB
FAC4
FB06
FB16
FAD6
FAD4
FB4D
FBB1
FB80
FB21
FB49
FBCD
FBBE
FAE3
FA7C
FC01
FF5E
02E4
04EB
0529
0482
03FD
0412
04A0
0542
0599
0585
0533
04F3
04EA
04F7
04DE
0491
0434
0403
0427
0495
0503
0523
04F6
04CD
04DA
04FF
050F
0511
0511
04D5
042F
038D
03D3
0526
0628
04F4
0138
FCF8
FAC0
FB23
FC62
FC85
FB66
FA69
FA83
FB27
FB33
FA87
FA26
FAC7
FBCF
FC21
FB92
FB0E
FB40
FBB3
FB93
FAEE
FAA1
FB16
FBAA
FB95
FB0A
FAE4
FB57
FBB7
FB8C
FB43
FB5C
FB7A
FAEF
FA24
FA9A
FD39
0106
0402
0523
050E
04EB
0516
0532
0512
04F4
0507
0524
051E
0504
04F8
04EF
04C5
0476
0435
0437
0475
04AE
04AD
047A
0451
0453
045E
043C
040B
042C
04AE
04F6
047D
03D0
0421
0582
061D
0400
FF97
FBA8
FA7B
FB7F
FC44
FB7A
FA39
FA2E
FB57
FC33
FBCE
FAC9
FA4E
FAA4
FB2C
FB63
FB6A
FB8B
FBAE
FB8E
FB49
FB52
FBCE
FC45
FC29
FB8A
FB02
FB00
FB59
FBA6
FBDC
FC2E
FC71
FC0B
FAE4
FA2F
FB8C
FF26
031F
0544
0537
0485
04A4
0562
058A
04AF
03BD
03BE
0496
0549
053A
04BE
0474
0480
0498
048F
0486
049B
04A3
046D
0421
0428
048E
04CC
046F
03CF
03B6
0441
04A0
043D
03BF
043E
0561
0524
021C
FD9E
FAAC
FAA9
FBED
FC1A
FAF8
FA3E
FAEF
FC0D
FC34
FB7B
FB0D
FB53
FB88
FB26
FACA
FB2D
FBE6
FBF8
FB57
FB06
FB99
FC5F
FC58
FB90
FB0C
FB68
FC16
FC33
FBB8
FB70
FBC3
FC14
FB99
FAA7
FAC8
FD33
013F
04A3
0598
049D
03C5
044B
0562
0588
0490
03C0
0413
050D
0581
0515
0472
042F
0433
0441
0472
04D2
04E8
0446
035F
0331
0405
04FC
0523
04A0
045D
04A9
04D1
0446
03A3
03F3
0510
055A
036A
FFC5
FC76
FB0D
FB3E
FB99
FB44
FAAE
FAA0
FB18
FB65
FB28
FAC6
FAC8
FB2B
FB7F
FB89
FB7D
FB91
FBB1
FBB7
FBB4
FBD3
FC00
FBF3
FB96
FB3F
FB49
FBA1
FBDC
FBC2
FB8D
FB98
FBE0
FBF3
FB85
FB11
FBC4
FE59
020A
04F3
05C9
0513
047D
04EC
05AF
05A7
04D8
0450
04A8
054E
056E
050E
04C7
04CB
04BF
0475
043C
044F
0469
0437
03EF
040C
0480
04AE
044B
03DA
03EB
044F
0472
044C
0472
051C
058A
049A
01F5
FE88
FBCD
FAAA
FADA
FB54
FB3F
FAA8
FA57
FAC8
FB7F
FB8C
FACE
FA35
FA94
FB90
FC18
FBBD
FB17
FAE0
FB20
FB70
FBA7
FBE3
FC03
FBB7
FB28
FB09
FBAA
FC67
FC66
FBBD
FB43
FB58
FB68
FB06
FAF3
FC7F
FFD4
036A
0576
05A4
050C
04BC
04C8
04C6
04AE
04D9
054F
0595
0549
04A8
044C
047A
04E2
050C
04D7
0475
0422
03FF
041D
0476
04D4
04EA
04A1
043A
0408
0418
0439
0448
0458
0489
04BA
047F
0360
013C
FE88
FC2C
FAF9
FB03
FB83
FB94
FB14
FAA3
FAB8
FB0A
FB05
FAA1
FA64
FAAD
FB3F
FBAA
FBD4
FBE2
FBD8
FBA1
FB6A
FB85
FBD5
FBC6
FB21
FA8D
FAD3
FBD0
FC8C
FC5C
FB8F
FADA
FA85
FA7F
FAF8
FC5E
FE9F
0100
02DE
043B
0546
05C1
055D
0473
03E7
042F
04E9
0572
059A
0583
0527
047B
03E3
03F6
049D
04FC
048E
03E3
03DB
046D
04CA
0491
044D
0484
04EB
04E2
0482
0487
0532
05D8
05C4
050D
041D
02CA
0096
FDB8
FB4B
FA3E
FA6A
FAF4
FB47
FB63
FB5F
FB23
FAC6
FAB2
FB22
FBAA
FBAE
FB35
FAE1
FB1E
FBA4
FBED
FBD6
FBA7
FB94
FB88
FB6D
FB59
FB61
FB6A
FB55
FB2A
FAF4
FAA2
FA68
FB13
FD75
0140
04BF
0630
0572
0412
03A3
044F
0522
0560
0518
04B1
0464
044E
0494
0522
0575
0520
0476
0440
04B6
052B
04FD
0475
0450
04A1
04C0
0455
03EE
0436
04FA
055C
04EF
03FB
02B3
00C9
FE26
FBA1
FA5A
FA8E
FB68
FBFB
FBFF
FBA1
FB15
FAA1
FAB1
FB66
FC1B
FBF3
FAF1
FA1E
FA42
FAF5
FB4C
FB07
FAA9
FAA1
FADC
FB35
FBBA
FC45
FC4C
FB88
FA96
FA62
FAF9
FBA4
FC46
FDD9
00FB
0479
063D
059D
0417
0386
042C
04E2
04CF
043F
03E4
03F1
043D
04BB
054B
057E
0511
0486
04AD
0586
061F
05C3
04EB
0497
04F5
0539
04DC
045A
0475
0519
0587
054C
0482
0325
00D2
FD91
FA7D
F912
F9B5
FB53
FC75
FC78
FBA9
FAB2
FA37
FAAB
FBE6
FCF0
FCB8
FB50
FA16
FA47
FB89
FC57
FBC5
FA72
F998
F9AE
FA48
FAE9
FB5A
FB6D
FAF5
FA40
FA0A
FAB5
FBC8
FCB6
FDD7
0008
0326
05AE
0643
0543
0442
0442
04E1
054C
0543
0505
04B6
0458
042B
0473
04E5
04D5
043A
03E1
045B
0521
055A
0513
0512
058C
05C2
053A
04A0
04EF
05F4
0671
05B3
0445
02C1
00CC
FDEB
FAEA
F96B
FA07
FB8D
FC5A
FBFD
FB25
FA77
FA18
FA32
FAFF
FC16
FC5B
FB56
FA20
FA46
FBD4
FD28
FCE1
FB6C
FA54
FA71
FB41
FBDB
FBE0
FB60
FA7D
F987
F923
F9BF
FB0E
FC7E
FE1A
006C
036B
05F5
06CB
05E3
0467
0388
03A0
046F
057D
0624
05BD
046F
036B
03CD
0533
060A
0566
0413
037C
03EF
048D
04B7
04B4
04CF
049F
03E1
0361
042D
05F6
071B
067E
04B2
02E0
0115
FE89
FB6F
F95F
F983
FB07
FC16
FBEE
FB4D
FB00
FAF1
FAD4
FAF2
FB9A
FC3B
FBEA
FACD
FA36
FB01
FC56
FCBA
FBE2
FAE1
FAB4
FB3F
FBD3
FC16
FC0D
FBA7
FAD5
FA01
F9E5
FACD
FC55
FE1E
003A
02AA
04C8
05C5
058E
04CF
0428
03CD
03E9
04BA
05E2
063D
050D
034A
02E4
046C
062B
0626
0480
032C
0371
049E
054F
0524
04B5
0459
03EC
03A8
043A
059A
0686
05DA
03F3
020C
007F
FE8E
FBFB
FA00
F9F3
FB74
FCB4
FC8D
FB8E
FAD6
FAA4
FA9D
FACD
FB81
FC51
FC3E
FB0C
F9D9
F9E8
FB0F
FBFA
FBD1
FB10
FAA5
FAD4
FB4F
FBD8
FC46
FC33
FB50
FA15
F99A
FA93
FCAD
FF24
0187
03AA
052B
05A2
054F
04FB
04F1
04B1
0401
03A8
046D
05A6
05BE
0457
0311
039A
0570
0672
0593
041A
03CA
04B5
057F
0554
04AD
0441
041D
0411
045C
0534
0603
05C1
0432
0214
0008
FDE2
FB84
F9C3
F99C
FAC8
FBD4
FBC6
FB10
FAB1
FADD
FB20
FB64
FC00
FCBF
FCAF
FB6D
FA11
FA0D
FB5B
FC80
FC53
FB36
FA61
FA6F
FB0E
FBB6
FC15
FBE6
FB0D
FA13
FA04
FB58
FD6A
FF5C
0124
0332
0542
0659
0610
0540
04EB
04F3
0493
03E1
03E1
04D7
057C
04A0
0306
029E
0402
0597
0596
0437
0333
0387
0484
0516
0516
04F9
04D8
0482
043B
0495
0577
05E1
04E4
028C
FF99
FCC3
FA87
F970
F9CB
FAFC
FBC6
FB93
FB0B
FB12
FB8F
FBC0
FB8A
FB9E
FC43
FCA9
FBFF
FAD2
FA96
FBC7
FD2C
FD4A
FC18
FAD8
FA96
FB4D
FC49
FCCE
FC5D
FAFD
F985
F941
FABE
FD2B
FF4F
00FA
02F1
054F
06DF
068C
04F9
03DC
03F9
0484
0496
046D
04B2
0513
049A
0354
02AC
0395
0516
0569
043F
0316
0344
046B
052B
04DE
0411
0387
0378
03D1
0495
0588
05E8
04F9
02C5
0003
FD68
FB62
FA4F
FA62
FB2E
FBBA
FB73
FAE5
FAF9
FBAE
FC17
FBB8
FB4E
FBB5
FC8B
FC9E
FB97
FA8E
FAB3
FBD7
FCB5
FC71
FB6B
FAA2
FAB9
FBA3
FCC8
FD42
FC6E
FABF
F9B5
FA84
FCDA
FF52
011D
02A8
0471
05D4
05C7
047D
037C
03D1
04DB
0560
0535
051C
054A
050C
0412
0351
03DA
0537
05C3
04C2
035C
032B
044A
056A
0578
04A5
03CB
0387
03F7
04E9
05CE
05D1
0472
021E
FFC7
FDE2
FC35
FAB3
F9F9
FA75
FB82
FBF2
FB76
FAD8
FACF
FB0F
FAED
FA8C
FAB2
FB80
FC0E
FB9A
FAA6
FA5F
FB25
FC2A
FC6E
FBC5
FACD
FA4C
FAA6
FBA5
FC77
FC27
FAA6
F947
F9B3
FC3A
FF7F
0206
039D
04E0
05E1
0605
053B
0474
0487
0512
051F
04A3
0493
0552
05E9
0557
0426
03DA
04EB
0617
05F6
04B7
03C5
040C
050A
05AB
0570
04AA
03FE
0405
04FD
065C
06DA
057A
0293
FF8A
FD5F
FBE5
FA90
F990
F98F
FA80
FB53
FB33
FA8E
FA69
FB00
FB97
FB97
FB48
FB3A
FB64
FB44
FABA
FA4C
FA7C
FB1A
FB78
FB29
FA5F
F9C5
F9FB
FB0C
FC23
FC1A
FAAE
F922
F945
FBA8
FF13
01DC
0387
04AE
05AE
0614
0595
04DA
04C4
053C
0560
04E0
047D
04E3
058E
056D
0471
03C9
045C
0599
062C
0596
04A6
0464
0507
05F5
066D
060A
04F9
0402
0418
055D
0696
0616
0367
FFD7
FD18
FBA7
FAE4
FA5D
FA5E
FB10
FBC4
FB9B
FAB5
FA1E
FA75
FB25
FB3D
FABA
FA76
FAEE
FB9D
FBAE
FB04
FA55
FA48
FAC5
FB22
FAE5
FA43
F9F0
FA68
FB4F
FBA9
FADD
F9A5
F998
FB9C
FEEB
01E3
03A6
0497
0555
05C6
057A
04AC
043E
049A
052F
0543
04F4
04EC
0552
058C
052E
04A3
04A8
0541
05B4
0578
04D9
048C
04DE
0585
05FE
05E4
0536
0476
0472
0567
0660
05D2
032D
FF9C
FCE3
FB9F
FB10
FA7B
FA26
FA98
FB6E
FB9C
FAE0
FA34
FA8B
FB7E
FBCD
FB01
FA0A
FA07
FAE5
FB90
FB4F
FA88
FA26
FA86
FB2E
FB67
FB04
FA8F
FAB7
FB81
FC1B
FBA3
FA4E
F98D
FAD1
FE08
01A4
0421
0543
05B8
05E8
05AA
04FD
0473
0492
051E
0564
052A
04EE
0518
056A
056A
051D
04F9
0538
0589
0582
0518
0495
044B
0464
04C7
0513
04D8
0434
03F7
04CA
05FF
05DF
0372
FFC6
FCDE
FB93
FB09
FA47
F9A4
FA10
FB60
FC2A
FB87
FA4E
F9F9
FAC8
FB8F
FB55
FA7D
FA18
FA82
FB1B
FB37
FAE7
FAB2
FADF
FB3E
FB80
FB88
FB76
FB8B
FBDB
FC13
FBB8
FADC
FA76
FBA2
FE74
01BE
0423
0544
05A1
05A2
053D
0489
0423
048A
055B
05B9
0556
04C8
04B6
050D
0544
0519
04D1
04BC
04DA
0502
0514
04F6
04A2
0464
04A6
053E
0553
046C
0368
03B1
0539
05E6
03B8
FF4F
FB87
FA61
FB0E
FB6B
FACB
FA58
FAF5
FBD6
FBB5
FAB3
FA2E
FAD0
FBB0
FBA5
FADA
FA70
FAE2
FB83
FB8D
FB26
FAF7
FB34
FB71
FB55
FB11
FAFB
FB07
FAF3
FAD4
FB3F
FCCC
FF80
02A2
051C
0625
05D6
0519
04D8
0536
0596
056B
04D5
0469
0475
04BA
04D6
04C0
04B0
04C6
04E2
04D1
0485
042F
0431
04BF
0578
058E
04B8
03D3
0423
0598
0646
043F
FFF3
FC10
FABC
FB65
FBD1
FAFD
FA0F
FA5E
FB7E
FBDF
FB09
FA33
FA88
FB8D
FBEC
FB4D
FAAD
FAE3
FB8D
FBC3
FB57
FAEB
FAE8
FB09
FAF6
FAEC
FB51
FBE2
FBD6
FAFA
FA4E
FB47
FE5A
0258
054D
0612
052F
0432
043B
0512
05A6
0558
049A
044B
04A6
0516
050A
04A2
0465
0488
04CB
04E3
04CC
04B6
04CA
050B
054B
0532
0494
03EB
041E
055A
0641
04EC
011A
FCE1
FAB4
FAE0
FB99
FB5D
FA9E
FAA5
FB7B
FBDB
FB28
FA63
FAC0
FBDA
FC35
FB4F
FA55
FA84
FB8D
FC19
FB97
FAD0
FAA8
FAFA
FB19
FAF0
FB03
FB6D
FB8E
FB03
FA91
FB96
FE8E
0250
04FD
059B
04D1
0416
044E
051B
057F
050A
0458
0452
050B
05A3
055B
047E
0401
0457
04FA
0523
04B3
0437
0432
04A1
0522
0554
0510
0497
047D
0516
05B4
04E5
01EA
FDDF
FAEE
FA38
FADC
FB47
FB0B
FAE6
FB3B
FB63
FAD7
FA3A
FA8E
FB9F
FC1B
FB5B
FA5C
FA75
FB85
FC25
FB9F
FAD7
FAF8
FBCE
FC28
FB8A
FACC
FACB
FB3B
FB42
FAEF
FB7C
FDD9
0163
045D
0594
054D
04AF
0493
04F3
054B
0547
0513
0506
052F
053A
04E9
0476
045E
04C6
053A
0522
047F
03EF
0408
04B3
0551
0553
04AD
03E7
03BA
0469
053D
04CA
0238
FE54
FB2B
FA30
FAEC
FBBC
FBA5
FB17
FAD9
FAEC
FAD3
FA96
FAB7
FB40
FB7D
FB03
FA77
FAC6
FBBB
FC22
FB6E
FA97
FACB
FBC6
FC2E
FB80
FAC4
FB0C
FBDE
FBDE
FAF4
FAD5
FD16
0121
04AA
0608
0593
04C8
0499
04DF
0513
050A
04E9
04CF
04BD
04BA
04CE
04ED
04FD
04FE
04F6
04DD
04A7
047A
0496
04FD
0544
04FA
0437
03B7
0427
0556
061C
052D
0242
FE7A
FB97
FA92
FAE8
FB51
FB20
FABB
FACC
FB40
FB74
FB27
FAD6
FAFC
FB59
FB5C
FB08
FAF7
FB5B
FBA0
FB46
FABC
FACC
FB66
FB9B
FAF8
FA57
FAB9
FBB9
FBEF
FB05
FAA7
FCB4
00D5
049A
05FA
053F
043A
041E
04A4
0502
0505
04F9
04F8
04DA
04A9
04B0
0502
0546
0528
04C3
0479
0476
0496
04B3
04D2
04F8
04FE
04C6
048F
04C5
0572
05E6
0523
02B3
FF3F
FC35
FABA
FABE
FB39
FB49
FAFD
FAF1
FB51
FB93
FB4C
FAD9
FAEA
FB77
FBBF
FB5F
FAE2
FAF5
FB63
FB6E
FAF7
FAB6
FB16
FB83
FB46
FABB
FADA
FB9A
FBC0
FAC6
FA34
FC24
007A
048D
05E8
04E0
03C7
040A
04F1
0531
04C4
0491
04E1
050E
04B6
045F
049C
051F
0524
04A0
0458
04BD
0547
053B
04B5
0470
04B4
04FC
04DB
04AF
050D
05AB
0551
0319
FF8B
FC47
FA9C
FA85
FB0A
FB53
FB43
FB30
FB45
FB5A
FB45
FB2A
FB3F
FB72
FB77
FB3D
FB0D
FB1D
FB3D
FB1E
FADD
FAEC
FB61
FBAF
FB5F
FAD1
FACB
FB4D
FB6C
FABF
FA72
FC3B
002D
042B
05F4
0567
045A
044F
0501
054B
04DE
0477
049D
04ED
04D6
047A
0470
04D2
051B
04EC
0498
0499
04D9
04E1
049E
0486
04D6
051B
04D4
0450
046C
0543
058A
03BE
FFF1
FC15
FA38
FA96
FBAA
FBF5
FB63
FADB
FAEB
FB3C
FB45
FB0E
FAF8
FB0F
FB06
FACB
FAB9
FB0A
FB6D
FB72
FB2E
FB20
FB62
FB7E
FB29
FAE0
FB3C
FBE8
FBD7
FAD6
FA52
FC05
FFD6
03AE
0585
054F
0499
0490
04F7
0507
04AF
048A
04DE
0540
053C
04FB
04ED
051B
0524
04DB
0498
04BB
051B
0538
04F0
04A6
04AF
04D7
04B4
0463
047B
0522
0564
03EA
007C
FC9E
FA51
FA3E
FB40
FBC3
FB54
FAB3
FAA1
FAFF
FB3A
FB1C
FAF7
FB06
FB1D
FB0C
FAF4
FB07
FB29
FB15
FADE
FAE4
FB3E
FB7E
FB4E
FB07
FB46
FBDE
FBDE
FAE4
FA21
FB67
FF10
0349
05BC
05C8
04CB
0468
04E8
0575
056F
0518
04EB
04EC
04CB
0488
047E
04D3
0533
0538
04F3
04CD
04EA
04FC
04C5
0483
0495
04D9
04CE
045D
0432
04D4
0587
04A9
0174
FD3C
FA63
FA0F
FB28
FBCB
FB4F
FA94
FA8E
FB14
FB5F
FB2F
FAFC
FB17
FB39
FB0C
FAC5
FAD5
FB2F
FB59
FB2B
FB10
FB58
FBA7
FB7A
FB01
FAF7
FB7E
FBC3
FB26
FA7E
FB83
FECA
02C9
0547
058B
04CA
0486
04F3
0542
0501
04A3
04B8
0513
0525
04CD
0483
04A2
04F0
04FE
04C8
04AF
04D9
04FC
04D8
04A3
04B8
04F6
04E0
0467
0439
04DD
059A
04CD
01AA
FD6F
FA79
FA00
FB17
FBE4
FB99
FAE2
FAA8
FAEE
FB25
FB14
FB0F
FB42
FB5E
FB22
FADD
FB04
FB7B
FBAA
FB57
FB00
FB25
FB8E
FBA6
FB64
FB55
FBA9
FBBB
FB07
FA52
FB3C
FE62
025F
0507
0582
04D9
0481
04D0
051D
04F9
04B8
04CB
0510
0514
04CC
04A6
04E0
052F
0526
04CC
0489
048E
04A4
0498
048C
04B7
04E9
04BC
043C
0410
04A8
0553
0497
01C2
FDEA
FB1C
FA72
FB26
FBA2
FB40
FAA8
FAB1
FB40
FB95
FB5D
FB06
FB03
FB30
FB22
FADE
FAD3
FB29
FB7B
FB6D
FB2F
FB2D
FB60
FB5D
FB18
FB11
FB8B
FBE9
FB73
FAA1
FB18
FDE6
0205
0522
05E2
050F
0460
0493
050B
0514
04D6
04D9
051B
051C
04B3
045D
048D
04FF
051C
04CC
048D
04B1
04ED
04D6
048E
0489
04C6
04C7
045E
0431
04DC
05BB
051E
0219
FDDE
FAD0
FA39
FB32
FBE1
FB7F
FAC4
FA9E
FB02
FB48
FB32
FB20
FB54
FB7F
FB42
FAD3
FABD
FB1A
FB6C
FB56
FB1B
FB2C
FB71
FB6F
FB13
FAEB
FB53
FBC1
FB70
FAAB
FAF6
FD72
015C
0491
059D
050B
0479
04C1
0554
055C
04DB
0481
04A6
04F0
04F2
04C7
04C6
04F3
04FD
04D1
04C0
04FB
0537
0515
04BF
04B7
0508
051E
049F
0423
0483
056E
0549
02D2
FEC6
FB64
FA3D
FAD6
FB8D
FB76
FAFC
FAD9
FB11
FB2C
FB08
FAF9
FB2E
FB58
FB22
FAC1
FAB0
FB09
FB63
FB63
FB2A
FB0E
FB17
FB09
FADE
FAEA
FB58
FBB6
FB6B
FAB4
FAD6
FCF6
00B1
042B
05B3
0549
0468
0454
04F0
054E
0512
04C8
04F2
0545
052E
04B8
0485
04D8
0530
050B
04AA
04AB
050A
0521
04B2
0458
049F
0522
051F
04B6
04CB
0579
0557
02FA
FEFA
FBA7
FAA0
FB3A
FBAF
FB42
FAB0
FAB9
FB1B
FB2C
FADE
FAB6
FAEF
FB38
FB45
FB33
FB2F
FB28
FB0B
FB05
FB2F
FB4A
FB20
FAFA
FB36
FB8B
FB42
FA76
FA93
FCEB
00EC
045E
059D
051E
047A
0483
04DC
04FD
04F7
0503
0503
04CF
049F
04C3
0517
052B
04FD
04FA
0533
052D
04B5
0460
04AF
052C
0505
0472
048C
057F
059A
0318
FE99
FAE5
F9F9
FB0A
FBE7
FB9A
FAF0
FAD7
FB2D
FB56
FB3F
FB36
FB41
FB23
FAED
FAFB
FB3F
FB38
FACA
FA8F
FAF0
FB71
FB64
FAF6
FAD9
FB0D
FADE
FA51
FAD2
FDA2
01DE
0508
05B2
04E1
046E
04C9
050C
04B6
0459
047F
04D7
04D3
0496
04A9
0507
0527
04ED
04E2
0540
0578
0515
048D
0492
04FA
050B
04C5
04E9
057C
050E
024F
FE18
FAE5
FA2A
FAEB
FB50
FAE7
FA98
FAEA
FB5A
FB57
FB1F
FB34
FB7B
FB81
FB42
FB28
FB42
FB25
FAB7
FA7A
FAC1
FB18
FB05
FAD3
FB0F
FB69
FB11
FA4E
FAD6
FDE1
0242
0554
05CB
04E4
0481
04FA
0560
053A
050A
0532
0545
04D4
043B
042B
049E
04EA
04C7
04A1
04CC
04FE
04E3
04B7
04CD
04F0
04CD
04BB
0546
05EA
0509
01C9
FD88
FABD
FA63
FB2F
FB71
FAFB
FAB1
FAEB
FB1D
FAED
FABE
FAF6
FB4B
FB43
FAFF
FB01
FB50
FB69
FB21
FAF5
FB38
FB86
FB66
FB16
FB1A
FB42
FAF0
FA6B
FB20
FE07
0219
0512
05BE
0502
047A
04A8
04F7
04F2
04CA
04CA
04E6
04F5
0506
0525
052A
04FB
04CF
04E5
050F
04EB
0496
0495
04F7
051B
04B0
046A
04FE
05AE
04AB
0145
FD1C
FA98
FA6A
FB34
FB78
FB2E
FB18
FB5E
FB7D
FB45
FB1D
FB39
FB3F
FAE9
FA91
FAB2
FB25
FB4F
FB0B
FAD5
FAFF
FB40
FB47
FB40
FB58
FB33
FA8A
FA26
FB85
FF0C
0322
0595
05C7
04FA
0499
04C4
04D2
048F
0469
049D
04E7
04F6
04D7
04BC
04B7
04CE
0511
0564
0568
04F2
047B
0496
050C
0510
0482
045B
0534
05E3
0475
0097
FC62
FA3D
FA73
FB57
FB7F
FB17
FAF1
FB22
FB2F
FB01
FB00
FB4E
FB8E
FB7B
FB4A
FB2E
FB05
FAB3
FA95
FB00
FB91
FB83
FADD
FA8A
FAFF
FB70
FB12
FAAF
FC0B
FF9A
038B
059C
057B
04BC
04AF
0519
0528
04D1
04AB
04DE
04FE
04D4
04AF
04D0
04F9
04DD
049A
0480
0498
04B6
04E2
0539
0568
04F5
0432
0434
0544
05E0
041C
000F
FC13
FA5B
FABE
FB62
FB2A
FAAB
FAC6
FB49
FB67
FB07
FACF
FB13
FB6D
FB6E
FB31
FB0D
FB0F
FB16
FB21
FB3D
FB40
FB0F
FAFE
FB6F
FBF3
FB92
FA55
F9F3
FC20
0059
041B
0583
0518
04AB
0508
0571
0531
04B4
04AF
04FC
04F8
049A
047A
04D1
0524
0509
04C3
04C5
04FC
0506
04D9
04BC
04A9
0459
0406
046F
0589
05D6
03C2
FFAD
FBDD
FA36
FA7D
FB1E
FB25
FAE4
FAE7
FB17
FB24
FB28
FB53
FB70
FB33
FAD8
FAD7
FB2B
FB53
FB26
FB12
FB5A
FB87
FB29
FABA
FB0C
FBD8
FBD9
FACA
FA6B
FCAD
0113
04DF
0606
052C
0468
04AA
0528
050A
04A3
04AC
0511
0533
04EE
04B4
04BE
04CB
04AB
049A
04C7
04F9
04EC
04C8
04D4
04E1
0494
043B
0491
0564
0522
0282
FE5B
FB15
FA2B
FADD
FB76
FB4B
FAF5
FAFB
FB17
FAEC
FAC3
FB04
FB7E
FBAA
FB70
FB2B
FB0D
FAF8
FAE8
FB10
FB66
FB82
FB3F
FB29
FBAF
FC30
FBAB
FA7E
FAA3
FD7A
01D6
0508
05B6
04FC
04A1
0509
055B
0524
04E0
04F3
04FA
048E
041A
0447
04F1
055A
0534
04F1
04F1
0504
04E6
04BD
04C1
04AD
0434
03D0
0450
054E
0502
0231
FDFD
FAEA
FA3A
FAE4
FB40
FAED
FAB4
FAFC
FB49
FB31
FB05
FB30
FB79
FB6D
FB1F
FAFF
FB1B
FB17
FADF
FACC
FB11
FB5B
FB6A
FB82
FBE3
FC10
FB69
FA8B
FB35
FE48
025C
051A
05AD
053F
0520
054F
051F
049F
0487
04FC
0544
04E5
0460
0466
04D4
050F
04FF
0509
0538
0521
04AD
0461
0487
049F
0431
03D3
046F
0577
04DF
0189
FD0C
FA3D
FA21
FB2C
FB7D
FAEC
FA91
FADE
FB30
FB05
FAC4
FAED
FB44
FB43
FAF4
FACA
FAE3
FAFD
FB10
FB56
FBBB
FBCD
FB75
FB49
FBA8
FBE9
FB47
FA79
FB74
FF01
0354
05C7
05AC
04A9
046C
04EF
0534
04FB
04E3
0537
0572
0537
04EA
0502
053E
0522
04CE
04BF
04E8
04C6
0448
040C
0467
04CB
04A4
0466
04D7
056F
046A
0103
FCE5
FA8D
FA95
FB61
FB5A
FAA7
FA5B
FABF
FB20
FB0C
FAD8
FAE6
FB05
FAF0
FAE2
FB20
FB62
FB40
FAEF
FB00
FB72
FBA4
FB57
FB1C
FB5F
FB8B
FAF1
FA54
FB8B
FF2A
0358
05A6
05A7
04F3
04E7
0546
053B
04CF
04B1
0500
0526
04DF
04AA
04E4
0526
04FA
04A8
04C4
052D
0538
04C3
046A
048C
04BA
0491
0489
052B
05A4
0439
007B
FC5A
FA38
FA70
FB5F
FB98
FB41
FB22
FB4D
FB3F
FAE6
FABD
FAFB
FB43
FB4F
FB56
FB7B
FB67
FAE8
FA84
FAD0
FB76
FB9B
FB2A
FAF8
FB6B
FBAD
FB05
FA79
FBFF
FFDE
03D4
0585
0508
0453
0492
0516
04EC
0460
0463
0501
0559
0501
048D
0497
04E0
04E5
04BC
04C8
04F2
04DB
0499
049E
04E9
04E7
047E
046C
051D
0572
03B7
FFE7
FC24
FA75
FAB2
FB3A
FB2E
FB0F
FB5D
FBAA
FB69
FAEF
FAF2
FB5D
FB70
FAFB
FAB8
FB1C
FB9C
FB8C
FB36
FB4C
FBB7
FBBA
FB36
FAEE
FB3D
FB5F
FAB4
FA4B
FC02
0009
0422
0600
05A8
04E2
04CD
04FF
04CF
0476
0485
04DF
04F7
04C5
04C3
0500
04F5
0479
0430
0491
0519
0507
0481
044D
048B
049B
0455
0480
056A
05BA
03A6
FF6E
FB8F
FA19
FA90
FB16
FAEC
FADA
FB69
FBE6
FB8B
FAC7
FA9D
FB27
FB88
FB4E
FB0A
FB40
FB8B
FB5B
FAF4
FAFD
FB66
FB8C
FB54
FB53
FBAB
FB94
FAB4
FA5C
FC62
009C
048F
0607
0562
04A0
04C8
0529
04FF
04A1
04BD
0522
0516
0490
0453
04B5
0518
04EB
0485
0488
04E0
04F8
04B5
048D
04AD
04B9
049A
04C8
0554
0514
02B7
FEBA
FB6A
FA7C
FB3B
FBB4
FB22
FA79
FAA7
FB4C
FB81
FB32
FB0D
FB52
FB85
FB4F
FB0E
FB2B
FB65
FB46
FAE4
FABF
FAF3
FB2D
FB49
FB7D
FBB9
FB7C
FAD1
FAF1
FD36
0134
04AF
05D8
0521
0466
049D
0521
0512
04A3
0492
04F4
0525
04D2
046D
047B
04D3
04FA
04DD
04CE
04EE
0509
04F8
04CE
04A5
0487
049E
0517
0585
04C3
0207
FE1F
FB1E
FA5B
FB2A
FBD3
FB8C
FB00
FAFF
FB59
FB55
FADC
FA94
FAE0
FB55
FB60
FB13
FAF2
FB22
FB3E
FB0B
FADF
FB28
FBB6
FBD4
FB38
FA9C
FB4A
FDE2
0190
0496
05B1
051D
0442
0445
0500
0571
0515
047C
0472
04F6
0555
052D
04DF
04E6
0519
04FF
049D
047D
04C7
04F3
0498
0435
0488
0531
04AE
0201
FE22
FB38
FA70
FB03
FB6A
FB23
FADA
FB21
FB9B
FB96
FB0F
FAA8
FAC1
FB08
FAF9
FAA5
FA8F
FAED
FB5C
FB6F
FB46
FB5A
FBAD
FBA8
FAF1
FA4B
FB2C
FE36
0235
050C
05A3
04D5
044A
04B0
0553
055A
04DD
0499
04CF
0501
04CF
0492
04D1
0563
0593
051D
0498
04A0
04F9
04EA
0467
044A
051B
05E7
04F3
01A8
FD7C
FAB0
FA3A
FB1B
FBB1
FB5E
FAC3
FAA9
FB0E
FB5A
FB3C
FAF2
FAD9
FAEE
FAEF
FACD
FAC8
FB04
FB44
FB39
FB04
FB0F
FB68
FB7C
FAE6
FA4E
FB27
FE28
0238
0537
05F7
0536
0494
04CF
0551
054C
04D1
048F
04D6
0538
0539
04ED
04BF
04CD
04DC
04D0
04E1
0527
054A
04EB
0451
0442
04FD
0588
0473
0160
FD9E
FB0C
FA6D
FAF0
FB48
FAFC
FA90
FA98
FAF9
FB33
FB14
FAEC
FB04
FB35
FB2B
FAEE
FADE
FB23
FB67
FB4D
FB05
FB12
FB74
FB82
FAD6
FA46
FB60
FEB2
02D1
057D
05C0
04B6
0422
049C
0556
0572
050D
04D3
0501
0532
051B
04F3
0506
052C
050A
04AF
0496
04E7
0520
04BE
0416
0413
04F1
0594
0479
0159
FD9C
FB18
FA6D
FACB
FB10
FAEA
FAC8
FB00
FB53
FB55
FB05
FAC7
FAD7
FAFE
FAEA
FAB1
FABB
FB25
FB86
FB6F
FB0F
FB00
FB68
FBAA
FB3D
FABC
FB9C
FE92
027B
0541
05DC
052A
04B4
04FB
0552
051D
04AC
04A3
0503
0537
0501
04D4
051B
0588
057A
04F2
049E
04E5
0546
050C
0462
043C
04FD
0597
046F
0123
FD28
FA7D
F9E3
FA7C
FAF6
FAE0
FAB5
FAF1
FB61
FB79
FB19
FAB2
FAB1
FAFB
FB23
FAFD
FACC
FAD3
FAF2
FAEC
FAD7
FB08
FB71
FB7F
FAEB
FA82
FBAD
FEE7
02E6
059A
061F
0562
04E5
0527
0580
054B
04C3
0491
04E0
053E
054E
0534
053A
054C
0522
04C9
04AD
04FB
0548
0513
0488
046A
04FC
0550
0401
00C0
FCEE
FA74
FA06
FAB1
FB1B
FAE1
FA98
FAC4
FB22
FB34
FAFC
FAEE
FB24
FB27
FAA5
FA11
FA29
FAF5
FBA4
FB90
FB13
FAF7
FB53
FB68
FADE
FAB3
FC56
FFE6
03AF
05BA
05AC
04D8
04A7
0535
05A7
0575
04F6
04BD
04DC
04FB
04FA
0512
0560
0593
054F
04C3
0489
04DC
053B
050E
0483
0465
04F0
051C
037C
FFF5
FC2E
FA1F
FA32
FB17
FB60
FAEF
FA9F
FAEB
FB5C
FB53
FAE7
FAB3
FAED
FB26
FB01
FABC
FACA
FB1D
FB37
FAF0
FAC5
FB25
FBAB
FB8A
FAC3
FA97
FC66
0010
03D0
05CD
05BE
04E6
049B
0505
055C
051B
049E
048F
04FF
055F
0544
04E8
04C6
04EA
04F7
04CC
04C5
0521
057D
053C
0484
0439
04C9
052F
03CF
005A
FC7D
FA55
FA62
FB46
FB8A
FB16
FAC6
FB0A
FB61
FB3E
FAD1
FAAE
FAF1
FB2C
FB1C
FB07
FB38
FB74
FB4A
FACF
FA9F
FB03
FB6E
FB25
FA6B
FA91
FCAB
0043
0397
052F
0516
0482
0479
04EE
0533
04F6
049A
049F
04FB
0538
0518
04DB
04D8
04FF
04FC
04BC
0494
04BB
04F1
04DC
04AD
04F4
05A3
0597
0396
FFD3
FC25
FA67
FABB
FBA3
FBB8
FB06
FA8A
FAC9
FB49
FB64
FB2A
FB1B
FB59
FB76
FB27
FAC2
FACB
FB35
FB72
FB45
FB1B
FB5C
FBAC
FB4E
FA5F
FA3F
FC48
002C
03E6
0596
0538
0465
0471
0531
0595
0522
0470
0441
0495
04DB
04D1
04C5
04FD
0538
0512
04A7
0479
04B4
04E4
04A1
044C
04A0
057D
058E
0385
FFB7
FC19
FA72
FAC1
FB8A
FB8F
FAF6
FAA8
FB03
FB81
FB8A
FB38
FB11
FB3F
FB65
FB36
FAE8
FADD
FB14
FB35
FB27
FB3D
FBA2
FBE1
FB67
FA86
FA9B
FCCB
009D
0422
05B1
0557
047E
0455
04C2
04F9
04B2
046D
04A2
0516
052D
04C8
046E
0492
04FB
051D
04D9
049B
04B2
04DD
04BD
0483
04BA
054D
051C
0301
FF43
FBB5
FA1B
FA89
FB8D
FBD3
FB57
FAF3
FB1E
FB75
FB76
FB35
FB1C
FB41
FB4F
FB1D
FAFC
FB3C
FB9A
FB8C
FB0B
FAB9
FB07
FB7E
FB52
FAA6
FAD9
FD23
0104
046F
05B2
050E
042C
0441
04FF
055A
04F3
0463
044D
0495
04BC
04A7
04AA
04E8
0508
04C8
0478
04A0
0527
0556
04D3
0445
048F
056A
0547
02EB
FF00
FBAA
FA7B
FB0E
FBC2
FB99
FB04
FAF4
FB83
FBEF
FBAD
FB16
FADC
FB1D
FB59
FB35
FAF8
FB0F
FB5E
FB67
FB0E
FADE
FB3F
FBB7
FB75
FAA1
FAB0
FCF3
00E4
0461
05B5
0533
0484
04A2
0507
04CF
0416
03C4
043F
04EA
050B
04C7
04C7
0529
0556
04EF
0471
048C
051E
0551
04D0
0456
04BA
059B
0567
02F7
FEF3
FB65
F9E5
FA56
FB54
FBB3
FB6D
FB33
FB6C
FBC6
FBC2
FB64
FB14
FB09
FB09
FADF
FAC5
FB0B
FB7F
FB89
FB04
FA9B
FAF0
FB93
FB78
FA9D
FA9D
FD12
016D
0526
063C
0532
0428
045B
0515
051D
0473
0412
046C
04E1
04CA
0475
049A
0537
0582
0512
0479
047E
04FF
052A
04B7
0469
04F6
05C8
0540
0270
FE56
FB1C
FA1C
FAC9
FB84
FB60
FAD5
FAD2
FB75
FBF0
FBA5
FAF2
FAB2
FB1C
FB8A
FB5D
FADA
FABE
FB37
FBAA
FB8C
FB1F
FAF9
FB1B
FAFE
FAAC
FB35
FD9A
015A
0490
05BD
0534
0486
04AB
0532
0531
049B
0437
0485
051C
054F
050F
04DB
04EF
04F2
049D
044D
048D
0535
056E
04CB
040E
0443
0532
0528
02BE
FE9A
FB10
F9DA
FA8E
FB6F
FB70
FAFF
FAF1
FB44
FB59
FAFB
FAB0
FAE7
FB52
FB62
FB16
FAF9
FB3C
FB65
FB06
FA88
FAB6
FB98
FC2E
FBAB
FAB8
FB16
FDC4
01C8
04F5
05F1
0547
0489
04A5
053C
0577
0521
04C4
04D1
0512
050C
04B6
0485
04C1
0522
0534
04F6
04C9
04D9
04E0
04B1
049F
04FE
0550
0460
0195
FDE6
FB25
FA49
FAAD
FB0B
FAE2
FAA9
FADA
FB3D
FB56
FB1B
FAEE
FB00
FB12
FAEF
FAC5
FAE4
FB3A
FB64
FB36
FB02
FB27
FB80
FB87
FB0E
FABE
FBA1
FE2D
01A9
049E
05F1
05BF
0517
04E9
0538
055B
04F4
046D
046C
04F7
056E
0554
04DF
049D
04BD
04F6
0506
04F5
04D8
04A0
0464
0498
056D
0603
04D3
0159
FD17
FA6C
FA3F
FB41
FB95
FAE6
FA62
FADD
FBB9
FBD2
FB0E
FA65
FA8F
FB2E
FB7D
FB55
FB26
FB32
FB47
FB42
FB42
FB45
FAF9
FA72
FAB2
FCE3
00C5
0468
05EF
0561
0469
0459
04F5
0541
04F5
04A4
04BC
04FC
04FF
04D4
04C2
04C7
04B4
049E
04BE
04EE
04C3
045C
047F
0571
05F7
0457
006B
FC45
FA33
FA7C
FB7A
FBB5
FB49
FB15
FB47
FB58
FB14
FAEB
FB27
FB6F
FB5E
FB2E
FB4E
FB94
FB6A
FADC
FAB5
FB51
FBD3
FB40
FA3C
FACC
FDFF
0261
054F
05AB
04B0
042C
0485
04E9
04D5
04A8
04D1
050E
04F1
04A1
0493
04B4
0481
03F2
03C1
0460
052B
0530
0498
0482
053C
0554
0329
FF21
FB94
FA56
FAEB
FB93
FB79
FB2D
FB45
FB6E
FB2B
FAD2
FB05
FB96
FBB1
FB36
FB06
FBAD
FC62
FC18
FB1E
FAC8
FB78
FBF4
FB44
FA84
FBD8
FFA2
03AA
058E
053E
0482
0487
04DA
04B7
0462
0491
052F
0564
04DD
0439
0417
043E
042C
0404
0440
04BB
04B7
0412
03C0
0484
0582
04D5
01BB
FDB0
FB03
FA84
FB16
FB56
FB16
FB02
FB59
FB90
FB38
FAA7
FA86
FAF8
FB83
FBC0
FBC1
FBBD
FBAD
FB8A
FB95
FBF3
FC31
FBAD
FAB8
FAD0
FD29
010D
044A
055E
04E2
047C
04D8
053E
0505
0496
04AB
0521
0542
04F0
04C7
050D
0526
048C
03CA
03CB
0470
04A5
0410
03B7
0464
0506
03A7
0005
FC46
FAA4
FB0F
FBAC
FB5A
FAB8
FABC
FB38
FB5D
FB17
FB07
FB4C
FB41
FAA0
FA31
FABF
FBD5
FC40
FBBC
FB53
FBC3
FC50
FBDD
FAEA
FB6B
FE6E
028B
0544
059E
04D5
0484
04E7
0527
04E5
04A3
04D8
0530
0522
04C5
04A2
04D6
04EE
04A6
045A
046B
0497
0464
0402
042C
04E4
04D5
02A3
FEBF
FB50
FA14
FAB4
FB83
FB80
FB1A
FB14
FB5E
FB5E
FAFC
FAB5
FAD0
FB03
FB0B
FB1D
FB6D
FBAE
FB80
FB2B
FB56
FBEA
FBF4
FB14
FA93
FC40
0029
0424
05F4
058A
049E
047A
04DC
04F2
04B0
049E
04D7
04ED
04BF
04B6
0504
0521
04A6
041D
0462
0541
057C
0489
038F
03EF
0517
04B7
0185
FD11
FA40
FA2C
FB4C
FBA8
FB13
FABB
FB27
FB99
FB5C
FADB
FAE8
FB74
FBB4
FB65
FB22
FB5B
FB96
FB3B
FAAD
FAD7
FBAC
FC05
FB5D
FB0E
FCF5
00F9
04BB
0616
0553
0474
04A6
053D
052B
0499
0472
04EC
054B
0507
0482
0453
0470
046E
0454
0482
04E3
04E6
047A
0464
0513
0577
03E4
0032
FC59
FA7D
FAB9
FB67
FB46
FAAE
FA90
FAFF
FB4E
FB33
FB13
FB2F
FB3E
FB0F
FB07
FB82
FC0C
FBDE
FB20
FAE2
FB8D
FC0D
FB47
FA10
FABC
FE4B
02DD
0586
0571
046D
0469
0551
05C6
0545
04AF
04C5
0520
0505
049A
048E
04ED
04FD
0476
0411
0471
0510
04FB
0458
0454
0541
0589
035D
FF25
FB6E
FA37
FAF2
FB96
FB27
FA74
FA79
FAFB
FB1E
FAC8
FAAB
FB1C
FB97
FB93
FB4C
FB48
FB79
FB68
FB16
FB0F
FB79
FBA5
FB1C
FABE
FC15
FF6C
031D
052D
054B
04BF
04AD
04FF
0515
04EA
04F2
0543
0562
050C
04A0
0484
0492
0472
044F
0499
0526
0535
048B
0407
0487
055D
04AE
019C
FD98
FB01
FAB4
FB73
FBA8
FB20
FAB7
FADB
FB19
FB00
FAD4
FB00
FB5F
FB79
FB49
FB3C
FB73
FB7D
FB21
FAE5
FB4F
FBE7
FBA3
FA97
FA76
FCD7
0119
04B3
05C6
04E6
0415
0461
051E
054C
04F6
04CF
0508
0527
04E5
04A1
04B4
04E2
04C6
0485
048F
04D2
04C5
0463
0472
054D
05CF
043E
006E
FC69
FA70
FABD
FB9E
FBAA
FB1B
FAE1
FB22
FB3D
FAF1
FAC0
FB0B
FB70
FB66
FB0F
FAF8
FB32
FB47
FB17
FB1E
FB93
FBC5
FB09
FA22
FAE4
FE1B
024D
050F
0578
04BA
0468
04C0
0502
04D6
04B9
0509
0562
053E
04C4
0488
04B5
04E8
04DF
04D6
04FC
04FA
0483
0416
048A
059F
05AA
0341
FF12
FB85
FA54
FAF4
FB98
FB57
FACF
FAD4
FB39
FB44
FADD
FAA5
FAF3
FB5B
FB62
FB2D
FB26
FB47
FB39
FB11
FB49
FBD0
FBCB
FAD6
FA29
FBA8
FF8E
03B7
05BB
0562
047D
0480
0516
052C
04AF
047D
04F2
0562
052D
04A9
048B
04D0
04EA
04B8
04B3
04FA
04FE
0471
040E
04AA
0596
04E3
01A4
FD5F
FAA5
FA5E
FB2E
FB70
FB07
FAE2
FB4C
FB90
FB31
FAB1
FAC4
FB45
FB7E
FB42
FB1B
FB56
FB89
FB4C
FAFB
FB2A
FB93
FB61
FAA0
FAD3
FD58
017E
04DF
05D1
0504
045A
04AF
0540
052B
04AC
0494
0503
0550
0514
04B0
049B
04B1
0493
0464
048E
04F7
0505
049C
047B
0513
0562
03BF
FFF7
FC0A
FA36
FAAA
FB98
FB83
FAC3
FA8E
FB2A
FBB9
FB8F
FB02
FABC
FADA
FB09
FB2F
FB6A
FB97
FB64
FAFF
FB13
FBC1
FC1F
FB62
FA61
FB1B
FE6B
02AD
0552
0588
04BF
049F
0526
0546
04AD
0431
047A
051B
0549
04FE
04D0
04F3
0503
04CB
04AC
04E2
04EF
0459
03B0
0407
0536
056D
0313
FEDE
FB55
FA26
FAA4
FB15
FAE3
FAD7
FB71
FC05
FBBB
FAE2
FA84
FAF6
FB75
FB57
FAED
FAE6
FB3C
FB60
FB41
FB64
FBE7
FC09
FB4E
FAB4
FBF9
FF7D
0377
05B6
05D3
052D
0500
0530
050E
0499
0471
04C6
0513
04F6
04BA
04C5
04EC
04C8
047B
0487
04E2
04DD
043F
03E2
049A
05A2
04FE
01C6
FD80
FAAB
FA33
FADE
FB25
FAD7
FABB
FB18
FB6E
FB61
FB3C
FB4F
FB5F
FB25
FAF3
FB4A
FBEC
FC03
FB5F
FADD
FB37
FBCC
FB6B
FA46
FA49
FCF8
0163
04E8
05ED
0542
04B4
04EF
053E
0508
04A6
04B0
04FD
04F9
0491
044E
0471
0490
0450
040C
0455
04FC
053B
04D9
049E
051E
057D
040F
006A
FC4E
FA03
FA14
FB13
FB80
FB42
FB22
FB5F
FB7D
FB32
FAED
FB1B
FB76
FB7A
FB34
FB2A
FB6F
FB81
FB2E
FB0A
FB81
FBF7
FB85
FA9D
FB18
FE1F
0272
0576
05E7
04E7
044A
048F
04ED
04D7
04A5
04BF
04F7
04F1
04CE
04E4
0516
04F8
0495
047A
04D1
04F3
0465
03CA
042A
053F
053D
02C5
FEAF
FB63
FA67
FB0B
FB9A
FB58
FAE7
FAFC
FB67
FB8C
FB4A
FB07
FB03
FB11
FB04
FB07
FB40
FB79
FB5E
FB1E
FB3E
FBC0
FBE3
FB3B
FABD
FC0C
FF7F
035F
0588
0593
04EC
04E1
0540
0520
0474
0419
0481
0516
052C
04EF
04E2
04FE
04E0
0497
049B
04E9
04DF
0453
0424
04FE
05D7
04AE
010F
FCFC
FACC
FAB8
FB28
FB02
FAAC
FAE4
FB74
FBA2
FB53
FB0C
FB05
FAF6
FAD0
FAF1
FB5E
FB81
FB1D
FADC
FB50
FBD7
FB7B
FAB8
FB6D
FE93
02BA
0570
05DE
0547
050F
0538
0520
04CA
04AE
04CB
04C2
04A1
04CC
0530
0537
04B7
044C
0476
04D1
04BE
0483
04D3
053A
0416
00B9
FCB9
FA65
FA43
FAEC
FB19
FADE
FADB
FB15
FB1D
FAF5
FB07
FB56
FB6D
FB2D
FB0E
FB4A
FB7A
FB56
FB41
FB7B
FB77
FAD1
FA88
FC45
002B
042A
0603
059A
04AC
0484
04DA
04EE
04C9
04D1
04EC
04CA
0496
04A9
04D9
04BC
0477
048D
04F4
04FF
048A
0472
0532
057C
0365
FF0D
FB13
F9B7
FA7F
FB57
FB4C
FB12
FB49
FB8F
FB64
FB19
FB34
FB7D
FB62
FB03
FB07
FB6E
FB80
FB10
FAE7
FB55
FB78
FAC8
FAA6
FCFE
017E
0563
0675
055D
046E
04B0
0534
0502
0483
0483
04D6
04DD
04A4
04A5
04D9
04D6
04A3
04A6
04D8
04C2
0474
04A8
0568
0538
0290
FE21
FA97
F9B6
FA96
FB3D
FB0F
FAD8
FB10
FB45
FB1B
FAE8
FB05
FB37
FB2B
FB0C
FB2E
FB60
FB42
FB14
FB64
FBDD
FB85
FA91
FAF0
FE00
026A
0560
05BF
04F3
04C6
0542
055D
04E0
049F
04FE
0557
051E
04C0
04C2
04E8
04C6
0495
04B0
04C3
0460
0408
048E
056C
04AE
014F
FCF6
FA6E
FA83
FB6F
FB6B
FABD
FA9C
FB22
FB6A
FB23
FAE6
FB15
FB55
FB4C
FB29
FB2E
FB34
FB1B
FB3B
FBC2
FBF9
FB24
FA31
FB4D
FF2A
039E
05DD
0589
0495
048A
050F
0524
04C1
0495
04CA
04DF
04A1
047A
04A1
04BE
04A9
04B7
04F4
04CC
0424
03F6
04E7
05B8
044C
0059
FC28
FA2C
FA7A
FB3E
FB42
FAF9
FB1B
FB67
FB57
FB24
FB48
FB8E
FB81
FB42
FB49
FB79
FB55
FAFA
FB15
FBA4
FBA1
FAA3
FA2F
FC48
00A0
047D
05C8
053B
04D0
051A
0536
04C2
046F
04B7
050B
04D4
046B
0478
04CE
04BF
045F
0466
04D6
04D4
044A
0464
058A
05EE
0378
FEC7
FAE6
F9E7
FACF
FB5E
FAEF
FA9C
FB0D
FB88
FB58
FAF5
FB0E
FB5B
FB49
FB0E
FB34
FB87
FB6F
FB1D
FB4D
FBE2
FBC9
FAC9
FA98
FD11
018A
052D
0625
056B
04F7
0538
054F
04E4
0493
04AD
04CE
04B2
04B0
0501
0533
04E5
048A
04BE
051F
04C9
03FC
03FA
04DC
04B7
01F2
FDB5
FAC1
FA3B
FAC9
FACD
FA5D
FA79
FB26
FB7F
FB3B
FB13
FB66
FB96
FB31
FAD3
FB11
FB6E
FB36
FAD1
FB1A
FBC9
FBBF
FB0E
FB92
FEA2
02E9
059B
05B0
04D6
04E2
0599
05B1
04FF
047D
049F
04DE
04CD
04AF
04C8
04DB
04B6
04AA
04FD
053C
04E0
0462
04A7
0535
042B
00AB
FC75
FA20
FA35
FB0A
FB20
FAA5
FA7C
FACB
FB12
FB23
FB40
FB69
FB51
FB16
FB3B
FBAA
FBA4
FB05
FAB7
FB41
FBB4
FB1D
FA7D
FBF9
FFFC
0435
0615
059C
04D3
04F9
0566
0541
04F0
051B
0565
0516
0476
0455
04B3
04CC
0475
0463
04E2
0534
04C8
0461
04DF
0553
039C
FF65
FB39
F9AC
FA78
FB58
FB22
FAAE
FAE7
FB62
FB48
FAC3
FAA3
FB11
FB6C
FB6A
FB6B
FB94
FB7A
FB0F
FAFB
FB70
FB8A
FACB
FA8E
FCB9
0116
050A
0662
059B
04D2
0507
0567
0515
0477
0456
04A1
04D0
04D7
04F5
0502
04C1
0481
04B0
0501
04CC
0442
0463
0550
055B
02CE
FE63
FADB
F9E9
FA8E
FAE7
FA9E
FA98
FB1E
FB8A
FB84
FB75
FB9E
FB9B
FB29
FACB
FB04
FB64
FB31
FABA
FAFA
FBC7
FBC9
FAC9
FAC8
FD9E
0233
0578
05F5
051E
04FA
0599
05B3
04F0
0453
047D
04C8
0490
0442
0479
04DF
04D7
049C
04CE
0537
051F
04A3
04AD
0535
049B
0191
FD40
FA5F
FA20
FB0D
FB3F
FAAD
FA7C
FAFA
FB67
FB5C
FB42
FB6E
FB99
FB81
FB5E
FB6D
FB6D
FB1E
FADB
FB16
FB66
FB06
FA80
FBA4
FF33
035F
05A0
0579
049F
048C
050A
0537
04FD
04EE
0524
051E
04B6
0462
0465
046F
0456
0476
04E6
050D
04A6
047F
053A
05CA
0442
0059
FC3B
FA4B
FAA2
FB70
FB73
FB14
FB0E
FB31
FB02
FAC2
FAEB
FB46
FB50
FB29
FB4D
FB9C
FB76
FAE3
FABE
FB54
FBB1
FB09
FA7B
FC1C
0020
0419
05AE
052F
0492
04C4
050E
04D2
0485
04C1
0536
053A
04D9
04AA
04D1
04DB
04AB
04AA
04EC
04EE
04A3
04C8
0583
0564
02F2
FED6
FB86
FA90
FB23
FB7F
FB28
FAEA
FB30
FB6B
FB34
FAF9
FB17
FB29
FADC
FAB4
FB30
FBCA
FBAF
FB21
FB15
FB8F
FB6D
FA6B
FA52
FD0B
01C7
0569
0603
04D6
0441
04C7
0530
04D7
046F
049F
0509
050E
04D3
04DE
0525
0523
04C4
047A
0475
046D
046A
04E1
0587
04DE
01E7
FDC9
FAE2
FA4F
FB09
FB86
FB62
FB35
FB53
FB70
FB55
FB37
FB31
FB0E
FADB
FB00
FB78
FB9D
FB34
FAF5
FB6C
FBDB
FB4B
FA66
FB3A
FEB0
0302
0583
0582
049C
045F
04A6
04A7
046D
047C
04BC
04BF
04A5
04E5
054D
0530
0487
042C
0496
050D
04CA
0456
04B7
055E
044B
00BD
FCAF
FAA7
FAD6
FB74
FB58
FB0F
FB56
FBC7
FBA3
FB21
FB0B
FB68
FB74
FAF9
FAB8
FB1F
FB8E
FB6A
FB1F
FB40
FB64
FAF6
FABF
FC67
0025
03F0
0593
0517
0452
046E
04DA
04C0
0463
0473
04D9
0508
04F4
04F2
04F4
04B6
0473
04A1
050D
04F8
045E
044B
053B
05B0
0396
FF27
FB31
F9FF
FAE8
FBB0
FB71
FB0D
FB49
FBB7
FBB1
FB59
FB29
FB1B
FAEA
FAC5
FB13
FB8E
FB82
FB02
FAF1
FB7B
FB96
FAC8
FA8F
FCCD
011C
04E1
0622
056E
04A1
0495
04C5
04BA
04B5
04DD
04CA
0461
0444
04C7
0540
0506
0493
04BB
053D
052C
048D
0481
054B
053D
0298
FE25
FABA
FA00
FAD4
FB43
FAFD
FAF3
FB64
FB97
FB3C
FAEC
FB1B
FB70
FB76
FB56
FB63
FB67
FB08
FAA3
FAD6
FB4A
FB03
FA41
FAF2
FE45
02B1
0571
05A7
04E4
04C7
052F
0529
04AB
047D
04CE
04F9
04BF
04B5
0519
0541
04C6
045A
04B3
0542
0521
04A4
04E1
058D
04AF
0128
FCAE
FA33
FA7D
FB96
FB94
FACE
FA9A
FB1B
FB66
FB26
FAF1
FB15
FB2D
FB04
FB00
FB58
FB86
FB1C
FAA4
FADA
FB50
FB07
FA75
FBA4
FF7A
03EE
0614
0577
0443
044C
0523
0568
04F3
04B7
0512
0554
050E
04C8
0500
053F
04E6
044A
042C
048E
04D4
04D8
04F3
04E1
0380
004E
FC97
FA70
FA7E
FB68
FBAB
FB34
FAD9
FAEF
FB0D
FAEF
FACA
FAD1
FAF4
FB19
FB40
FB50
FB27
FAFB
FB41
FBEA
FC22
FB69
FAD2
FC3B
FFF4
03EE
05D5
0584
04BB
04BC
0520
0507
0493
0485
04F5
0536
04FA
04C0
04E6
04FF
0493
0411
043D
04EA
051D
0492
0444
04F6
05A7
0467
00C5
FCAB
FA74
FA80
FB43
FB5F
FAF9
FAE7
FB48
FB81
FB4A
FB0E
FB28
FB53
FB2D
FAEC
FB19
FBA4
FBDA
FB6E
FB05
FB4D
FBD9
FBA5
FAC5
FADF
FD64
0195
04FC
05EF
0520
046B
04A7
0523
050E
0498
046D
04A8
04D7
04C6
04B4
04C5
04C0
048C
047C
04C8
0506
04AC
0416
0444
0552
05BD
03CD
FFBB
FBCF
FA1E
FA8C
FB5D
FB55
FACD
FAB7
FB35
FB9B
FB80
FB36
FB34
FB6F
FB8F
FB82
FB7A
FB7F
FB66
FB37
FB3B
FB74
FB5C
FAAC
FA35
FB6E
FECA
02CD
0553
05A5
04F2
04AF
0508
0534
04D9
047A
048F
04CF
04B9
046C
0469
04B0
04BB
0461
0433
0499
051A
050A
04A7
04D2
057F
052B
028C
FE69
FB23
FA37
FADE
FB5B
FB14
FACA
FB14
FB81
FB6E
FB0B
FB02
FB67
FBA0
FB61
FB1E
FB47
FB8C
FB5F
FAEC
FAE7
FB61
FB7B
FAC9
FA75
FC39
0022
040E
05C9
0550
047A
049E
0542
0551
04C5
0489
04F4
054F
04FA
0465
0460
04DF
051E
04D3
048A
04B3
04E7
04B1
047C
04F7
0592
0492
012D
FCF6
FA70
FA61
FB4C
FB82
FB00
FAC7
FB24
FB5C
FB04
FAAD
FAF2
FB72
FB6D
FAF4
FACE
FB39
FB8F
FB4E
FAEA
FB08
FB5E
FB1D
FA78
FAFD
FDC9
01DE
04EF
05BE
0525
04AF
04CF
04E8
04A4
0474
04C0
052A
0523
04C8
04B1
04FC
051D
04C4
0471
04B8
0546
054B
04C0
0491
0525
054D
0367
FF86
FBC8
FA2E
FA9B
FB59
FB50
FAF5
FB17
FB8B
FB98
FB26
FADA
FB05
FB3D
FB20
FAFD
FB3B
FB8A
FB50
FAB8
FAA3
FB47
FBA2
FAF4
FA44
FB8F
FF4B
037A
05AB
057D
049A
047E
04FA
0513
049A
0441
0475
04D4
04E2
04BB
04C0
04EE
04F6
04CE
04C4
04F1
04FF
04C0
04A8
0530
05C7
04F2
01EA
FDD2
FAE2
FA3E
FAFE
FB78
FB24
FAD3
FB37
FBD6
FBD1
FB38
FAEF
FB56
FBC2
FB7E
FAE1
FAC1
FB3A
FB92
FB5B
FB0D
FB20
FB2E
FAC1
FAA7
FC74
0054
043C
05F4
057B
04B3
04D8
0549
04FC
0439
0419
04BE
0521
04B1
042D
0469
04FC
04FA
0475
0458
04D4
0502
0469
0401
04CB
05D9
04E1
0121
FCAE
FA45
FA5E
FB28
FB27
FAB2
FAC8
FB5E
FB97
FB38
FAF4
FB3E
FB94
FB62
FAF8
FB0A
FB85
FBAA
FB4F
FB34
FBC9
FC3F
FB91
FA5B
FAAC
FDB6
021A
0530
05C2
04F8
048E
04DF
0517
04CF
0492
04D9
0539
0513
0498
0482
04F5
0537
04CE
0439
0432
048F
0492
0430
0444
0519
0564
037F
FF93
FBCF
FA2F
FA8D
FB44
FB4A
FB05
FB1D
FB62
FB3F
FACB
FAAF
FB19
FB72
FB50
FB19
FB57
FBCA
FBC4
FB45
FB1A
FB9B
FBFB
FB6C
FAB1
FBA4
FEF9
0308
056E
058A
04D5
04C9
0543
0544
04A7
0451
04C9
056A
0559
04BC
0466
0496
04BD
0485
0462
04B7
050A
04B8
041F
0445
0513
04D7
0228
FDFB
FAEB
FA5B
FB25
FB61
FAC8
FA87
FB2D
FBCF
FB85
FAC8
FAB3
FB57
FBB7
FB52
FAE2
FB22
FBA7
FB9A
FB1E
FB1E
FBB3
FBD1
FAF9
FA96
FC90
00BB
0491
05E8
0530
047A
04CD
0551
0512
0476
0475
0504
0531
04A8
0437
048A
051C
050A
0474
0449
04C3
0505
0483
0410
04A6
0586
0495
00F8
FC8E
FA1A
FA4D
FB67
FBA2
FB1A
FAF2
FB6A
FBA1
FB25
FAA6
FAE1
FB7C
FB9E
FB3E
FB18
FB71
FBA5
FB3D
FACC
FB15
FBB8
FBA2
FAD8
FB0B
FDA7
01D4
0511
05DC
0511
047C
04BF
0514
04DE
0480
049F
0516
0543
04F8
04A8
04A2
04AB
0488
0479
04C8
052B
0516
04A2
0493
0523
0533
034D
FF88
FBD9
FA36
FAA0
FB70
FB62
FAC9
FAA6
FB26
FB86
FB44
FACD
FAC7
FB28
FB6C
FB64
FB5C
FB70
FB55
FAFA
FAD4
FB25
FB5F
FAE4
FA65
FB9B
FF38
0385
05E5
059F
0474
0450
0523
0588
04F8
045C
048E
0529
0549
04EA
04B9
04EA
04F8
04A6
047E
04DF
0536
04E3
0465
04C7
05B8
054C
022B
FD9A
FA6D
FA09
FB20
FBA1
FB1D
FAA6
FAE5
FB4F
FB3F
FAFD
FB22
FB86
FB7D
FAFC
FAC1
FB2E
FBA1
FB66
FAD6
FADC
FB72
FB85
FAAC
FA54
FC56
0088
047B
05F5
0538
0456
04A0
0574
059E
050D
04A3
04C3
04E4
0499
044B
048A
0514
0533
04D0
0492
04CD
04FC
04AC
0464
04DE
057F
047E
0116
FCEA
FA84
FAA0
FB9E
FBB1
FADE
FA62
FAC6
FB4C
FB44
FAFF
FB17
FB67
FB56
FAE7
FABF
FB16
FB5D
FB27
FAEE
FB4C
FBD5
FB8F
FAAA
FAEC
FDB4
01FE
0527
05B3
04AF
041E
049D
0533
0511
049E
04A5
051C
055E
0533
0507
051A
051D
04D2
0497
04D0
0521
04DC
042B
0415
04EF
0559
0387
FF8B
FBA4
F9FE
FA89
FB7B
FB93
FB2E
FB28
FB7C
FB7C
FAFF
FA9B
FAB2
FAEE
FADB
FAAA
FACE
FB38
FB66
FB3B
FB2F
FB79
FB8B
FAFF
FAA8
FC07
FF6D
0336
0554
055C
04A5
0481
04E9
051B
04E6
04C9
0504
0531
04FE
04C3
04FB
0572
0581
0502
0491
049D
04CB
049C
0463
04D8
05AB
0532
023F
FDE4
FABA
FA37
FB4B
FBE7
FB58
FA96
FA93
FB04
FB24
FAED
FAEC
FB34
FB3C
FADE
FAAF
FB0F
FB7A
FB50
FAEB
FB21
FBCB
FBBA
FA95
FA0B
FC25
0094
0498
05EB
0511
0441
049A
0553
0566
04FC
04D6
0504
0503
04C1
04C2
0529
0553
04DF
0464
04A2
053F
053A
047E
0433
0506
05BD
0458
008D
FC7A
FA7B
FAC5
FB9A
FB8D
FADD
FA8E
FADB
FB24
FB06
FADC
FB0C
FB5B
FB53
FB05
FAF3
FB3C
FB5F
FB0D
FAC0
FB05
FB79
FB3F
FA8F
FB0C
FDF6
0242
0558
05C4
04A6
041B
04BF
0573
0550
04D4
04DC
0545
0543
04B5
0450
047E
04CA
04BF
04AA
0504
0575
0540
0491
047B
0541
0562
032C
FF09
FB64
FA19
FAAD
FB4D
FB12
FA9B
FAB2
FB2A
FB5C
FB30
FB16
FB39
FB4D
FB2F
FB29
FB68
FB91
FB40
FABF
FAB7
FB37
FB71
FAE3
FA75
FBCD
FF5E
0383
05F3
0603
050D
04B0
0524
0579
051E
048B
046B
04AF
04D2
04B2
04A8
04CE
04D5
04A5
04A1
04FA
0539
04E7
047B
04CC
0586
04F3
01F1
FDB3
FAD0
FA72
FB45
FB63
FAA0
FA36
FAC4
FB83
FB96
FB34
FB1A
FB5C
FB6C
FB21
FAFA
FB3E
FB81
FB5D
FB31
FB7E
FBE9
FB97
FAA3
FA86
FC93
004F
03C1
0563
0561
04F2
04E1
050D
051B
0506
04FC
04FC
04DA
0493
045A
0461
0494
04B1
049F
0494
04C4
04FF
04D4
043A
03E5
048F
05C9
05E4
037C
FF2D
FB5E
F9FD
FABB
FBB4
FBA5
FAFA
FAC0
FB1F
FB58
FB04
FAAC
FAF7
FBA4
FBE6
FB81
FB1B
FB48
FBC1
FBD0
FB5C
FB10
FB5A
FBB4
FB4F
FA6B
FA7F
FCC6
00B5
0448
05D9
0588
04C0
0497
04F1
051D
04E1
049F
049B
04A2
0478
0453
048E
0502
0513
0486
03FA
0433
050B
0580
04FC
0434
044B
0531
054A
031B
FF1A
FB79
FA05
FA8B
FB61
FB5E
FAD4
FAB3
FB35
FBBA
FBBF
FB7F
FB74
FB96
FB77
FAFF
FAAB
FAE1
FB58
FB7B
FB3C
FB2E
FB99
FBE6
FB53
FA4A
FA6E
FCFE
013E
04E0
0627
056F
0478
046C
04EC
050C
04A8
0467
04A7
04F7
04CF
0467
0467
04EE
0554
0513
0486
0466
04C1
04E5
0476
041A
04A2
05A3
0573
02E5
FEC1
FB45
FA07
FAA4
FB7A
FB7E
FB01
FAD4
FB1A
FB44
FAFE
FAAD
FAE0
FB7B
FBCF
FB7A
FAEC
FAC5
FB0D
FB3F
FB22
FB1F
FB89
FBE6
FB78
FA8E
FAB5
FD2E
0145
04B4
05D5
0527
0470
04A9
053E
053E
04BB
0482
04DD
052D
04E1
0455
0453
04F1
056A
0533
04B4
04A6
0503
050B
0471
03F6
0475
0576
0540
02A7
FE84
FB23
FA13
FAD4
FBA9
FB87
FAE2
FABA
FB3A
FBA6
FB71
FAF2
FAD8
FB33
FB6C
FB25
FAC5
FADC
FB4B
FB6B
FB10
FAD5
FB38
FBB8
FB72
FA9A
FACB
FD55
017E
04E8
05E7
0510
0440
0479
0519
051A
0485
0437
049D
052D
0535
04C9
048C
04C2
0503
04ED
04B4
04C4
0509
04FF
0489
0453
04EE
05B9
0518
022C
FE06
FAE8
FA22
FAFF
FBCA
FBAF
FB35
FB25
FB6C
FB64
FAEB
FAA0
FAFD
FB9C
FBB9
FB3B
FAD6
FB11
FB8D
FB94
FB21
FAE8
FB49
FBA8
FB3A
FA67
FACE
FD8C
01C1
0520
061C
0540
044D
044A
04CD
0501
04D2
04CC
0520
054F
04F1
045B
0436
0495
04DE
04A8
0448
044D
04A7
04BC
045B
042D
04D6
05C0
0553
0294
FE73
FB1D
F9FB
FA89
FB3A
FB2D
FAD2
FAE5
FB54
FB73
FB0B
FAAB
FAE0
FB70
FBB3
FB7F
FB4E
FB7C
FBC4
FBB9
FB7B
FB89
FBE2
FBD4
FAFD
FA33
FAFB
FDE6
01C9
04B7
05B8
0562
04F5
050A
0549
0533
04D9
04B1
04E3
0515
04E6
047C
0455
0492
04C7
0494
043D
044B
04B5
04CC
0448
03E2
0466
054E
04DE
0204
FDD8
FAB8
F9FA
FACA
FB71
FB3A
FAC0
FAB7
FB02
FB1D
FAF4
FAEF
FB48
FBAD
FBB0
FB5B
FB24
FB4A
FB8A
FB81
FB41
FB34
FB7D
FBA8
FB44
FAC9
FB89
FE5B
025F
057C
0653
0579
049A
04A0
0516
0531
04F1
04E3
051F
051C
0499
041B
043D
04C3
04EB
047D
0422
046B
04FC
050D
0490
0466
0517
05C8
04D1
018E
FD4F
FA40
F97E
FA49
FB1E
FB35
FAEE
FAE6
FB1D
FB24
FAE6
FACF
FB2B
FBA4
FBB0
FB52
FB17
FB53
FBA9
FB96
FB34
FB1E
FB7C
FBA0
FAF1
FA1D
FAD3
FE04
028E
0603
06DB
05BF
049B
0491
0529
0557
04E6
048C
04CA
053A
0530
04AB
044E
047B
04D9
04E9
04B7
04A5
04BE
04A6
0458
046A
052A
05B7
0490
0140
FD30
FA76
F9E7
FA98
FB22
FB15
FAED
FB0D
FB37
FB18
FADC
FAF4
FB5D
FB94
FB49
FADB
FAE0
FB57
FBA0
FB59
FAF5
FB1C
FBA9
FBBD
FB03
FA89
FBDD
FF3F
0318
056C
05B2
0509
04B4
04E4
0507
04E7
04DD
0520
0550
04FD
0466
043D
04BB
0547
0531
049A
0448
0499
0502
04CF
0431
041D
04F1
0594
0457
00DD
FCCF
FA64
FA46
FB2A
FB7E
FB06
FAA6
FAEB
FB54
FB31
FAAD
FA8F
FB16
FB9F
FB89
FB15
FAFB
FB5C
FB9D
FB5D
FB16
FB6E
FC1A
FC12
FB0A
FA4B
FB95
FF1F
031A
0564
058F
04ED
04D2
053D
0555
04D5
046A
04B5
0565
05A2
052D
04A3
0496
04D3
04C8
046A
0442
0495
04E6
04A3
040D
0409
04D9
0564
041F
00C9
FCF0
FA92
FA4B
FB09
FB68
FB1B
FAD6
FB19
FB83
FB6E
FAE2
FA8B
FACF
FB4B
FB70
FB42
FB3E
FB86
FBA9
FB5C
FB06
FB3D
FBCC
FBCD
FAF9
FA7B
FBEC
FF7B
0368
05A0
05A7
04C2
0467
04CC
0527
04F5
0497
04A4
050F
053C
04E3
046F
046A
04C5
04FC
04D7
04B1
04D7
04FD
04B1
0430
044E
0534
05A6
0412
0066
FC7D
FA65
FA72
FB3D
FB6A
FAF6
FAB4
FAFA
FB47
FB28
FAE9
FB14
FB9B
FBD9
FB76
FAEA
FADF
FB4E
FB87
FB32
FAD8
FB22
FBCC
FBD5
FAF6
FA6C
FBE0
FF75
0354
056A
0563
04A5
048A
050B
054E
04FF
04A5
04BC
050A
050C
04BD
0494
04CE
0513
04F8
049D
0480
04C4
04FC
04C2
045A
046E
0514
054C
03CE
0075
FCC0
FA8F
FA6E
FB3B
FB90
FB31
FAEF
FB4A
FBC5
FBA2
FAF4
FA82
FAAF
FB11
FB27
FB1A
FB50
FBAA
FB9A
FB11
FAC1
FB2B
FBBF
FB7F
FA7C
FA3C
FC35
000F
03C8
0598
0577
04B8
0475
04A9
04BD
0486
0470
04C4
0535
0547
0504
04E4
051A
0535
04C2
040D
03E2
047E
0526
0513
0493
04B5
05AA
0603
040D
FFE2
FBB3
F9BE
FA3E
FB88
FC05
FB9A
FB2B
FB33
FB51
FB1A
FAC4
FACB
FB2D
FB68
FB35
FAF1
FB17
FB8E
FBC5
FB82
FB39
FB58
FB88
FB16
FA25
FA11
FC2A
001E
03F0
05C8
058C
04A7
045B
04AE
04EE
04CE
04AB
04D5
050D
04F4
04A1
0485
04BC
04E3
04B1
0471
04A3
052D
055A
04D3
044C
04B7
05D6
0601
03CA
FFB5
FBFB
FA71
FAE1
FBA0
FB81
FADB
FAA6
FB15
FB7B
FB57
FB00
FB0D
FB75
FBA6
FB63
FB20
FB50
FBAC
FB87
FACE
FA4A
FA9A
FB47
FB46
FA78
FA40
FC21
FFE8
039A
0559
052C
0496
04B7
053E
0547
04BC
045C
049C
0503
04EF
0481
046B
04E2
054A
0518
049C
0490
0508
0555
050C
04BE
0530
060C
05D2
0368
FF83
FC26
FABE
FAF2
FB61
FB45
FAF3
FB04
FB62
FB81
FB3B
FB0D
FB58
FBC0
FBA1
FAF6
FA72
FA9B
FB16
FB2C
FACB
FA98
FAF9
FB63
FB0C
FA36
FA55
FCA1
0098
0437
05CD
056F
0489
0448
04A5
04E8
04C4
048F
04A3
04D6
04D1
04A9
04BC
0517
0549
0507
04AA
04C3
053F
0577
051D
04CE
053B
05F2
056C
02B2
FEA7
FB63
FA41
FACA
FB88
FB97
FB3E
FB29
FB6C
FB8F
FB4C
FAF8
FB03
FB50
FB54
FAE4
FA82
FABE
FB61
FBA2
FB35
FAC6
FB05
FB8D
FB61
FA85
FA85
FCC9
00B7
041A
056F
053B
04F9
0531
0545
04CA
0443
0453
04C2
04EE
04BB
049E
04D3
0510
0514
04FE
04FE
04F5
04CA
04BD
050B
0558
050B
045B
0432
04BA
049B
026F
FEAE
FB7E
FA6F
FAFF
FB95
FB72
FB19
FB19
FB42
FB36
FB18
FB2C
FB4C
FB28
FAE4
FADC
FB00
FAEF
FAAC
FABA
FB44
FBAC
FB67
FAEC
FB1E
FBD9
FBFF
FB49
FB35
FD5F
0144
0488
058E
04FF
048B
04CD
0512
04D4
0488
04BA
0525
0539
04FB
04E4
0510
0520
04EA
04B0
04A2
049B
0488
04A9
0506
0512
046C
03CF
045B
05B1
05A6
02A6
FDEB
FA7D
F9FC
FB31
FBEB
FB81
FAEE
FAF1
FB24
FAF7
FAA4
FAAE
FAFD
FB1E
FB0E
FB22
FB55
FB50
FB1C
FB34
FBAF
FBEA
FB70
FAD1
FAE0
FB54
FB23
FA68
FAE8
FDE9
0231
0517
0573
0496
044F
04D1
0522
04E4
04BE
0514
0564
0533
04DE
04F1
0537
051E
04B7
0492
04C2
04C6
047B
046D
04DD
0526
04AF
0428
04B6
05DD
0564
0203
FD64
FA84
FA6B
FB72
FBAF
FB14
FABF
FB08
FB3B
FAEE
FAA7
FADF
FB34
FB22
FADC
FAE7
FB29
FB24
FAE0
FAEC
FB61
FB9E
FB4B
FAF9
FB39
FB89
FB09
FA42
FB15
FE69
02A1
0530
055D
04A7
0492
050A
052C
04DA
04BC
050B
0541
050A
04CE
04E7
0508
04D2
0494
04CC
0537
0521
048C
0447
04B4
0522
04EB
04A3
052D
05DF
04B2
00E6
FC79
FA2F
FA87
FB93
FB9D
FAEB
FAA5
FAF1
FB05
FA9F
FA6B
FAD3
FB50
FB4D
FB10
FB20
FB5A
FB4A
FB12
FB39
FBA4
FB98
FAEF
FA84
FAEC
FB5D
FAD7
FA24
FB6A
FF59
03CA
05FC
059F
04AC
04A6
0529
053C
04F9
0519
0587
057D
04DF
0487
04E3
053D
04E8
0461
0480
050C
051B
0493
0461
04EC
055F
04F7
0460
04B2
0553
0433
0085
FC41
FA0B
FA4C
FB33
FB47
FAD1
FAB7
FAFB
FB09
FACD
FAC4
FB03
FB17
FAEA
FAFC
FB76
FBAA
FB23
FA85
FAB0
FB59
FB7A
FAED
FAB9
FB68
FBFC
FB70
FAB5
FBFC
FFCA
03E9
05D3
0574
04AD
04AD
04F1
04C7
0490
04FA
05AF
05B7
04F5
045B
0488
04FD
0508
04D2
04E1
051B
04FC
0498
0484
04D4
04E9
0486
046B
0516
0568
0398
FF9D
FBC2
FA3B
FAD0
FB95
FB6A
FAE3
FAD8
FB1E
FB13
FAC4
FAC2
FB1B
FB3E
FAF4
FABB
FAF0
FB33
FB1E
FAFF
FB46
FBAA
FB86
FAFD
FAE7
FB70
FBA8
FAFA
FA9B
FC6B
006A
0444
05D3
0561
04C8
04F8
0550
051E
04B9
04C2
0510
050D
04BE
04BF
0532
0579
0536
04DB
04DF
04F4
04A4
043F
046B
0500
0523
04AA
047E
051F
054F
034A
FF3A
FB83
FA2B
FAB7
FB3D
FAE5
FA79
FABB
FB3D
FB3D
FAE0
FAD9
FB42
FB71
FB0E
FA98
FA9C
FAF5
FB2C
FB36
FB46
FB43
FB01
FACE
FB1D
FBA4
FB87
FABC
FAC0
FD17
0139
04B9
05D0
051C
047C
04CD
0569
058F
0553
0521
04FB
04B5
0482
04B2
0514
051C
04C5
04A3
04F5
053B
0506
04C0
04F9
0561
052B
0470
0445
0504
052F
02FC
FEC9
FB1B
F9F1
FABB
FB82
FB52
FACB
FAAC
FAD8
FAE7
FAEA
FB1F
FB4B
FB0A
FA96
FA95
FB19
FB74
FB42
FAFD
FB22
FB57
FB10
FAA6
FADE
FB88
FB7F
FA86
FA54
FCC6
0149
050B
060A
0514
044D
048D
0507
0510
050A
0569
05C4
057A
04CD
048D
04E5
052D
0502
04CE
04F5
0525
04F4
04AE
04D8
0536
0524
04BE
04D5
0569
04FD
0242
FE1F
FB1E
FAA0
FB80
FBD2
FB36
FAB2
FADB
FB27
FB0F
FADF
FB08
FB46
FB13
FA9B
FA91
FB0B
FB53
FB04
FAA6
FACB
FB1F
FB0B
FAC2
FAF1
FB79
FB75
FAD4
FB0F
FD91
019D
04C8
0596
04E7
047B
04CF
0520
04F3
04B0
04B4
04BE
0488
046C
04DA
0582
05A1
051B
04A2
04AF
04EC
04F6
050A
056C
05AB
0536
0480
0496
055F
0515
0242
FDE8
FABD
FA3C
FB37
FBA7
FB16
FA8F
FAC2
FB36
FB49
FB1F
FB2D
FB69
FB6B
FB2C
FB04
FB0A
FAFA
FAD2
FAEC
FB44
FB49
FAC3
FA66
FAD4
FB6F
FB1E
FA3C
FACB
FE17
02AB
059B
05B1
0482
0429
04E9
059A
059C
0565
0556
0520
0494
0435
047E
0502
04FA
047F
046E
0510
0596
0554
04BC
0497
04CB
04C5
04A6
0519
05C8
0504
01BC
FD49
FA68
FA45
FB6C
FBCE
FB17
FA63
FA62
FAAE
FAC7
FACC
FAFC
FB25
FB08
FAE1
FB1C
FB97
FBC0
FB73
FB20
FB09
FAED
FABC
FAEC
FB9A
FBE0
FB03
FA06
FB17
FEE9
0365
05BC
056D
0479
049B
0568
0594
0506
04C1
052E
059C
057C
0531
0546
0573
051E
0474
043B
049F
04F2
04CE
04AF
0500
0541
04E2
0469
04C1
0569
047E
0106
FCA4
FA0F
FA1D
FB2B
FB72
FAF6
FAB9
FAEF
FAF6
FA9F
FA7B
FAD6
FB2B
FAFD
FA9E
FAA7
FB05
FB2A
FAFF
FB06
FB62
FB8F
FB52
FB33
FB84
FB98
FADD
FA55
FBE5
FFD5
03F1
05C3
0543
047E
04CD
0582
057A
04ED
04D8
054D
0578
050F
04C7
0524
05A0
0580
04F3
04C1
050C
052F
04DB
0486
0486
0480
0442
0468
0545
05A0
03B1
FF91
FBBB
FA76
FB54
FC05
FB4F
FA3D
FA34
FAFA
FB60
FB11
FABE
FACD
FAD8
FA94
FA60
FA9B
FAF7
FAF8
FACE
FAFE
FB5E
FB40
FAB4
FAB4
FB99
FC44
FBB7
FAFD
FC48
0013
0420
05E3
054A
045A
047B
0520
053A
04DB
04C7
0514
0538
050E
050D
055D
058E
0559
0520
0542
056D
0524
04B1
04C9
0549
0535
044E
03B8
044C
04E6
0377
FFB9
FBE0
FA2D
FA95
FB4F
FB47
FAF8
FB13
FB54
FB33
FAE5
FAEF
FB28
FAFF
FA82
FA61
FAD5
FB38
FAFE
FA8F
FA9A
FAF8
FB02
FAC8
FB10
FBDB
FC0B
FB26
FAB9
FCCC
0119
04E9
05FF
04F7
041C
0487
054F
0558
04DC
04B3
04F0
050A
04E9
04F8
0551
0583
0554
0518
0514
050B
04BA
047C
04C7
0543
0521
046F
0437
04D6
04E9
02CD
FEE2
FB74
FA48
FAE3
FB91
FB76
FB0B
FAE2
FAE0
FAC5
FACA
FB23
FB76
FB51
FAE7
FAC6
FAF5
FAFE
FAC5
FAC9
FB44
FBAB
FB6D
FAEC
FAFB
FB82
FB88
FAE2
FB08
FD70
016C
0499
056E
04BD
0453
04CF
0564
055E
050E
0507
0530
0516
04B7
047C
048E
04AF
04BF
04DF
050E
0505
04B3
047E
04B1
04F8
04D6
0488
04C0
0552
04CF
0221
FE2F
FB38
FA84
FB41
FBCC
FB85
FB00
FACE
FACC
FABF
FAD0
FB2A
FB75
FB4C
FAEB
FAEA
FB5C
FBB3
FB89
FB2D
FB1F
FB5B
FB78
FB50
FB19
FAE7
FA9A
FA85
FB98
FE59
01EE
04A9
0592
0523
0484
045D
049D
04F5
0538
054C
051F
04D9
04C1
04DD
04E3
04B2
0486
0491
049D
046F
0450
04B4
0562
0585
04D6
0439
04A5
0586
0500
0217
FE11
FB3C
FA89
FAFA
FB35
FAFE
FAEC
FB36
FB6C
FB3B
FAEC
FAE4
FB0D
FB0D
FAEA
FAFB
FB53
FB93
FB7C
FB4D
FB65
FB9F
FB78
FAD3
FA4B
FA80
FB38
FB8D
FB16
FAA9
FBA3
FE6E
01E5
0455
0503
04A9
0478
04DD
0558
055D
0501
04C1
04CE
04E9
04E0
04DC
0512
0551
0534
04B5
0455
047C
04EF
0523
04F8
04D4
04F8
0517
04DC
0499
04E2
0568
04D0
0222
FE3A
FB3B
FA77
FB32
FBBA
FB56
FAC2
FAD1
FB4D
FB78
FB2A
FAEB
FB0B
FB2F
FAF8
FAA7
FAC0
FB39
FB79
FB38
FAE6
FB01
FB58
FB57
FAF2
FAC5
FB1C
FB65
FAF6
FA4C
FAF2
FDDA
0200
0522
05E1
04F8
0432
0478
052E
0552
04D0
0470
04AF
052C
0546
04F8
04C6
04EE
0521
0510
04DF
04DB
04F6
04EB
04C1
04D5
052F
054E
04E5
0480
04E5
05B9
055C
029C
FE55
FAE0
F9CE
FA8B
FB5F
FB59
FAEE
FAE2
FB34
FB56
FB1D
FAED
FB0E
FB40
FB28
FAE8
FAEB
FB3F
FB6F
FB21
FAA3
FA89
FAEB
FB46
FB3A
FB10
FB34
FB6D
FB1E
FA75
FACC
FD58
0177
04E2
05E1
04FE
0433
0495
0562
0563
049A
0417
0477
0528
055A
050E
04DF
050D
053B
0524
0501
0519
0538
0508
04B7
04C4
052B
0540
04A7
040D
0468
0573
0578
0310
FEE9
FB5D
FA28
FADA
FBAE
FB98
FB17
FB11
FB82
FBA3
FB23
FA9C
FAB6
FB36
FB60
FAFB
FA99
FAB6
FB0F
FB1D
FAE3
FAD7
FB23
FB66
FB5B
FB54
FBA9
FBF5
FB7A
FA70
FA5C
FC9C
00A6
0441
05A3
050E
0437
0448
04F0
0542
0506
04D1
0504
0545
051A
04B0
04A2
0517
057D
0553
04DC
04B5
04EF
04F8
047F
0404
0424
04A7
04CF
048B
04A0
0558
0583
0397
FFC0
FC21
FAB0
FB34
FBDA
FB7F
FAB7
FA93
FB0F
FB4D
FAF2
FA8B
FAA1
FAFF
FB23
FB0B
FB1E
FB6E
FB8F
FB41
FAE9
FB0F
FB97
FBE0
FBA3
FB53
FB71
FBBC
FB84
FAC4
FAA2
FC66
FFED
0370
0523
04EB
0442
046B
0537
05A1
054F
04E7
0507
0564
0551
04CA
0476
04A8
04E8
04B9
045F
0472
04E9
051C
04BF
045A
047C
04D6
04B3
042B
0432
0526
05C0
0430
0051
FC35
FA2F
FA96
FBC0
FC0C
FB6B
FADD
FAE6
FB18
FAF4
FAB5
FADB
FB52
FB89
FB4A
FB09
FB30
FB86
FB90
FB5E
FB67
FBB4
FBAD
FB05
FA69
FABE
FBC3
FC2A
FB5D
FAA4
FBF3
FF95
039A
05BD
058E
047E
0411
0471
04D0
04B7
047A
0491
04E7
0509
04CF
048C
049C
04E8
0512
04EF
04BB
04B9
04CF
04C4
04A3
04AB
04CD
04B7
046C
047F
052D
0581
03F1
003D
FC40
FA45
FAA9
FBAC
FBAB
FAE9
FAB8
FB72
FC21
FBF5
FB5D
FB38
FB85
FB84
FAE9
FA5F
FA8A
FB21
FB6B
FB43
FB25
FB4D
FB64
FB20
FADA
FB14
FB9E
FBAF
FB00
FA91
FBDF
FF43
034A
05E6
0638
052C
0451
0459
04C3
04D4
0487
045F
0489
04AF
0496
0485
04CC
0537
054C
04FD
04C1
04DE
0507
04E0
049B
04A4
04E1
04BE
0436
041C
04F1
05B1
048E
010A
FCDB
FA55
FA21
FAE8
FB28
FACA
FABA
FB56
FBF5
FBE3
FB59
FB18
FB5D
FBA9
FB7F
FB0C
FAD0
FAE7
FAF8
FAD8
FAD4
FB32
FBAB
FBBC
FB6D
FB46
FB81
FB94
FB0D
FA9B
FBAF
FED5
02B6
053E
05A0
04F1
04B2
052C
0587
052A
047C
043C
0489
04DF
04DC
04A8
0498
04AE
04AE
0493
04A1
04F2
0538
0524
04D3
04A4
04A5
047F
0413
03E5
047A
053E
04A2
01B9
FDA2
FAB8
FA3B
FB2D
FBB5
FB35
FA91
FAA4
FB27
FB5A
FB2E
FB35
FB92
FBB6
FB4F
FAE6
FB16
FBA2
FBC4
FB53
FAF8
FB2E
FB90
FB83
FB2E
FB46
FBEB
FC46
FBAB
FAD3
FB68
FE37
0224
0515
05D8
050D
0448
046E
0511
0546
04DF
0480
04A9
050E
051D
04CE
049F
04CD
04F7
04C1
0470
0482
04E2
04FA
04A8
0479
04C3
0506
04B0
0426
0446
04E0
0469
01BD
FDD1
FAF4
FA66
FB30
FB98
FB26
FAB0
FAE1
FB5F
FB84
FB43
FB08
FB02
FAFF
FAE5
FAF5
FB55
FBB1
FB93
FB0E
FABB
FAF5
FB5F
FB62
FB02
FADB
FB46
FBBC
FB7F
FADA
FB4F
FE07
0231
0574
062F
0512
0423
047A
055E
0590
04EE
0462
0488
0500
0527
04F3
04D0
04DB
04D4
04AF
04BC
0523
057F
055E
04E6
04AA
04DC
0501
04B4
045A
04A4
0549
04D8
0232
FE17
FAC2
F9C6
FA9B
FB7B
FB64
FAE2
FAE3
FB59
FB7F
FB17
FAC5
FB0E
FB90
FB9C
FB38
FAFF
FB27
FB37
FAD1
FA5C
FA70
FAED
FB29
FAFA
FB02
FBA1
FC2D
FBC5
FAD6
FB10
FD9A
019C
04ED
0618
0588
04BB
049E
04EF
0506
04C7
049D
04C9
0502
04E4
0488
0468
04BC
0525
052D
04F6
04FC
0554
0586
054D
0505
0515
0537
04E0
043A
0417
049A
0475
0242
FE71
FB36
FA35
FAD6
FB55
FAF4
FA7C
FABB
FB61
FB9E
FB58
FB26
FB51
FB6D
FB1D
FABA
FAD1
FB4A
FB7D
FB24
FAAE
FAA0
FAE5
FB06
FAE1
FAD6
FB27
FB7D
FB57
FAF7
FB88
FDF6
01AB
04CA
05E5
054C
0489
04A4
0538
0558
04E5
0496
04CE
0519
04F7
04A8
04C4
053B
0563
04F7
0485
04AB
0531
0561
050F
04C4
04D8
04EB
049F
0463
04EB
05D1
057B
02BE
FE70
FAE4
F9C0
FA8F
FB88
FB85
FAE2
FA92
FADB
FB39
FB42
FB23
FB31
FB54
FB3D
FAF8
FAE8
FB28
FB4A
FAF9
FA9F
FAE3
FB9C
FBE0
FB49
FAA4
FAE1
FBA3
FBA4
FAA9
FA55
FC79
00C1
04B9
0645
0598
048B
0469
04F6
0551
0530
04E9
04C8
04BD
04A9
04A0
04C8
0506
051E
0500
04DF
04E5
04FB
04EE
04C1
04A7
04B6
04BB
0483
044B
0491
0540
053B
0350
FFB0
FC20
FA5D
FA75
FB13
FB2C
FAF6
FB16
FB78
FB76
FAF2
FA9D
FAF3
FB81
FB8D
FB21
FAE4
FB10
FB2E
FAEF
FAC0
FB29
FBDA
FBED
FB2B
FA80
FAD6
FBC9
FC15
FB5C
FAF4
FC88
0022
03DE
05C0
058B
04AC
047B
04F3
052F
04CA
044C
0457
04D4
052D
0517
04CA
049A
049C
04C0
0504
054A
0547
04D4
0446
0426
047C
04BE
049F
0489
04FB
0587
04FD
02AB
FF41
FC48
FACE
FAB7
FB2F
FB88
FB96
FB81
FB76
FB82
FB8E
FB7A
FB45
FB0E
FAEC
FADE
FAE3
FAF9
FB06
FAEC
FAD3
FB11
FBA1
FBFB
FBAC
FB19
FB14
FBB1
FBF1
FB29
FA6F
FBBC
FF7B
03A6
05D0
05A0
04B2
0466
0499
0496
0461
0487
0509
0546
0501
04B7
04C9
04D6
0471
0400
0448
0539
05E3
05A0
04D8
0466
048E
04E0
04F6
04D8
04B4
0498
049F
04E9
0521
045A
01F4
FE8F
FBBA
FA8E
FAD2
FB7B
FBC3
FB9E
FB57
FB1D
FAFC
FAF9
FB0E
FB27
FB3A
FB51
FB5C
FB32
FAD6
FA9A
FABC
FB07
FB19
FAF7
FB0E
FB82
FBD4
FB8B
FAFC
FAE4
FB49
FB4C
FA8A
FA30
FBEB
FFC7
03AF
0574
04FE
0415
0425
04F5
057F
056B
051F
04DD
0480
041E
043B
0506
05CE
05BB
04F3
046C
04A7
051C
0517
04B5
0491
04D9
052B
053B
0522
04FC
04BE
0495
04EA
058D
0536
02B0
FE99
FB40
FA50
FB20
FBCB
FB7D
FAFE
FB25
FBAD
FBCA
FB53
FAD1
FAA1
FAA9
FAD4
FB3D
FBB3
FBAC
FB0A
FA6F
FA71
FAD5
FB08
FB02
FB1B
FB3F
FAFE
FA76
FA70
FB2E
FBAF
FB0C
FA43
FB7B
FF37
0340
0517
04B5
0411
0463
0503
04FB
0493
04A8
052E
054A
04C4
0460
04AC
052C
0544
0525
0543
0563
04FC
044D
042F
04D5
056C
054B
04D9
04D4
0520
0523
0508
059A
0694
061E
02EB
FE44
FAFF
FA71
FB4B
FB9C
FB12
FABA
FB1E
FB8F
FB5E
FADC
FABF
FB0F
FB43
FB25
FAF8
FAF1
FAF6
FB01
FB36
FB87
FB94
FB31
FAC7
FAC3
FAEB
FAB6
FA3D
FA35
FAC5
FB08
FA63
F9E4
FB61
FF2C
034B
0572
055B
049C
0484
04E2
04F8
04C7
04D4
0524
0530
04CC
046A
0460
0471
044C
042D
047C
050D
0554
053F
0551
05B7
05EE
059F
0542
0557
0575
04EF
0431
0478
05CC
0623
0386
FEC6
FAFE
FA28
FB2B
FBBD
FB43
FADA
FB31
FB92
FB42
FAB7
FACE
FB70
FBBE
FB6E
FB23
FB4E
FB84
FB41
FAC4
FA8E
FA99
FA96
FAA9
FB15
FB82
FB45
FA81
FA2C
FAAB
FB0A
FA6C
F9CF
FB46
FF2B
033A
050C
04C4
045C
04DF
057E
0545
049A
0475
04E0
050E
04B2
0462
048C
04CD
04BF
04B6
051D
0599
057F
04E8
049C
04E4
0535
0521
0509
055A
05AC
0557
04C0
04FF
05FC
05D8
0309
FE93
FB3D
FA8B
FB61
FBC2
FB31
FAAB
FADD
FB3F
FB1C
FAB3
FABB
FB45
FBAD
FB87
FB1E
FAE5
FAEB
FAFA
FAF0
FAD7
FAC0
FAC5
FB06
FB60
FB59
FAB9
FA1F
FA6F
FB7F
FBF9
FB1D
FA2F
FB5F
FF1E
0342
0549
04FB
0438
046C
051C
052D
04A6
0476
04F2
056E
0554
04F0
04D6
04FE
04FB
04CA
04D3
051F
0537
04EC
04B2
04E7
0535
0520
04D4
04CA
04ED
04BD
0461
04AE
05A6
05A5
0304
FE84
FAFF
FA4F
FB5B
FBCD
FB07
FA60
FACE
FB8D
FB70
FAAC
FA6F
FB1C
FBCB
FBB2
FB26
FAE7
FB00
FB00
FAD7
FAD4
FAFE
FB13
FB10
FB32
FB6B
FB4C
FACE
FA9B
FB12
FB79
FAF2
FA39
FB5D
FF2B
03B1
0626
05EE
04DD
04BA
055A
0592
0511
0498
049F
04B9
047D
043E
0472
04DF
04FB
04C7
04B8
04EF
0511
04EE
04C8
04D5
04EA
04E5
0509
0586
05DD
056D
0490
0461
0506
04E6
026B
FE38
FACD
F9DF
FAAE
FB55
FB1C
FAD3
FB29
FBA8
FB8E
FB04
FACD
FB1F
FB71
FB62
FB35
FB48
FB7E
FB80
FB4D
FB26
FB13
FADE
FA8F
FA7A
FAB8
FAEF
FAED
FB02
FB65
FB9D
FB2B
FAC0
FBFF
FF82
0399
05CE
0584
046F
0448
04E2
0503
046C
041A
04A9
0567
0562
04C1
0467
0499
04C3
048E
046C
04C3
052D
0519
04BE
04C2
053B
0597
0579
0523
04D9
0484
042D
045A
0521
053C
030C
FED5
FB18
F9FD
FB03
FBF1
FBA1
FAE6
FADD
FB52
FB5F
FAEB
FAB1
FB06
FB60
FB4B
FB1D
FB3F
FB74
FB4F
FB00
FAFF
FB3F
FB4A
FB0B
FAEE
FB18
FB23
FADD
FAB9
FB14
FB60
FAF2
FA88
FBF4
FFB6
03CD
05B5
0537
044A
0474
0539
055D
04D0
048C
04FA
0565
052B
04AA
0490
04D3
04F0
04CC
04C7
04FB
0519
04F9
04DA
04E3
04D4
0482
0447
048B
04FF
04FA
048C
0496
054D
0553
0310
FED4
FAF3
F971
FA16
FB20
FB5F
FB20
FB1C
FB54
FB55
FB11
FAEB
FB0A
FB29
FB1E
FB1C
FB49
FB6B
FB3B
FAE4
FAD4
FB1C
FB60
FB63
FB51
FB59
FB5B
FB42
FB48
FB8D
FBA1
FB1D
FAAF
FBE2
FF50
036C
05CF
05C0
04C7
049D
053D
057D
04F9
0480
04BA
053E
0552
04FE
04D8
0503
0509
04B4
0466
0474
04A8
04C1
04EC
054A
0571
04FD
0455
043F
04B6
04E3
0468
040F
0477
04A2
02CF
FEF6
FB57
FA0B
FAB5
FB60
FB15
FA97
FAC0
FB3B
FB3B
FAC8
FA96
FAD6
FB05
FADE
FAD2
FB30
FB88
FB5B
FAF0
FAEB
FB53
FBA1
FB94
FB6C
FB4D
FB07
FAAA
FABC
FB6C
FBF6
FB96
FB03
FC12
FF6B
0356
057F
0571
04AD
048F
04F7
051C
04E1
04CE
051B
0563
055A
052E
0511
04E2
0497
0485
04D5
0514
04C2
042E
0419
049F
0505
04D2
0486
04C9
0548
0521
045A
040B
04A0
04BC
02A8
FEB7
FB48
FA3C
FB07
FBB6
FB59
FAB6
FABA
FB2D
FB41
FAD7
FA8B
FAB7
FB09
FB25
FB26
FB45
FB66
FB53
FB32
FB4E
FB85
FB61
FADC
FA8A
FACF
FB53
FB96
FBAA
FBDF
FBF8
FB73
FAC8
FB89
FEAE
02F3
05D0
0623
0535
04DD
055E
05A9
052E
0481
044F
047F
04A5
04C0
0507
0554
054A
0506
0509
055E
056B
04F3
0487
04AE
0504
04E4
0473
045A
04A2
04A3
0436
042A
04E1
0513
0304
FEF5
FB55
FA19
FAAF
FB3F
FB13
FAE8
FB3B
FB7F
FB2A
FAA0
FA90
FAE4
FB02
FAD8
FADF
FB21
FB03
FA5F
F9FE
FA78
FB35
FB49
FAD8
FAD1
FB74
FBFB
FBE0
FBA2
FBD3
FBFA
FB60
FAB2
FBBF
FF29
032A
056A
057B
04D6
04B8
04F8
04F6
04C1
04D1
0527
0557
054D
0563
05A0
058E
0508
04B5
0520
05D5
05E3
052C
0489
0498
0505
052A
04FC
04D5
04B2
0447
03D8
0426
0516
0516
02A8
FE6A
FADB
F9D2
FAB2
FB82
FB4C
FACE
FAED
FB68
FB6C
FAE1
FA79
FA97
FAD2
FAAC
FA51
FA44
FA9A
FAE8
FAED
FADB
FAEE
FB10
FB11
FAFC
FAEF
FAEB
FAFE
FB4F
FBC6
FBDB
FB4B
FAE6
FC1D
FF5E
033C
05A8
05FC
055C
0511
053C
054D
0524
0511
0525
0520
04F4
04E8
050C
0514
04E5
04E3
0551
05B3
0569
04BF
04AB
0558
05B9
0512
041F
0416
04E8
0573
0537
04EC
0505
0488
0231
FE7D
FB83
FA98
FAEA
FAEF
FA5E
FA0B
FA5E
FACF
FAE9
FAEA
FB30
FB8B
FB99
FB6D
FB62
FB6D
FB2C
FA9B
FA44
FA75
FAC8
FAD0
FACA
FB21
FB98
FB91
FB15
FADE
FB3D
FB89
FB20
FAAD
FBBD
FEDF
02B2
0537
05C2
054F
0519
0565
05A8
0578
04FC
04A6
04B2
04EA
04ED
049A
0436
042B
0494
051B
0553
052A
04F4
04F7
051C
051C
04E6
04AB
049D
04BA
04D2
04B7
046C
043C
048C
0555
05D3
04E8
0227
FE7B
FB89
FA4E
FA61
FAAB
FA9C
FA87
FAD4
FB48
FB5F
FB10
FAE0
FB23
FB7C
FB69
FAFC
FACB
FB12
FB5D
FB31
FAC7
FAB6
FB0D
FB3A
FAF4
FABB
FB21
FBDB
FC17
FBA4
FB3B
FB69
FBAA
FB2C
FA45
FA81
FCE8
00A0
03AC
04DD
04B2
0469
04B1
0551
05BD
05B4
055D
0506
04DE
04E0
04DF
04C6
04AF
04C1
04EF
0500
04E2
04C4
04CF
04EF
0507
0510
04F8
049C
041C
03F2
0468
0504
04FD
0452
0405
04BC
0578
045A
00E6
FCEC
FAB3
FAA6
FB4E
FB4B
FAB4
FA65
FAA8
FB00
FB01
FAD9
FADE
FB04
FB0F
FB04
FB1C
FB61
FB91
FB73
FB1D
FAD1
FACC
FB19
FB8D
FBE0
FBE7
FBAB
FB4D
FAF4
FAD4
FB24
FBC8
FC22
FBA3
FABF
FB03
FDA3
01D7
0541
0631
0547
0477
04C0
056A
056B
04DA
049A
0501
056F
0548
04C1
0476
048C
04A8
049F
04A6
04D9
04F1
04B1
0461
0474
04D5
04EB
0470
03F0
0425
04E7
053F
04AA
03EB
041B
04FF
04E5
0277
FE74
FB22
FA13
FAC1
FB7F
FB62
FADD
FAB5
FAF2
FB19
FB05
FB09
FB56
FBA5
FB9F
FB54
FB21
FB30
FB49
FB28
FAE1
FACF
FB24
FB9C
FBCD
FB9D
FB5C
FB60
FB94
FB9E
FB6E
FB63
FBB0
FBDE
FB78
FB1B
FC49
FFA1
03B0
0621
061E
0501
0492
0514
0576
0519
048B
047F
04C7
04CF
0494
0490
04DA
0504
04D3
0495
0498
04A9
047E
0453
049B
052E
0543
0485
03B1
03BA
0486
0513
04C7
0435
0451
052E
05A4
045D
012A
FD54
FAA3
F9F1
FA9D
FB4B
FB3A
FAC9
FABA
FB21
FB67
FB30
FADA
FADB
FB15
FB24
FB14
FB50
FBDC
FC1A
FB96
FAC6
FA8D
FB1E
FBC4
FBDB
FB9D
FB9F
FBE0
FBD8
FB5C
FAF1
FB03
FB35
FAF2
FA8C
FB41
FDE2
0199
0489
058C
052B
04C2
0501
0581
05A0
0554
0507
04FB
050C
04FE
04C7
047A
042F
0404
041C
0469
04A0
0487
044E
0458
04AB
04D3
0482
0414
0420
04B9
054B
054D
04E3
04A7
04F0
0550
04D9
02DC
FF93
FC33
FA2F
FA14
FB05
FB92
FB2C
FA83
FA6A
FACF
FB0C
FAF9
FB07
FB6E
FBB6
FB6D
FAEF
FAF7
FB8D
FBF1
FBB1
FB4B
FB62
FBCB
FBDB
FB72
FB24
FB49
FB82
FB5E
FB1F
FB50
FBCA
FBB8
FADC
FA5D
FBC5
FF3E
0327
0589
05D6
0519
04B4
050A
0570
0534
047A
0402
043C
04D1
0529
051B
04F4
04E7
04D0
048A
0451
0474
04D3
04F7
04BD
0486
049D
04C2
0497
0440
0430
046E
047D
042C
0414
04C5
059A
04F9
0206
FDE1
FAC7
F9F3
FAB5
FB7E
FB84
FB28
FB0C
FB3E
FB61
FB53
FB5A
FB9C
FBCC
FB89
FAF1
FA86
FA8D
FAC4
FAD5
FAD8
FB1B
FB96
FBE0
FBC8
FBA6
FBD8
FC19
FBDA
FB2E
FAE3
FB6A
FC0D
FBC3
FAC7
FAC0
FD08
0106
0490
05F9
057E
049F
0476
04E3
0534
051A
04D5
04B1
04A7
0484
0450
0457
04BD
0539
0565
053A
0510
0517
0510
04B8
0444
0431
0498
04FB
04ED
04A2
0492
04B4
048D
0419
040F
04D2
0562
0414
0083
FC5E
F9EA
F9D8
FAE4
FB75
FB36
FAE4
FB03
FB48
FB3D
FAFA
FAEC
FB23
FB3A
FAF7
FAA8
FAC4
FB44
FBA5
FB9A
FB65
FB65
FB79
FB3C
FABC
FA8F
FAFE
FB87
FB7D
FB07
FAF7
FB8C
FBF2
FB62
FA92
FB4B
FE59
026A
0542
05EE
054F
04C4
04CE
0511
0534
053F
054B
053F
0501
04BC
04AC
04D0
04F3
04F3
04DC
04C5
04B2
0499
0479
0463
047C
04CC
0519
0512
04BC
0485
04B8
0513
051A
04DF
04FD
057F
0535
02CE
FEB6
FB2B
FA05
FACC
FB80
FB09
FA2C
FA20
FAD8
FB4F
FB11
FAC3
FB09
FB95
FBA9
FB38
FAE4
FB0C
FB58
FB5B
FB32
FB39
FB6D
FB72
FB27
FAE5
FB02
FB4D
FB4E
FAF8
FAC5
FB06
FB60
FB39
FAAF
FACD
FCA0
0003
0386
059B
05E0
053D
04CE
04EC
0533
0536
04EF
049D
0469
045A
046F
04A6
04DB
04DE
04AC
0485
04A8
0504
0541
0532
0507
0505
0522
051B
04DE
04BD
04F5
053A
0500
0458
0415
04C1
057C
0488
013C
FD18
FA74
FA31
FB12
FB60
FACD
FA59
FAC0
FB98
FC0C
FBE5
FB86
FB3A
FAFE
FAD3
FAE0
FB1A
FB37
FB0D
FAD6
FAE5
FB1E
FB1A
FABA
FA6E
FAA9
FB47
FBB5
FB99
FB2F
FAFB
FB32
FB86
FB83
FB44
FBB3
FDC2
0133
046D
05D7
0560
046E
0445
04C8
0509
04B9
0476
04BA
0525
0529
04EB
04F7
054D
055C
04EA
0480
04AB
0532
056E
053C
0517
053D
0548
04E2
0470
048C
050E
0526
048D
040D
046F
0536
04D2
0250
FE8B
FB7B
FA67
FAE4
FB95
FB97
FB14
FAB6
FAD2
FB33
FB7A
FB88
FB68
FB20
FAB4
FA5C
FA61
FAC7
FB2B
FB3A
FB14
FB17
FB50
FB61
FB11
FAB0
FAB8
FB14
FB31
FAD1
FA88
FAFE
FBE7
FC31
FB6F
FACC
FC07
FF78
0366
059B
0586
048E
0452
0504
05A1
0578
04EB
04B3
04E9
051D
051C
0526
055F
057B
0532
04C2
04A9
04EC
050D
04CC
0484
049E
04E8
04DF
0485
046C
04DF
055F
0543
04B0
0484
0526
05B0
04AE
01B1
FDF1
FB3E
FA6B
FACE
FB2B
FAF9
FAA3
FAAF
FAFD
FB0C
FAC9
FAAC
FAFD
FB53
FB2E
FABC
FAA8
FB29
FB9F
FB6E
FAD9
FAA0
FAF1
FB3A
FB25
FB1C
FB79
FBC2
FB4F
FA73
FA4E
FB33
FBEB
FB38
F9C5
F9D9
FCD2
016A
04F3
05FF
0565
04CD
04E9
053A
052E
04E0
04C5
04FE
053C
0540
051B
04FE
04EC
04C5
048E
0478
04A1
04E1
04FB
04ED
04EF
0513
050F
04AB
043D
0463
0523
05AF
055C
04A9
04B5
05A3
05EB
03E2
FFC7
FBE0
FA3D
FAC8
FBBA
FBC3
FB2D
FAEB
FB2C
FB45
FACE
FA39
FA36
FACA
FB5B
FB7B
FB55
FB3E
FB3D
FB29
FB12
FB33
FB86
FBAD
FB6A
FAFD
FAD7
FB00
FB16
FAE5
FAC7
FB1B
FB99
FB87
FACC
FA73
FBD1
FF0B
02AF
04FB
055B
04B3
043C
045B
049C
0493
046F
0498
0503
0539
04F8
049A
049C
04F1
0512
04BC
045C
0477
04EC
0523
04EC
04C3
0504
0550
0511
0476
044C
04DC
0566
052B
0490
0487
04EC
0449
019B
FDE8
FB52
FAD1
FB5B
FB79
FAFB
FAC0
FB38
FBC9
FBCA
FB6B
FB45
FB6E
FB72
FB2D
FB04
FB44
FB9D
FB8D
FB24
FAEE
FB2E
FB76
FB3C
FAA7
FA6D
FAE7
FB89
FB8A
FAE6
FA70
FAC9
FB7D
FB92
FAEE
FAE2
FCDC
00A0
0430
05BB
0552
0488
048D
051E
054A
04D1
044B
043C
0476
0492
048B
049B
04C5
04D0
04BF
04D9
0532
0575
0553
04F9
04D4
04F2
04F3
04A9
046D
0499
04F4
04F9
049D
0469
04AD
04FD
04D1
0467
047D
0510
04DC
02A4
FED4
FB70
FA21
FAA8
FB72
FB6E
FAF1
FAD4
FB36
FB7D
FB4C
FAF4
FAF1
FB3A
FB5F
FB1E
FAAF
FA72
FA8E
FAE4
FB37
FB54
FB2D
FAF2
FAEF
FB34
FB71
FB5C
FB18
FB06
FB35
FB48
FB08
FACF
FB0E
FB87
FB6E
FA99
FA34
FBBE
FF54
033C
056F
0577
049B
045D
0505
05B8
05B0
0509
046E
0442
0467
04A2
04E7
0534
055C
052A
04BB
0479
04AA
051D
0565
0552
0511
04E0
04D7
04F4
0527
0545
0519
04BF
04A1
04F3
0540
04EA
0426
03F7
04CE
0569
03E3
FFFC
FBCC
F9C0
FA24
FB31
FB5B
FADC
FACD
FB6D
FBE3
FB95
FAF5
FAC8
FB1A
FB5C
FB46
FB17
FB0A
FAFE
FAD2
FAB5
FADB
FB19
FB17
FADF
FAD2
FB11
FB3D
FB06
FAB0
FAAF
FAF2
FAF8
FAAF
FAB8
FB7B
FC4C
FC1D
FB17
FAF2
FD3C
0163
0502
0639
055E
0441
0414
048F
04E1
04D9
04D3
04EC
04DA
0489
0463
04BC
054D
057D
0525
04B3
048E
04B0
04E3
051C
055A
0565
050E
0499
0495
051A
0590
0566
04D7
048F
04B2
04AB
0429
03CE
0454
0530
04AF
01DA
FDD5
FAF3
FA64
FB38
FBB6
FB47
FAAC
FAA7
FB06
FB27
FAF1
FACF
FAEB
FAFB
FAD0
FABF
FB18
FB91
FB96
FB1C
FABB
FADD
FB2F
FB27
FAD6
FAC9
FB21
FB60
FB2F
FAED
FB18
FB7B
FB7F
FB27
FB23
FBAE
FBFB
FB51
FA7B
FB58
FEA3
02CC
0573
05D1
051C
04CB
050B
052E
04F4
04CF
0507
053B
0500
048A
0467
04B6
0503
04F5
04B0
0488
048F
04A6
04CB
0509
0535
0509
0498
0463
04B9
0542
055C
04F3
0498
04B2
04E7
04B0
043B
044F
050D
0546
0387
FFD6
FC0A
FA18
FA48
FB34
FB79
FAFF
FA97
FAC0
FB2F
FB63
FB50
FB3F
FB4D
FB50
FB26
FAF2
FAE5
FB01
FB23
FB37
FB42
FB48
FB4C
FB61
FB90
FBB3
FB89
FB1B
FACF
FAF8
FB59
FB67
FB07
FAC8
FB1A
FB90
FB63
FABE
FB0B
FD85
0191
0505
0638
0583
0486
0454
04A9
04D0
04B6
04C2
050A
0532
0511
04F7
0520
054A
0515
04A2
046A
048C
04AA
0484
0462
049B
0502
051A
04DD
04BF
04F3
050E
04BD
0467
04A1
052C
0526
045E
03D9
0471
0548
0461
00FC
FCC8
FA41
FA2A
FB25
FB96
FB45
FAEF
FAF8
FB13
FB10
FB35
FBA9
FBF6
FB9E
FAE5
FA8A
FAD5
FB42
FB4B
FB11
FB02
FB1C
FB08
FAC5
FAC9
FB41
FBA4
FB63
FACB
FAB5
FB52
FBD6
FB95
FB03
FB18
FBD4
FC1C
FB5D
FAC8
FC3C
FFF7
03F2
05DE
0570
045E
043E
04FC
0575
0518
0471
0439
0478
04BA
04C4
04BA
04BE
04C2
04C4
04ED
053E
0560
0510
048D
0463
04B6
0510
050A
04D9
04EB
052E
0522
04B2
0474
04CF
053B
04EF
041D
03EC
04CA
0554
039F
FF9D
FB92
F9D8
FA87
FBBB
FBEA
FB45
FADA
FAFB
FB21
FAF4
FAD2
FB1B
FB84
FB87
FB28
FAE8
FB08
FB42
FB48
FB2C
FB1F
FB0E
FADA
FAB8
FB01
FB89
FBB3
FB3D
FAB8
FACA
FB46
FB70
FB18
FAE4
FB3A
FB79
FAE2
FA13
FADC
FE27
0283
055E
05A1
048E
040B
0494
053B
0531
04BD
0490
04CA
0507
050B
0503
050A
04F6
04B6
048E
04C2
0521
0538
04EF
04A8
04B0
04DF
04E5
04CE
04D6
04EA
04B2
0439
041C
04C5
05A4
05B5
04D2
0416
0476
053F
0489
0167
FD36
FA60
F9F4
FADF
FB73
FB38
FAEE
FB26
FB81
FB6A
FAFD
FADD
FB40
FBAB
FBA5
FB47
FAF5
FAD1
FAC0
FAD1
FB30
FBB0
FBC3
FB3A
FAAF
FAE3
FBB8
FC45
FBF8
FB41
FAE0
FAEE
FAF7
FAE5
FB19
FB94
FB99
FACB
FA4D
FBF1
FFFA
044B
065A
05C2
0460
0408
04B9
053C
04F4
0471
045A
048F
049E
048E
04BF
052E
055F
050D
048F
0463
0494
04CB
04D7
04C7
04A3
045C
041A
043B
04D4
055B
0542
04B2
045F
048D
04AD
043F
03B7
03FA
04EA
0502
02DF
FEFC
FB76
FA04
FA71
FB3F
FB6B
FB35
FB4C
FBBC
FBF1
FB95
FAFE
FAB5
FAD8
FB1B
FB40
FB45
FB37
FB0A
FAC1
FA98
FACF
FB53
FBC1
FBC8
FB7E
FB3C
FB44
FB9D
FC16
FC5F
FC33
FB9E
FB20
FB45
FBE7
FC23
FB62
FA6E
FB0B
FE22
0277
059B
063A
052E
0446
0453
04CB
04F8
04EA
050B
054F
0542
04D9
049E
04EF
056F
0583
0522
04CB
04CC
04E4
04BE
046A
0431
041E
040A
03FC
042F
0496
04C8
0490
044B
046B
04C2
04BB
0453
0440
04D9
0523
03A5
0035
FC88
FA90
FA92
FB34
FB3C
FABF
FA8A
FADF
FB45
FB53
FB2F
FB1B
FB09
FACF
FAA1
FAD5
FB50
FB8B
FB45
FAE7
FAFC
FB73
FBBC
FB91
FB3D
FB1F
FB2A
FB28
FB34
FB8F
FC0A
FC15
FB90
FB23
FB6C
FBFD
FBD1
FADC
FAA0
FCAF
00B7
048B
063B
05D5
04DD
0475
0484
0483
047C
04CD
0565
05B0
0563
04E5
04C2
04FB
0526
050A
04DA
04C1
04A0
045A
0424
0444
0498
04B7
0481
0456
0484
04D5
04DD
04A4
0497
04CF
04D5
045D
03ED
0446
0513
04C4
022C
FE15
FAC3
F9C5
FA8E
FB63
FB49
FABB
FA9A
FAF7
FB44
FB37
FB1B
FB33
FB50
FB28
FADF
FAE0
FB42
FBA5
FBB2
FB79
FB3E
FB16
FAF6
FAF4
FB32
FB88
FB93
FB42
FB03
FB37
FBA2
FBBC
FB83
FB81
FBE4
FC06
FB5F
FAB6
FBB5
FF01
031D
05BF
0612
0543
04DE
052C
0565
0515
04B1
04C6
0531
0565
0532
04E4
04B5
0495
0474
0476
04AA
04D3
04B7
047F
0488
04D5
0501
04D6
04A3
04C1
04FF
04E4
046F
0435
0481
04D0
0481
03E2
03F7
04FC
0593
03F6
000D
FBD7
F993
F9A9
FAA5
FB08
FAB1
FA74
FAC5
FB3B
FB54
FB2D
FB30
FB63
FB63
FB0A
FAB5
FAC3
FB0E
FB24
FAF3
FADB
FB1C
FB77
FB94
FB87
FBA2
FBD8
FBBA
FB2B
FAAF
FACA
FB4F
FBA5
FBA1
FBA0
FBBE
FB84
FAD5
FAC9
FCDA
00F0
04EA
0698
05E5
04A6
0465
04F8
0558
0535
0518
054F
0571
0525
04C3
04CF
0522
0527
04C3
0484
04C9
0535
053C
04E9
04B8
04CE
04D3
0498
0478
04BD
0511
04F0
0478
044D
049F
04DB
048A
0421
045A
04DF
0447
01B0
FE09
FB48
FA70
FAC8
FB03
FABF
FA8C
FAD9
FB55
FB6E
FB0F
FAA2
FA82
FAAA
FAE6
FB0C
FB07
FAD8
FAA5
FAB1
FB0B
FB66
FB6D
FB2A
FAFC
FB0F
FB26
FB02
FADD
FB24
FBBE
FC00
FB8C
FAF3
FB0E
FBBD
FBEB
FB0D
FA4B
FB84
FF22
0353
05C6
05EA
051A
04C4
0501
0519
04D6
04B8
0506
0559
053E
04EA
04E5
0534
0550
04F6
0492
04A9
051D
0568
054F
0515
04FD
04F5
04DC
04CA
04E4
0507
04F8
04C8
04BF
04D5
04A9
0428
03D9
0431
04CC
04DB
0454
041F
04B6
0510
0383
FFDF
FC06
FA1B
FA65
FB5D
FB98
FB1A
FABD
FADF
FB10
FAE5
FA8A
FA6F
FAA8
FAF1
FB11
FB09
FAF1
FADB
FADB
FAFA
FB19
FB09
FAD7
FAD3
FB28
FB91
FB9C
FB43
FAF7
FB05
FB3D
FB43
FB20
FB26
FB59
FB62
FB2B
FB32
FBD3
FC82
FC3D
FB11
FAA0
FCA0
00CD
04D5
068A
05E3
04A2
0445
04BF
0526
0511
04D8
04D5
04EB
04E2
04DA
050C
0560
0575
052F
04D8
04B9
04C4
04CA
04C8
04D9
04E9
04C9
0482
0466
049E
04EE
04FE
04C5
047C
043E
03FC
03D8
041A
04B3
0511
04CB
0452
0471
0509
04BC
025E
FE82
FB31
F9F8
FA84
FB59
FB77
FB0C
FAB4
FAA8
FAC3
FAEA
FB21
FB52
FB54
FB2F
FB24
FB4C
FB70
FB5A
FB22
FB05
FB0C
FB0B
FAF7
FAED
FAFA
FAFA
FAE2
FAE1
FB20
FB6F
FB7E
FB5E
FB76
FBE1
FC21
FBC8
FB30
FB1C
FB9D
FBD5
FB2A
FA72
FB5A
FE7C
0272
051E
05AC
0512
04AC
04D6
0506
04E1
04AA
04BC
04F1
04E0
0480
0437
0451
049F
04C8
04C0
04C1
04EB
051B
0525
0517
0512
051B
0514
04F5
04D2
04B9
04AA
04A8
04BE
04CE
0498
0418
03B6
03DC
0451
046E
040D
03E3
048D
0551
0487
0175
FD7E
FAE2
FA7C
FB24
FB5D
FAFE
FAE1
FB60
FBDD
FBC2
FB5D
FB55
FBA9
FBBC
FB44
FAB3
FA8A
FAB5
FAD8
FAE8
FB16
FB4F
FB40
FAE3
FAA8
FAE4
FB5F
FBA6
FBA9
FBA6
FBA3
FB6A
FB18
FB30
FBD0
FC48
FBE7
FB0A
FAB7
FB32
FB8F
FB1E
FAC4
FC35
FFC1
0395
0594
0574
04A5
0465
049B
049D
0457
0441
0484
04BF
04B1
04A2
04E3
053F
053B
04D3
0484
04A9
0512
0552
0541
0501
04B6
046C
0439
043B
046A
0490
0494
049E
04CF
04F4
04CA
0475
0469
04BD
04F5
04AA
0441
0480
0556
056E
036E
FF9C
FBE1
FA06
FA22
FAE0
FB23
FAFB
FB04
FB60
FB97
FB5C
FAFA
FADF
FB08
FB1D
FAFB
FADE
FAF2
FB10
FB01
FADD
FAE8
FB2A
FB61
FB58
FB29
FB16
FB33
FB5E
FB6E
FB50
FB09
FABE
FAB4
FB0B
FB7C
FB94
FB54
FB44
FBAD
FBFC
FB6B
FA62
FA91
FD3D
0185
04F7
05F6
052D
0475
04B0
0547
0562
050E
04E0
0500
0516
04F2
04D4
04F4
051E
050D
04D8
04C2
04C7
04AC
0477
0475
04CB
0530
0551
053A
0524
0510
04D6
0493
049D
04ED
0506
04A2
0442
047E
050E
0503
042F
03AE
047C
05C2
0557
022A
FDBB
FAAA
FA16
FADE
FB57
FB18
FAD7
FB06
FB41
FB11
FAA8
FA8E
FADD
FB31
FB40
FB2C
FB2F
FB3F
FB36
FB1C
FB13
FB19
FB08
FAE4
FAE0
FB0D
FB34
FB23
FAFF
FB08
FB33
FB39
FB14
FB19
FB70
FBB2
FB72
FAF8
FB05
FBAF
FC09
FB5F
FA96
FB8D
FEED
0308
056B
0567
0487
0481
0559
05E2
0584
04E9
04D8
0527
052A
04BD
046C
0497
04F3
0515
0504
0505
051D
051A
04F6
04E1
04DF
04BC
047A
0476
04E5
0569
0571
0502
04A7
04A1
0495
0447
041B
047B
0503
04EA
0447
042F
0519
05AE
03FA
FFE4
FBBB
F9E2
FA6B
FB71
FB7F
FAE3
FAAA
FB08
FB54
FB28
FADE
FAE2
FB0E
FB02
FACA
FAC4
FB0B
FB5C
FB7E
FB84
FB7F
FB54
FAF6
FAAA
FAB9
FB0B
FB3F
FB34
FB2C
FB50
FB63
FB33
FB06
FB40
FBB6
FBC7
FB4D
FAF8
FB69
FC1D
FBF1
FACF
FA4F
FC2A
0020
03FE
05CA
0598
04F9
0504
056B
0566
04EE
04A2
04CF
0514
0504
04C4
04B9
04EA
0501
04D4
04A7
04BF
0500
051E
0508
04EA
04E0
04D9
04CB
04C9
04D3
04C5
0491
0471
049A
04D5
04C2
0475
046E
04D4
0515
04B3
0431
0484
057F
056C
02D7
FE8D
FB17
FA25
FAF4
FB93
FB3A
FAB6
FAD9
FB51
FB50
FAD0
FA7E
FAB3
FB04
FAFF
FAD2
FADD
FB11
FB15
FAEA
FAE9
FB27
FB4E
FB2A
FB03
FB2D
FB7A
FB7D
FB32
FB07
FB2A
FB47
FB24
FB15
FB69
FBC2
FB82
FADD
FAC6
FB90
FC31
FB8C
FA40
FA72
FD62
01BE
04EF
05BB
052C
04E3
0543
058E
0547
04D5
04C8
0511
0543
053B
052F
0539
052F
0500
04DB
04E7
04FB
04E4
04BE
04D4
0527
055E
0539
04E6
04B8
04BB
04BC
04B1
04BF
04DE
04BF
044B
03F9
0449
04FB
053B
04C2
0459
04CE
0580
04B1
0183
FD4D
FA74
FA00
FAD2
FB42
FAEF
FAA9
FAF8
FB6B
FB6B
FB19
FAFD
FB2A
FB35
FAF8
FACF
FAFE
FB32
FB02
FA96
FA73
FAB4
FAEF
FADD
FABF
FAE2
FB18
FB06
FAC9
FADB
FB53
FBAF
FB93
FB4F
FB57
FB80
FB5B
FB10
FB44
FBF9
FC30
FB45
FA51
FB5B
FEED
031E
0575
0573
04A5
048B
0511
0549
04ED
0492
04A2
04D8
04D7
04C3
04F1
0546
0562
0536
0518
0534
0546
0517
04E1
0501
0561
058D
054D
04E9
04BA
04BB
04C0
04CD
04FC
051B
04DF
046C
0452
04C0
0513
049F
03C5
03AE
04B4
0574
0415
0070
FC81
FA72
FA8F
FB5F
FB88
FB19
FAEC
FB53
FBC1
FBAD
FB37
FADD
FAD2
FAE6
FAEB
FAEB
FAF2
FAE7
FAC0
FAA5
FAC2
FAFC
FB17
FB01
FAE5
FAE9
FAFC
FB0F
FB2F
FB65
FB7E
FB4A
FAF6
FAE4
FB1D
FB37
FAFF
FAE4
FB66
FC22
FC1D
FB34
FADC
FCC1
00B2
0478
0602
056C
047C
047A
0516
055A
050F
04C3
04CD
04E4
04BB
0486
049D
04F3
0530
0531
0516
04F6
04C8
04AA
04DA
054D
058A
0537
04A0
0465
04A6
04E3
04C0
0489
04AA
04FE
050B
04D1
04CA
0511
0511
0465
03B4
03F9
04EE
04D9
0268
FE6B
FB2D
FA1E
FA9D
FB1D
FAF2
FAA5
FACD
FB37
FB54
FB04
FAA4
FA7D
FA81
FA90
FAAE
FAE0
FB0C
FB1F
FB33
FB5F
FB81
FB62
FB13
FAEC
FB1F
FB75
FB92
FB6F
FB4A
FB45
FB3D
FB1D
FB13
FB3D
FB60
FB2A
FACB
FAD2
FB61
FBC4
FB4F
FA93
FB2E
FE0F
0227
053F
0621
059B
053B
058C
05DC
058A
04EA
04BB
0519
057D
058E
0587
05A9
05C0
0573
04DD
0475
0477
04A0
04A3
048C
0493
04BA
04D6
04DB
04E2
04E5
04B8
046E
0467
04D6
0562
058F
055B
0525
0504
04AD
0427
041B
04E6
058C
0459
00D9
FCC3
FA63
FA48
FB00
FB08
FA70
FA3E
FACC
FB54
FB19
FA65
FA0C
FA54
FACB
FAFE
FAF8
FAF7
FB02
FAFF
FAF8
FB0E
FB3C
FB5C
FB60
FB63
FB69
FB52
FB1A
FAFD
FB27
FB63
FB5D
FB1F
FB0A
FB44
FB75
FB46
FAE8
FADD
FB36
FB71
FB3D
FB03
FB53
FBF4
FC09
FB5C
FB21
FCD7
007F
0441
061D
05CB
04B7
0457
04D3
055C
055F
0513
04EF
050F
0533
052F
0512
04F7
04E5
04E3
0504
0545
0570
0554
04FA
04A0
046E
045E
0464
0484
04B1
04C3
04B2
04B0
04EB
0533
051F
04A1
043A
045D
04D4
04FF
04B4
046C
0483
04A8
046D
041F
0477
0551
053F
02F7
FEFD
FB73
FA06
FA72
FB33
FB4E
FAFB
FAD5
FAF5
FB15
FB1E
FB30
FB47
FB29
FAD3
FA98
FAB1
FAF2
FB10
FB10
FB22
FB3F
FB2F
FAF9
FAEF
FB35
FB7C
FB6B
FB29
FB2C
FB7F
FBA9
FB5E
FAFA
FB01
FB58
FB71
FB28
FAFE
FB55
FBC4
FBA9
FB20
FAF3
FB6C
FBCD
FB53
FA9C
FB4C
FE38
0239
052C
05F3
0545
048F
0486
04E2
0522
052F
052D
052C
0526
052B
054C
056A
0552
0509
04D7
04E9
051B
0528
050B
04F1
04EB
04D3
049D
047E
04A7
04EA
04F1
04BE
04B6
0500
053B
04FF
0480
045C
04C4
0529
0505
0496
047F
04CA
04E3
0492
0477
0507
056F
0425
00C8
FCEC
FA9F
FA63
FAFC
FB1B
FAB8
FA8C
FAD6
FB27
FB2C
FB13
FB15
FB11
FAD9
FAA5
FACD
FB36
FB60
FB14
FAB5
FAAE
FAE1
FAF1
FADF
FAFD
FB53
FB77
FB2A
FACB
FADB
FB42
FB72
FB39
FB05
FB35
FB7D
FB5F
FAFC
FAF5
FB7C
FBFE
FBEC
FB86
FB61
FB6A
FAFD
FA1F
FA1B
FC4B
0059
0437
060B
05D6
0507
04C4
0506
0537
052B
0523
053B
053A
0505
04D7
04E8
050E
04FF
04C6
04BC
0505
0557
055E
0525
04F3
04DD
04C0
049A
049F
04DE
050D
04E3
0490
048A
04E3
0525
04F5
0499
0499
04FF
0549
0525
04D7
04BF
04C1
0496
0477
04E0
057D
04F4
0242
FE3A
FB08
FA16
FAC1
FB5A
FB1A
FA9F
FAA7
FB0C
FB33
FB04
FAF1
FB25
FB49
FB1A
FADC
FAED
FB31
FB3A
FAF8
FAD0
FB00
FB43
FB48
FB31
FB4D
FB84
FB74
FB0F
FACC
FB01
FB5C
FB55
FAE7
FA9A
FABD
FB09
FB24
FB2C
FB63
FBA4
FB8C
FB2C
FB13
FB76
FBB9
FB4C
FAD5
FBD5
FEED
02CC
0553
05AD
04E3
0472
04C2
0531
053E
051E
0530
055E
054C
04F4
04B4
04C1
04EA
04EA
04D3
04E5
0527
0560
0566
054C
052E
0507
04D8
04D1
0516
056C
0561
04D9
0448
0432
0493
04F6
0511
0503
04F1
04BD
044E
03EB
03F9
0463
04AA
04A2
04C1
0548
0565
03C7
0047
FC8C
FA8F
FAAA
FB7F
FBAB
FB26
FACA
FAF1
FB20
FAE2
FA77
FA5C
FA98
FAD0
FAD9
FADE
FAF4
FAF5
FACC
FAB2
FAD6
FB03
FAE9
FAA0
FA9B
FB04
FB74
FB84
FB5E
FB70
FBBF
FBDE
FB9A
FB4E
FB68
FBC1
FBDF
FBA1
FB5D
FB4B
FB2E
FADA
FAA1
FAE1
FB4C
FB2F
FA9D
FAD8
FD16
00EC
046D
05FD
05C0
050E
04DA
04FF
04F8
04C3
04BF
0500
0530
0510
04D2
04C2
04E1
0501
051A
0546
0577
056A
0506
048E
0455
045B
0468
046B
048D
04D2
04F0
04B4
045B
0458
04BD
0523
052C
04F3
04CA
04C3
04B3
049B
04AF
04E6
04E2
047E
0441
04B8
0563
04C9
0205
FE11
FB14
FA4F
FB13
FBC8
FBAC
FB39
FB12
FB2C
FB23
FAF3
FAF7
FB45
FB87
FB77
FB44
FB3D
FB5F
FB6B
FB4F
FB37
FB35
FB22
FAEE
FAD2
FB00
FB4B
FB61
FB41
FB43
FB83
FBAC
FB70
FB0C
FAF3
FB2A
FB41
FB07
FADB
FB19
FB83
FB99
FB61
FB5F
FBB1
FBB4
FB07
FA8C
FBCC
FF26
0315
0587
05CF
04F9
045A
044F
0470
047D
04A3
04F8
0538
051E
04CB
0494
049C
04BF
04DB
04F3
0504
04F3
04C1
04A0
04B3
04D6
04CC
04A4
04AB
04FA
053E
0528
04D7
04B8
04E6
0506
04CC
046C
0456
0493
04BD
049C
047B
04AC
04FD
04FD
04BF
04D6
055A
0546
0363
FFD2
FC46
FA75
FA78
FB08
FB18
FACA
FAC3
FB14
FB43
FB16
FAE2
FAFE
FB45
FB61
FB53
FB59
FB7C
FB77
FB30
FAE9
FADC
FAEA
FADE
FAD6
FB0F
FB6F
FB91
FB5F
FB41
FB86
FBE2
FBCC
FB48
FAEB
FB06
FB39
FB0C
FAAF
FAAB
FB11
FB62
FB59
FB4B
FB86
FBAD
FB33
FA87
FB11
FDB6
0195
04AE
05CC
0574
04FC
050B
0547
0530
04D8
04A6
04C0
04EC
04F4
04E7
04E8
04F4
04F2
04E5
04E7
04F9
0506
0504
0501
04FF
04E7
04B3
0493
04BD
0514
0535
04EB
047C
0452
0472
048A
047B
0483
04CF
051B
0510
04D0
04C4
04F9
04F9
0497
0467
04EC
0575
0474
014E
FD64
FAD3
FA5D
FAF1
FB34
FAEB
FAB0
FACC
FAE8
FACB
FABB
FAFA
FB49
FB48
FB0F
FAFD
FB20
FB2E
FB09
FAFB
FB2F
FB5C
FB2E
FAD2
FAC4
FB1C
FB61
FB3D
FAFD
FB1A
FB7E
FBA9
FB6A
FB1E
FB15
FB1C
FAE6
FA9D
FABB
FB4A
FBBD
FBA9
FB68
FB8E
FBF5
FBD3
FAF7
FA8D
FC14
FF96
0352
0562
0585
0507
050E
0576
0579
04FE
04A9
04D6
0517
04EE
0499
04AB
0523
0567
052B
04DB
04F3
053E
0532
04D9
04CC
053E
0595
0551
04CA
04B2
050A
0531
04DF
048F
04B3
0506
0503
04BC
04BA
0508
0513
049D
0437
0468
04C2
048B
03FE
0413
04E6
04FF
02E5
FF14
FBC7
FAA0
FB18
FB86
FB24
FA91
FA8A
FAE4
FAFE
FABB
FA94
FADC
FB46
FB56
FB06
FAC0
FACC
FAF9
FAEF
FAB0
FA91
FAC2
FB10
FB2A
FB0B
FAFB
FB25
FB53
FB41
FB01
FAEE
FB27
FB68
FB6A
FB43
FB34
FB55
FB86
FBA6
FBA9
FB8C
FB64
FB5F
FB90
FB9F
FB26
FA7F
FAFF
FDAB
01BE
04FF
05EF
0541
04C2
0537
05D7
05BE
052C
04FA
054E
0582
052F
04BF
04BA
0501
051B
04F3
04DF
0507
0534
0532
050F
04ED
04CF
04B6
04BB
04DF
04F4
04D0
04A2
04B3
04F1
04F3
04A6
047A
04B9
0503
04D0
0450
0439
04BB
051B
04AA
03DF
03DF
04EB
05A6
0458
00D5
FCCD
FA4B
F9F7
FADF
FB9D
FB94
FB25
FAEF
FB0E
FB22
FAF0
FAAD
FAA7
FAD3
FAE3
FABB
FA99
FAB5
FAF2
FB04
FAE1
FACE
FAF5
FB34
FB5B
FB68
FB6E
FB6A
FB5C
FB60
FB7F
FB8F
FB67
FB2C
FB2A
FB5E
FB71
FB3E
FB1B
FB59
FBAF
FB92
FB24
FB18
FB90
FBB7
FB03
FA83
FC06
FFDD
0410
063A
05F0
04D6
048A
0515
0585
0564
050A
04D9
04C8
04B0
04A0
04B3
04DC
04FD
0515
052E
053E
0537
0525
0526
0531
051D
04E4
04BE
04CC
04E6
04D3
049B
046A
0458
0461
0486
04C1
04E8
04D8
04A1
0483
049B
04CA
04E8
04FA
050A
04FE
04C5
0493
049D
04AB
0457
03D4
03EC
04C0
050B
033F
FF7A
FBC1
FA09
FA59
FB28
FB4A
FAF1
FACF
FAF9
FB00
FAC5
FA97
FAAC
FADA
FAF0
FAF2
FAEE
FADC
FABB
FAAB
FAC5
FAF2
FB02
FAF3
FAEF
FB07
FB1A
FB0D
FAFC
FB0C
FB37
FB66
FB8A
FB8A
FB49
FAED
FAD4
FB28
FB8C
FB8B
FB29
FADE
FAF2
FB2E
FB4A
FB5B
FB95
FBC6
FB9E
FB52
FB73
FBEB
FBE7
FB2E
FB09
FD03
00DF
0479
05F3
058F
04F4
051C
058B
057A
0502
04BA
04C6
04D2
04BE
04C4
04FD
0536
054E
055E
0577
0571
0531
04EB
04E9
051A
0524
04E4
04A9
04BF
0500
0512
04DF
04A1
048B
04A0
04C9
04E5
04D6
049D
046B
0464
0478
0482
0486
04A2
04C6
04B2
0464
043D
047E
04C5
048B
041A
044A
0515
0504
02BB
FED8
FB94
FA7B
FB01
FB80
FB2B
FA8D
FA60
FAA0
FAE2
FB06
FB2B
FB40
FB21
FAEB
FAD7
FAE0
FADC
FAD4
FAF2
FB23
FB1E
FAD4
FA9A
FAB4
FAED
FAE8
FAB6
FACB
FB46
FBAE
FBA1
FB58
FB3C
FB4D
FB47
FB2D
FB3D
FB80
FBB2
FBB0
FB9E
FBA4
FBAC
FB9C
FB8F
FB9B
FB8B
FB32
FAE4
FB19
FB8A
FB5E
FA92
FAA0
FCF4
00FA
0470
05B0
0534
049E
04C6
0533
053D
04FA
04DA
04E6
04DD
04C6
04E1
052D
0562
054F
050B
04C5
04A2
04B7
04F3
051B
0500
04BD
049E
04B9
04D4
04BC
04A0
04C9
0517
051F
04D2
0497
04AA
04BD
0488
0446
0452
048D
04A2
049B
04CC
0528
052B
04AE
0446
0479
04DE
04B3
042E
0452
0524
04FA
026B
FE55
FB35
FA74
FB2D
FBB1
FB74
FB1F
FB29
FB3E
FB08
FACB
FAE3
FB23
FB1F
FAE2
FAC9
FAED
FB0D
FB0B
FB0D
FB32
FB64
FB85
FB91
FB8A
FB62
FB22
FAF7
FB05
FB30
FB3B
FB23
FB17
FB22
FB1D
FB0A
FB23
FB6B
FB8E
FB6E
FB5F
FB9F
FBD6
FB9A
FB27
FB1A
FB82
FBBC
FB71
FB37
FBA2
FC20
FBA2
FA84
FABB
FD8D
01B8
04AE
0554
04C3
0483
04DC
0521
0500
04D8
04F3
051B
0510
04F6
04FF
0506
04DA
04A0
0495
04A4
049B
048F
04B4
04EF
04F3
04B9
0495
04B9
04F2
04F1
04BE
0497
048A
046F
0442
0438
0459
046C
0462
047D
04CF
04FA
04C0
0478
0484
04AF
0482
041D
0425
04B5
050A
04A4
0439
04C0
059F
04DD
0195
FD72
FAF8
FAD3
FB86
FB93
FB00
FAA7
FAD4
FB12
FB10
FB06
FB2D
FB5C
FB58
FB37
FB24
FB12
FAEB
FADE
FB12
FB54
FB5B
FB38
FB30
FB44
FB36
FB01
FAEF
FB33
FB96
FBBE
FBAB
FB99
FB9E
FB91
FB72
FB74
FB93
FB7D
FB22
FAE5
FB08
FB3A
FB23
FAF9
FB25
FB88
FBA2
FB74
FB98
FC2D
FC4E
FB47
FA1F
FAF1
FE68
02A1
051E
0552
04AC
0481
04CD
04ED
04C8
04B8
04D8
04E4
04C5
04BE
04F7
0535
053D
052F
0534
052C
04F2
04B4
04AE
04C8
04C8
04BF
04E9
0535
0544
04EB
0475
0441
044A
044F
044D
0474
04B4
04BB
0488
0484
04D8
051F
04FD
04B9
04BF
04F1
04E3
049E
0499
04DA
04CC
0436
03E8
04A9
05A8
04ED
01B3
FDA5
FB25
FAD5
FB66
FB88
FB30
FAF8
FB07
FB05
FAD3
FAB6
FAD6
FAFD
FAF9
FAEF
FB0C
FB31
FB2D
FB12
FB10
FB20
FB27
FB33
FB5B
FB78
FB5A
FB1F
FB15
FB4D
FB7B
FB61
FB20
FAFE
FAFC
FAF0
FAEE
FB28
FB74
FB5F
FAE4
FA95
FACD
FB26
FB26
FB05
FB43
FBB9
FBC1
FB48
FB10
FB7B
FBBF
FB02
FA18
FB10
FEA6
02FE
058A
05B5
04FC
04C7
050D
051D
04E1
04CF
0501
0518
04E3
04B7
04D6
0501
04E3
0495
046E
0479
048C
049D
04C4
04EA
04E4
04C3
04C5
04F4
050E
04E6
04A9
049D
04C5
04F0
050B
052C
053C
0508
04A8
0486
04BB
04E1
04B8
0491
04C3
050C
04F2
0492
047A
04B9
04AE
041B
03D5
04A3
05A1
04C6
0164
FD51
FAFE
FADE
FB6E
FB62
FAE8
FABF
FAEE
FAEE
FAAB
FAA0
FB06
FB6E
FB6A
FB26
FB07
FB15
FB1C
FB23
FB4D
FB7B
FB6F
FB30
FB01
FAF8
FAEA
FAC7
FAC0
FAF9
FB47
FB65
FB5B
FB5F
FB75
FB70
FB58
FB6A
FB93
FB6B
FAEA
FAA3
FAFE
FB91
FBBA
FB86
FB81
FBBE
FBB7
FB3C
FAE9
FB2B
FB5B
FAB0
F9F3
FB1C
FED2
0320
0579
0571
04BE
04C5
053B
0542
04E6
04E1
055B
05AC
0565
04ED
04C8
04D9
04C5
04A3
04C1
050C
0531
0523
051E
0525
04FD
049C
0450
0455
0487
049F
0499
04AB
04DE
0502
0505
04FC
04D8
0473
0409
041A
04AA
050D
04D6
047B
0498
04FC
04FF
049E
048A
04FB
0535
04B7
0443
04CF
0594
0470
00AF
FC66
FA37
FA64
FB06
FAC2
FA24
FA37
FADA
FB21
FACB
FA84
FABC
FB0A
FAEF
FAA2
FA9B
FACF
FAEE
FB00
FB40
FB95
FBAE
FB91
FB8B
FBAA
FBA0
FB48
FAE9
FAD7
FB05
FB2C
FB3D
FB65
FBA3
FBC1
FBC2
FBDE
FC00
FBC6
FB33
FAE1
FB1F
FB68
FB36
FADD
FB06
FB8B
FB9F
FB23
FAF8
FB9A
FC20
FB8C
FAD0
FC22
0001
040F
05AC
04F9
0432
04A3
057A
058F
0522
0530
05CD
0612
058D
04E1
04B6
04D6
04B5
046C
0475
04CA
04FD
04E2
04BC
04AA
0489
0449
0421
0439
046E
0485
047D
047E
048E
0493
048E
0499
04A4
0484
0458
0477
04D0
04E7
049F
047D
04D2
0525
04F1
048C
04A6
0517
04FD
0437
03E3
04B4
0552
039A
FF88
FBB6
FA69
FB10
FB8D
FB0E
FA94
FAEA
FB73
FB4D
FAB7
FA8F
FAEF
FB23
FAE2
FAC5
FB3C
FBC6
FBC0
FB67
FB5C
FBA1
FBA9
FB53
FB13
FB2E
FB55
FB31
FAEC
FAEB
FB2F
FB5C
FB42
FB1A
FB23
FB54
FB8F
FBD6
FC19
FC19
FBCA
FB71
FB3E
FB0C
FAC9
FABC
FB13
FB75
FB79
FB52
FB7E
FBD7
FB8F
FA94
FA57
FC6B
0066
03EF
0542
04EB
049B
04F9
0559
052C
04C1
0491
048F
0481
047F
04C1
0517
051D
04D7
04BB
04EF
0514
04F0
04DB
0516
0545
04F6
046C
044C
04AA
04F3
04C4
0469
044F
0469
0464
043C
043F
0474
0484
0452
0438
0470
04AE
04A0
0474
0482
04B4
04BA
049E
04A5
04C3
04AE
0489
04E6
05BA
05B0
035C
FF2F
FB7A
FA20
FABB
FB77
FB4B
FAC0
FAA9
FAFD
FB1F
FAD5
FA7F
FA79
FAAC
FAC5
FAB1
FAAC
FAE8
FB50
FB9E
FB95
FB40
FAF8
FB0E
FB69
FB9A
FB72
FB35
FB2C
FB3D
FB31
FB21
FB4F
FBAF
FBEB
FBDE
FBCB
FBE9
FC04
FBC6
FB50
FB1F
FB53
FB8B
FB81
FB5D
FB49
FB1B
FAD2
FAEA
FBA8
FC4D
FBD1
FA8A
FA67
FCF2
0144
04C6
05E3
056E
0512
053A
0526
0489
041E
0488
0551
0594
0529
04BF
04D1
0514
0509
04BE
04AD
04FF
0558
055F
051F
04D8
04A7
0483
0469
0472
04A7
04E8
0503
04EE
04C9
04B9
04B6
04A2
0476
044A
0432
0433
044F
0485
04B9
04B8
0488
048D
0519
05A5
04DB
01EA
FDCE
FAC2
FA22
FB25
FBF0
FBAA
FB03
FAE3
FB33
FB43
FAF5
FAD7
FB2C
FB75
FB35
FAB2
FA8F
FAE9
FB43
FB4D
FB3F
FB5F
FB8B
FB73
FB18
FAD0
FAC9
FADF
FAF5
FB27
FB87
FBD5
FBC6
FB71
FB34
FB3C
FB5C
FB6B
FB7F
FBAF
FBCC
FBA3
FB64
FB78
FBDD
FBFC
FB7D
FB19
FC23
FF08
0287
04C6
051D
0489
045C
04DC
0553
0543
04F8
04F4
0526
051E
04C6
0485
049B
04C7
04C0
04A7
04C9
0510
0517
04C4
047A
048F
04D3
04E1
04B5
04A3
04C5
04CF
0495
0460
047C
04BD
04C3
048E
0480
04BA
04E8
04C1
0480
0483
04AD
0497
044E
045A
04CA
0495
0296
FF0E
FBC4
FA53
FAA9
FB69
FB8D
FB44
FB3C
FB8E
FBB8
FB76
FB21
FB26
FB65
FB71
FB38
FB1B
FB55
FB9E
FB93
FB47
FB28
FB60
FB9B
FB81
FB39
FB29
FB64
FB97
FB92
FB85
FB9B
FBAD
FB89
FB5B
FB73
FBC4
FBE3
FB9E
FB48
FB3E
FB69
FB80
FB90
FBD1
FBFA
FB77
FA8E
FAC1
FD4A
0164
04BD
05CC
0540
04D4
0539
05AD
0570
04DE
04BA
0504
051A
04C1
046B
047B
04B2
04A3
0456
0434
0460
0495
0495
047D
0484
04A0
04A9
04A8
04C0
04DF
04C4
046C
042D
044E
04A6
04D5
04BF
049F
049E
048F
043F
03E2
03DD
0430
0465
0443
043F
04CF
0558
0466
0145
FD2F
FA63
F9ED
FAC2
FB2C
FAC5
FA80
FB03
FBBA
FBC3
FB36
FAE7
FB2C
FB7F
FB66
FB26
FB44
FBA2
FBB2
FB54
FB07
FB1D
FB4B
FB3C
FB28
FB6D
FBD8
FBDE
FB77
FB34
FB6A
FBA8
FB65
FAD9
FAB6
FB25
FB93
FB9B
FB99
FBF7
FC5F
FC37
FBAA
FB7E
FBE5
FC0C
FB6E
FB05
FC85
002F
0420
061D
05D7
04E5
04B4
0528
054B
04D3
0466
0491
0510
0547
051C
04F2
0502
0512
04E4
04A6
04A3
04CD
04CE
048F
045C
0474
04B2
04D5
04E3
0509
0535
051A
04B4
046F
049E
04F8
04F1
0489
044D
0482
04C5
04AF
0477
048C
04C4
0492
0406
03FC
04C2
051C
0357
FF80
FBBE
FA1E
FA7B
FB0A
FAAB
F9F3
F9E7
FA84
FAFA
FAEB
FAD1
FB14
FB71
FB79
FB46
FB47
FB83
FB9B
FB67
FB35
FB3F
FB4D
FB17
FACC
FAD7
FB37
FB74
FB4E
FB23
FB5E
FBC6
FBC4
FB3F
FAD5
FB01
FB77
FB97
FB4F
FB24
FB57
FB8A
FB6A
FB42
FB85
FBED
FBB8
FB03
FB43
FDC4
01DD
053C
063A
0570
04AF
04D7
0547
052F
04C2
04B3
0513
054B
050F
04C8
04D8
04F9
04BF
045C
0463
04EB
0560
0553
0507
04F5
0513
04FB
04A7
048B
04D7
0515
04CA
0438
040C
0471
04D9
04CB
047F
0474
04B6
04E3
04CB
04AD
04B3
04A6
045E
0435
048A
04CF
03B8
00B1
FCE8
FA65
FA13
FAF6
FB79
FB18
FA8E
FA8C
FAE0
FAFC
FAD6
FAD8
FB27
FB62
FB40
FB07
FB18
FB5B
FB5F
FB0B
FAC7
FAEE
FB53
FB8B
FB78
FB51
FB2F
FAF3
FAA6
FA9A
FAFE
FB80
FBAB
FB76
FB43
FB56
FB94
FBD2
FC0B
FC3A
FC2B
FBCA
FB6B
FB74
FBAE
FB76
FAC8
FACB
FCBB
005E
03F6
05DE
05F9
0569
0528
0544
055A
054D
054C
055E
055A
0535
051B
0524
0527
04F8
04AA
0475
0471
0482
048F
04A0
04BA
04C8
04B4
049B
04AA
04D8
04E4
04B1
047E
0496
04EC
0527
0516
04E0
04BD
049F
0468
0442
047E
0500
0524
049A
0406
044D
0527
04FD
0297
FEB9
FB87
FA5E
FAA2
FAE0
FA8F
FA41
FA67
FAA6
FA92
FA6C
FAB3
FB41
FB74
FB26
FAE8
FB33
FBB3
FBCE
FB7D
FB45
FB59
FB5B
FB06
FAB2
FAD2
FB3A
FB5C
FB20
FAFB
FB31
FB67
FB3A
FAE1
FAE9
FB5B
FBAC
FB8A
FB52
FB73
FBB1
FB8B
FB1D
FB1D
FBB6
FC0E
FB60
FA68
FB02
FE13
0245
0537
05D9
0532
04DA
0539
0596
056E
0516
0509
0523
04F8
0499
0488
04EE
0548
051B
049D
046C
04AE
04F6
04F1
04D8
04F8
0531
052A
04EB
04D4
050E
054A
0544
0528
053E
0567
054B
04EE
04C0
04EB
0507
04B7
0449
043F
0480
0479
041A
0421
04F1
0582
0428
0099
FC9F
FA69
FA6B
FB42
FB80
FB06
FA95
FA9C
FADC
FB08
FB29
FB55
FB61
FB1F
FAC4
FABA
FB13
FB71
FB81
FB51
FB27
FB18
FB0D
FB06
FB18
FB3D
FB40
FB0E
FAD8
FAD2
FAD7
FAA1
FA3C
FA0C
FA4C
FAB6
FAEC
FB05
FB5A
FBE1
FC14
FBB1
FB35
FB3C
FB8D
FB59
FA97
FA99
FCBF
00A7
0438
05AA
0531
0469
046F
0505
0562
0543
04F8
04B9
047F
045D
048B
04FD
053E
04F7
046E
0437
047A
04E0
0521
0553
0592
05AA
0560
04E8
04B7
04E7
0512
04F5
04DA
0523
059D
05A7
0511
0468
043D
046D
0470
0437
0442
04C9
054E
054B
050C
0537
0593
04D3
020D
FE24
FB34
FA85
FB62
FC25
FBFE
FB61
FB08
FB0B
FB1D
FB2B
FB60
FBA5
FBAC
FB63
FB21
FB1E
FB1C
FACA
FA57
FA3C
FA91
FAE5
FAE2
FAC5
FAF0
FB4D
FB68
FB25
FAF7
FB2C
FB72
FB4D
FAD7
FA9F
FAE5
FB3F
FB39
FAF4
FAE0
FB17
FB55
FB7F
FBC3
FC13
FBEC
FB1B
FA83
FB99
FEC3
02A5
0540
05CD
0532
04BF
04DF
0514
04F3
04A7
048A
04A3
04C6
04EB
052A
0568
0560
0507
04BF
04E3
0554
059A
0581
0548
053F
0554
0545
050D
04E3
04D7
04B5
0466
0434
046E
04ED
053C
0528
04F8
04FC
0522
052D
0513
04F1
04B5
043A
03CB
03FB
04BF
04E9
032C
FFB0
FC3E
FA8E
FAAF
FB46
FB3C
FABE
FA8D
FAD3
FB0F
FAE2
FA7F
FA4C
FA62
FA97
FACC
FAFB
FB11
FAFA
FACB
FAC0
FAEC
FB1C
FB18
FAF4
FAF0
FB18
FB33
FB1E
FB01
FB17
FB59
FB83
FB73
FB4B
FB39
FB3D
FB3D
FB3F
FB5F
FB8D
FB90
FB5D
FB40
FB74
FBB4
FB8C
FB31
FBAD
FDDB
013A
0422
0554
0525
04ED
0573
063A
065D
05B4
04E0
047C
0497
04ED
0543
0573
055A
04F8
0497
0487
04BE
04E7
04D8
04C9
04F4
0530
052B
04E2
04A8
04AD
04C1
04A8
0473
0460
0473
047B
046A
0472
04AD
04E3
04DD
04BB
04BE
04D3
04A2
0435
0425
04C7
0557
0465
015F
FD78
FAB1
FA06
FABD
FB6D
FB68
FB07
FADA
FAF7
FB1A
FB1A
FB03
FAE5
FABD
FA9C
FAAA
FAEB
FB2B
FB39
FB27
FB30
FB60
FB85
FB7A
FB57
FB44
FB45
FB43
FB3D
FB43
FB4A
FB3F
FB3A
FB75
FBE9
FC23
FBC3
FB11
FABD
FAFA
FB33
FAF4
FAE2
FC43
FF6B
0304
0536
0577
04D6
0493
04D6
04FA
04AF
0464
048A
04F7
052B
0504
04D1
04D6
04F4
04F2
04D5
04CB
04DE
04F0
04EF
04E6
04D8
04BE
04A0
049E
04B3
04AD
0471
0442
0473
04E7
0515
04B5
042D
040C
0448
045C
0425
042D
04C1
050C
03AB
0059
FCA1
FA7A
FA6B
FB41
FB9C
FB3F
FAD8
FAD8
FB03
FB07
FB00
FB2B
FB6A
FB61
FB05
FAB7
FACD
FB31
FB8D
FBAF
FB9E
FB6C
FB29
FAFA
FB07
FB3B
FB45
FB03
FABA
FAC5
FB1B
FB5A
FB4C
FB21
FB19
FB29
FB31
FB51
FBB7
FC19
FBDF
FB20
FB12
FD06
00CA
0478
062C
05C3
04B5
045C
04C1
0519
04F7
04A9
0495
04B6
04D1
04D9
04E4
04E8
04C9
049E
04A4
04E4
050F
04E2
048A
046B
049C
04D2
04CC
04A6
04A4
04D7
050F
0526
0519
04EF
04B1
0482
048C
04B9
04AC
0448
040A
047C
0534
04CD
0248
FE60
FB23
FA05
FA99
FB52
FB46
FAD3
FAB5
FB04
FB4C
FB50
FB49
FB68
FB7B
FB46
FAF0
FAD4
FB02
FB31
FB2A
FB11
FB23
FB63
FBA0
FBB7
FBA6
FB71
FB1B
FAD1
FACF
FB1A
FB6B
FB83
FB72
FB68
FB60
FB40
FB2F
FB81
FC12
FC19
FB1D
F9FF
FA8E
FDAF
0220
057E
0679
05C7
04F9
04C8
04D5
04B7
049D
04DF
0551
056E
0512
049F
0476
048B
0499
0486
046C
0464
046E
0491
04D1
0502
04E4
0486
044E
0485
04EA
0504
04C2
0487
0494
04AB
047D
0439
0443
0486
0485
0435
0447
0528
05E6
04CD
0157
FD1D
FA6D
FA13
FAE3
FB51
FB0C
FAC3
FAEC
FB40
FB50
FB1A
FAD5
FA8D
FA44
FA38
FAAA
FB5E
FBB7
FB79
FB1B
FB25
FB7D
FB9F
FB63
FB2A
FB3C
FB5A
FB34
FAFC
FB26
FBAD
FBFE
FBC4
FB60
FB52
FB82
FB8A
FB75
FBB6
FC3C
FC34
FB33
FA55
FB71
FEF9
032B
05B8
0603
054E
04F4
0517
0524
04F9
04FC
0544
055B
04F9
047C
045E
0484
047F
0459
0495
0559
0605
05FA
0569
050F
0529
0539
04DC
046F
0486
050D
0563
0535
04DC
04B8
04B1
047F
043C
0430
043E
0409
03B4
03F0
04D6
0521
0345
FF5E
FB7E
F9B4
FA0F
FAF9
FB35
FAF9
FB04
FB54
FB52
FAD4
FA6B
FA84
FADE
FB05
FB08
FB3C
FB8D
FB7E
FAF4
FA82
FAB0
FB3C
FB76
FB2D
FAD7
FACD
FAD5
FA99
FA4B
FA64
FAE4
FB45
FB2F
FAF5
FB0F
FB7A
FBE1
FC27
FC62
FC58
FBA5
FAA2
FAB7
FD16
0126
04B8
0613
0586
04B6
04AA
050A
051D
04E9
04F1
0548
0573
052B
04C9
04B9
04E6
04F3
04DC
04EC
0524
0521
04AB
042D
043E
04E6
0594
05CE
05A3
055F
051E
04DA
04AE
04B5
04C6
0492
041B
03C8
03D3
03FF
0408
042D
04CB
0568
04B8
01F8
FE22
FB34
FA49
FAB2
FB05
FABA
FA5B
FA73
FAD0
FAFA
FAEC
FAF9
FB37
FB5F
FB4B
FB30
FB3E
FB50
FB2E
FAF8
FAFF
FB44
FB65
FB27
FAC9
FAAA
FACE
FAEE
FAEB
FAE3
FAE1
FAC4
FA96
FAAC
FB35
FBCC
FBE6
FB9E
FBA0
FC21
FC62
FBB8
FADB
FB87
FE8D
02A4
058E
0648
05B9
054A
055C
0564
0515
04C8
04DC
0522
0536
050F
04F1
04F9
0502
0502
0520
0555
0548
04C5
0426
03FE
0464
04DF
0505
04E8
04CA
04A9
046E
0452
04AB
054D
0587
0506
0459
043E
049A
04AB
043F
041E
04CB
054F
03F6
0064
FC60
FA1B
FA07
FACA
FB15
FAEF
FB07
FB6F
FB8A
FB0D
FA78
FA69
FAD2
FB2F
FB39
FB11
FADF
FAAC
FA92
FACA
FB48
FB9C
FB77
FB29
FB3C
FBAC
FBD9
FB6C
FADD
FAD6
FB47
FB89
FB53
FB1A
FB4D
FBA9
FBAC
FB70
FB7F
FBD8
FBBF
FAF3
FA9A
FC40
FFE8
03A5
0581
0560
04C1
04D0
0551
0577
0523
04DB
04E3
04EE
04BB
0492
04D3
0560
05B7
0595
0534
04DE
04A4
0481
048C
04CB
04FD
04E2
04A2
04A0
04EB
0522
0504
04D3
04E7
050A
04B7
03FB
038D
03E2
0476
0484
0433
046B
0550
0581
0379
FF83
FBC5
FA25
FA84
FB4B
FB61
FB07
FAF4
FB39
FB61
FB38
FB09
FB10
FB28
FB1A
FAFE
FB08
FB2B
FB2E
FB10
FB06
FB24
FB32
FB07
FAC9
FAB9
FACF
FADA
FADC
FB0F
FB73
FBB5
FBA8
FB98
FBE0
FC44
FC33
FBA1
FB3F
FB88
FBEE
FB8A
FA9D
FAC2
FD38
0141
04A0
05CC
0539
0476
046E
04D6
050F
04FD
04E9
04F2
04FC
04F7
04F2
04E6
04BB
048F
04B3
053B
05C0
05B9
051C
0463
0405
0412
0457
04AA
04DD
04BF
045E
042B
048D
053F
0579
04ED
0449
0460
04FE
051A
045B
03C1
0456
0573
0511
0211
FDB9
FA87
F9BC
FA7A
FB35
FB5C
FB5D
FB89
FB9C
FB58
FB05
FAFC
FB1F
FB06
FAA9
FA78
FAB7
FB23
FB55
FB49
FB47
FB67
FB7B
FB6B
FB62
FB86
FBB7
FBC1
FBA7
FB8B
FB67
FB20
FAE1
FAFA
FB61
FB87
FB1E
FAAF
FB03
FBF1
FC46
FB58
FA4C
FB2F
FEA2
02E5
0588
05CD
04FC
0496
04CB
04DE
0480
0436
047E
050F
0548
04FE
049C
0483
04AA
04D2
04DA
04CD
04B9
04AC
04B9
04DC
04EC
04CA
0498
0496
04BA
04B6
046B
042C
0446
047F
045C
03EB
03DC
048C
0552
0540
0473
041C
04DA
0580
0425
006C
FC42
FA02
FA2F
FB4E
FBCB
FB7B
FB32
FB67
FBBB
FBB0
FB4D
FAF8
FAE6
FB05
FB36
FB6A
FB82
FB55
FAF5
FAB2
FAC7
FB13
FB4F
FB62
FB69
FB6E
FB5C
FB38
FB35
FB6B
FBA7
FBB2
FBAA
FBDB
FC3A
FC55
FBEB
FB63
FB49
FB86
FB79
FAFA
FAF4
FC8B
FFBC
0321
0536
05A3
052D
04B2
0480
0482
04A9
04EB
0518
0506
04D7
04D7
050C
0523
04E0
047C
045D
048F
04BF
04B7
049E
04AB
04CB
04BE
047E
0447
0443
0463
048F
04CA
0505
04FF
0499
0427
0422
0476
0489
0415
03C0
0450
0559
0538
02C5
FED3
FB87
FA40
FA7F
FAE3
FAD6
FACA
FB27
FB96
FB8C
FB1B
FAD0
FAE7
FB19
FB25
FB39
FB8A
FBDA
FBBF
FB42
FAF3
FB32
FBB6
FBF3
FBC7
FB88
FB71
FB62
FB2F
FAFB
FB03
FB40
FB79
FB90
FB92
FB76
FB23
FACA
FAE0
FB7B
FBEC
FB80
FABE
FB4A
FE31
0266
0583
062D
0548
04B6
052E
05CB
058C
04A8
041D
045A
04E2
0516
04F3
04CD
04BC
049A
046D
046F
04A5
04BE
048A
0446
044F
049D
04D1
04C0
0496
0478
0446
03F6
03E5
046B
0536
0585
0529
04D8
0521
0543
03BC
0032
FC46
FA1F
FA3D
FB33
FB7F
FB10
FACF
FB19
FB53
FAFC
FA74
FA75
FB0C
FB93
FBA4
FB85
FB98
FBC4
FBB0
FB64
FB3C
FB56
FB60
FB20
FAE2
FB02
FB5B
FB7B
FB4F
FB47
FB9A
FBDE
FBA8
FB49
FB68
FBF2
FC00
FB3B
FAD6
FC86
0061
0456
062D
05B4
0499
0458
04D7
0524
04F1
04C9
0506
054A
0525
04CA
04BB
0507
0535
0504
04BD
04B5
04C3
048E
042F
041D
047E
04E9
04FC
04D8
04D0
04E0
04C7
04A0
04DC
057B
05C1
0526
043E
0420
04C0
0483
0204
FDF6
FAB3
F9D1
FA9F
FB54
FB29
FACB
FAEC
FB3D
FB1A
FAAB
FAAE
FB47
FBAC
FB3B
FA69
FA34
FADD
FBAE
FBF5
FBC3
FB8A
FB6E
FB48
FB28
FB51
FBAD
FBBC
FB42
FAC0
FAC7
FB29
FB38
FAD6
FAAF
FB2A
FB9A
FB32
FA86
FB63
FEAE
02F8
05C0
0609
0519
04AD
050C
054A
04F4
04AB
0504
0596
0593
04F9
0490
04C2
0516
04FC
04A9
04B4
051C
053C
04C3
0430
0426
048F
04D6
04CA
04C9
0506
052A
04EC
04A6
04D9
054D
0544
04A7
045E
04FE
0581
041A
0069
FC59
FA40
FA7E
FB64
FB5C
FA82
F9FD
FA49
FAD1
FAFA
FAE8
FB09
FB52
FB5F
FB22
FAF9
FB1B
FB51
FB63
FB74
FBA9
FBB8
FB40
FA7D
FA2D
FA9C
FB32
FB38
FAD5
FAC5
FB37
FB7C
FB1B
FAA4
FAE8
FBA6
FBBA
FAE3
FA9E
FCA2
00AA
0467
05E0
055A
0498
04AC
051B
051B
04CF
04E6
0574
05CD
057C
04E6
04AC
04D9
0500
04EA
04CF
04D4
04CC
049E
048D
04D5
0532
052F
04E0
04DA
054A
0592
0520
0463
0459
052E
05DB
0587
04C6
04CB
057D
051F
0255
FE14
FAE0
FA2E
FB10
FBA4
FB3E
FAAC
FAB5
FB0F
FB10
FAC3
FAC0
FB2F
FB7F
FB42
FACA
FAB2
FAFF
FB2F
FB01
FACC
FAF3
FB53
FB80
FB59
FB21
FB0A
FB06
FB0F
FB41
FB8E
FB8D
FB07
FA7E
FAB8
FB9E
FC12
FB56
FA5E
FB22
FE6A
02AC
0581
05FD
0542
04DE
0525
055E
051F
04CF
04E6
0534
0533
04D6
0490
04AD
04F8
051C
0518
051F
0534
0529
04FA
04D7
04D2
04BF
0486
0462
0490
04E9
0504
04D2
04B2
04D8
04EA
048E
042D
0496
05B4
060E
041A
0011
FBFD
F9D7
F9C4
FA68
FAA1
FA83
FAAA
FB2B
FB86
FB71
FB35
FB2B
FB41
FB35
FB09
FAFC
FB17
FB1C
FAEB
FABF
FAD3
FB0B
FB23
FB1F
FB42
FB87
FB8F
FB2A
FAC6
FAEA
FB74
FBB0
FB5B
FB15
FB83
FC3E
FC3B
FB62
FB2B
FD21
00F4
0484
05FE
058C
04C5
04BD
052D
055A
0538
0545
05A1
05D1
0579
04DF
048C
049B
04BC
04C0
04C9
04ED
04FA
04C8
0491
04A8
04FF
052C
0504
04D8
04F2
051B
04ED
047F
0450
0487
04A7
044E
03F3
0449
04F1
0463
018F
FD65
FA36
F972
FA65
FB51
FB59
FAFE
FAF6
FB27
FB0D
FAA0
FA64
FAA0
FAFF
FB11
FAE5
FAE1
FB24
FB63
FB60
FB38
FB2A
FB41
FB59
FB68
FB78
FB7D
FB54
FB0D
FAEE
FB13
FB3C
FB2A
FB12
FB60
FBEE
FBF7
FB26
FA86
FBCB
FF65
03AE
0653
0693
05B1
0542
0582
0599
0519
0498
04C4
0564
05B8
057A
051D
0514
0543
0554
053D
052B
051D
04E9
049E
048A
04BB
04DB
04A3
0452
044E
0480
047D
0441
0456
04FF
059A
0563
04A5
0488
0565
05D4
03FF
FFE3
FBA9
F985
F99F
FA5E
FA81
FA3C
FA54
FAD2
FB0D
FAC7
FA83
FAB2
FB05
FAEE
FA7E
FA55
FAB2
FB23
FB35
FB13
FB26
FB5F
FB54
FAF8
FAC4
FB01
FB55
FB4E
FB1A
FB32
FB80
FB68
FAD1
FA87
FB18
FBCE
FB7E
FA6B
FA85
FD47
01BE
0546
063E
0570
04BB
04EF
0572
0598
058C
05B8
05F0
05AF
04F1
0459
0464
04D9
052B
0532
0535
0559
0563
051E
04BF
049A
04B3
04C3
04B2
04B3
04DE
04F8
04CC
049A
04C9
0536
053E
04B7
0466
0501
05CC
04F3
01A7
FD62
FA93
FA25
FAD3
FAF6
FA60
FA0A
FA6A
FAE4
FAD4
FA81
FA92
FB0B
FB5B
FB3B
FB08
FB1B
FB4F
FB57
FB41
FB4B
FB63
FB41
FAF0
FAE5
FB52
FBBA
FB93
FB0E
FAE3
FB48
FB97
FB41
FAA4
FA96
FB28
FB7A
FB03
FAAD
FC0E
FF79
034D
0583
05B1
0520
050F
0573
0594
054B
0527
0570
05B0
056A
04E5
04C6
0519
0547
0500
04AE
04BF
04FB
04E7
0495
0489
04DD
0511
04D4
0490
04C2
0527
0509
0465
0413
048D
0523
04F5
0451
0463
0553
058B
035C
FF2B
FB52
F9CA
FA51
FB1F
FB0F
FA8A
FA73
FADA
FB15
FAD9
FA93
FAB5
FB0D
FB1C
FADE
FAD2
FB37
FB98
FB65
FABF
FA56
FA8D
FB1A
FB86
FBB3
FBBD
FB9B
FB43
FAFC
FB1C
FB71
FB63
FAD5
FA8C
FB30
FC2A
FC3C
FB63
FB63
FDD5
01F6
0536
05F0
0503
0475
0506
05C2
05AB
050B
04CD
0525
0574
054D
0501
0501
0533
0535
04FF
04E6
0510
0531
04F9
0486
0434
0430
0459
0494
04DD
050C
04DF
0464
0423
0484
0525
0532
048A
0411
0488
0530
0443
0100
FCD9
FA2B
F9E2
FAD5
FB69
FB43
FB11
FB31
FB41
FAF1
FA9B
FAB8
FB14
FB17
FAAB
FA63
FAA4
FB17
FB33
FB08
FB0F
FB62
FB9E
FB82
FB53
FB5D
FB76
FB4E
FB15
FB49
FBE1
FC23
FBA3
FAFE
FB20
FBDD
FC06
FB23
FA8B
FC23
0007
0414
0604
05A6
04AA
0483
0510
0566
0536
04F7
0505
0522
0505
04E0
04FF
0541
0541
0500
04EA
052D
055E
0519
04A0
048B
04EA
0526
04D9
0468
046B
04D4
0506
04C7
0485
049B
04AF
044B
03C6
03F9
04D6
04E9
02CB
FEEF
FB74
FA0E
FA78
FB27
FB2B
FAD8
FAD2
FB0B
FB0F
FAD8
FACF
FB16
FB4D
FB23
FAD4
FAC8
FAFB
FB10
FAE5
FACB
FB01
FB55
FB72
FB4F
FB1F
FAF9
FAE0
FAFE
FB81
FC21
FC3A
FB9A
FAFA
FB35
FC0F
FC4F
FB58
FA53
FB2B
FE69
0278
0530
05D9
0573
053A
0566
056B
050C
04B6
04D2
0528
052A
04BB
044E
0451
04B0
0503
0514
0503
04F8
04EF
04D9
04C5
04BC
04A4
046A
0448
047C
04D5
04C9
043E
03D6
0425
04D4
0502
0481
0431
04B3
052C
03EC
007E
FC85
FA2F
FA16
FAFB
FB6D
FB23
FABD
FAB0
FAE0
FB09
FB27
FB50
FB68
FB42
FAEF
FABF
FAE4
FB3D
FB88
FBB2
FBCE
FBE1
FBCD
FB7F
FB26
FB15
FB55
FB85
FB4B
FAE0
FAD4
FB40
FB84
FB23
FAC0
FBBF
FEBF
02A4
0570
061C
0557
0490
0483
04E9
052F
0526
04FA
04E6
04F9
051B
0524
04FB
04B5
0487
0495
04D2
0505
04FF
04C4
0482
0461
0464
0468
0451
043B
045D
04B2
04D8
048B
042D
046D
052E
0520
02FE
FF21
FB7F
F9DD
FA3B
FB28
FB74
FB2F
FAFF
FB11
FB08
FAB8
FA6B
FA71
FAB3
FAE7
FAFC
FB1D
FB56
FB76
FB50
FB0D
FB08
FB51
FB8C
FB68
FB13
FB09
FB69
FBC1
FBA8
FB59
FB61
FBC1
FBBE
FB04
FA9D
FC27
FFD8
03CF
05D2
057F
0463
040F
0495
0511
0513
04FE
0530
056A
0547
04EA
04C3
04E9
0508
04FB
0500
053E
0566
051A
0483
0439
047F
04DA
04AC
0414
03DE
0472
052E
0520
044F
03D5
0479
055B
0498
0168
FD44
FA91
FA3E
FB13
FB65
FAF1
FAA8
FB12
FB96
FB71
FAD9
FAA2
FB0F
FB74
FB38
FAA3
FA72
FACF
FB30
FB2F
FB09
FB27
FB73
FB7C
FB34
FB0F
FB5E
FBC9
FBC2
FB53
FB1B
FB64
FBA2
FB38
FA99
FB32
FDE6
01D7
0500
0612
057C
04A6
046C
049C
04B9
04B7
04D1
04FB
04F1
04B6
04B0
0512
057A
056C
0505
04DF
052C
0559
04D8
0405
03D1
047F
0535
050F
0450
0406
048D
050B
04B1
03FE
0424
052A
0568
0347
FF46
FBAB
FA3C
FAA8
FB5E
FB6E
FB36
FB4D
FB95
FB87
FB1D
FAE2
FB24
FB7F
FB62
FAD9
FA7E
FAAF
FB1E
FB47
FB24
FB19
FB53
FB82
FB53
FAF8
FAED
FB45
FB86
FB57
FB0F
FB3C
FBBC
FBC5
FB11
FAA4
FBFB
FF56
0332
0598
05DD
04FC
0457
0469
04BF
04D0
04A2
048A
04A6
04CB
04D3
04D7
04FF
0534
0534
04EC
04A4
04A4
04D1
04D9
04B5
04B7
0503
0540
0514
04B1
0493
04BF
04B2
043B
0403
04A9
057B
04C9
01CA
FDCF
FB0F
FA76
FB0B
FB68
FB33
FAFC
FB1B
FB3F
FB0E
FAC4
FADC
FB55
FBA8
FB74
FAFD
FACD
FB08
FB4A
FB30
FAE0
FADA
FB40
FB8C
FB3F
FAAA
FA99
FB30
FBAD
FB78
FB0B
FB36
FBC8
FBAA
FAA2
FA48
FC71
00CA
04C1
062D
056C
0478
047E
04FF
0517
04C1
0491
04C0
04EE
04CD
0488
0479
04B0
04F6
051F
0523
0505
04D0
04A3
0495
049B
049F
049D
049C
04A1
04BC
04E9
04F4
04AA
0454
0491
056E
05C2
040D
0038
FC29
FA16
FA5D
FB61
FB93
FAFD
FAA1
FAE0
FB30
FB26
FB0F
FB56
FBC3
FBC2
FB37
FAA9
FA9B
FAEF
FB30
FB36
FB43
FB84
FBB6
FB89
FB1F
FAF4
FB3E
FB9C
FB8B
FB1F
FB03
FB7A
FBD3
FB49
FA78
FB2B
FE50
028C
0564
05C2
04D5
0465
04D7
053D
04F4
0478
048A
0514
056D
0549
04FA
04D8
04DC
04DA
04CD
04CB
04D4
04D3
04BA
049B
049E
04CF
0503
04FC
04B3
046E
0470
04A4
04B9
04AD
04DC
0541
04D3
0272
FE89
FB30
FA1B
FADD
FBA7
FB7C
FAFA
FB02
FB5C
FB3F
FAA0
FA4E
FAB1
FB30
FB28
FADC
FAFD
FB83
FBBC
FB51
FABC
FA9A
FAEA
FB3D
FB59
FB68
FB8E
FB9A
FB4D
FAD2
FAAD
FB1F
FBB8
FBBE
FB18
FAC4
FC28
FF93
0385
05DB
05D6
04B4
041F
0479
04F3
04F6
04D3
0501
0553
054F
0504
04F8
054A
0566
04E6
0448
044E
04ED
055A
051F
04AE
04AC
0507
0524
04CC
0477
0490
04C5
0484
03F6
0404
050B
05F0
04F1
0196
FD71
FAB8
FA3B
FAED
FB54
FB02
FA9A
FAA8
FB03
FB3B
FB39
FB2C
FB1F
FAFB
FACF
FACE
FB00
FB28
FB1C
FB03
FB1E
FB6A
FB9A
FB7B
FB36
FB1B
FB3C
FB5A
FB40
FB09
FB0D
FB6A
FBBF
FB85
FAEB
FB2A
FD77
0175
0517
067B
05B8
0494
046B
04EC
0506
048E
0462
0500
05C3
05D2
0546
04E6
04FD
051B
04E6
04A8
04C8
051D
052B
04E1
04AC
04C6
04D7
048E
0434
044C
04B9
04D1
0454
03F1
046C
055E
053D
02E1
FEF3
FB8B
FA45
FADC
FBAE
FB85
FAA5
FA23
FA7B
FB1D
FB45
FAF0
FAB7
FAE5
FB1F
FB02
FAC2
FAD0
FB27
FB43
FAEB
FA97
FAD1
FB6B
FBBA
FB81
FB3F
FB66
FBB3
FBA4
FB59
FB69
FBDC
FBE1
FB0B
FA6A
FBBF
FF5D
0373
05C8
05EA
053D
0517
056D
0574
04FB
049F
04C8
0518
0508
04B0
0494
04E0
0533
053A
0518
051A
0537
051F
04BE
0469
0476
04C7
04EF
04BD
047B
047F
04AA
0492
042D
040D
04A6
0564
04CA
01F0
FDC6
FA83
F99F
FA87
FB79
FB70
FAE8
FACF
FB39
FB73
FB1A
FA9D
FA91
FAE7
FB1E
FB06
FAEE
FB15
FB41
FB29
FAF5
FB0B
FB6B
FB9E
FB5A
FAF6
FAF8
FB52
FB7F
FB4E
FB35
FB90
FBE1
FB67
FA77
FAA9
FD3A
0162
04CF
05DE
0514
043E
0467
050E
0540
04E6
04AF
04F9
055B
054B
04DE
049D
04C5
0501
04ED
049E
0477
0499
04BB
049F
0477
0497
04E7
04FB
04B1
0476
04A8
04FB
04E1
046A
0462
0516
0572
03E0
003A
FC57
FA50
FA75
FB51
FB80
FB0A
FACD
FB18
FB64
FB40
FAF3
FB05
FB6E
FBA5
FB6B
FB1B
FB21
FB60
FB6C
FB31
FB13
FB5E
FBCD
FBD0
FB4F
FAD2
FAD6
FB33
FB6B
FB6C
FB93
FBE9
FBD2
FAF6
FA3D
FB47
FEA2
02CC
0576
05BE
04D6
0471
04F4
0579
0543
049A
0440
0471
04C8
04D8
04AD
0499
04B3
04C7
04A5
0469
044E
0464
048D
04AF
04D7
050A
051E
04E7
0486
045D
0490
04BA
047F
0432
047B
0521
04BE
0233
FE36
FAF6
F9F8
FAB3
FB75
FB61
FB07
FB2B
FB9B
FBA4
FB2C
FADB
FB26
FBB9
FBF2
FBB0
FB5A
FB43
FB4B
FB2B
FAED
FAE7
FB3E
FBA4
FBB4
FB72
FB36
FB31
FB38
FB30
FB52
FBD0
FC42
FBE4
FACC
FA70
FC67
0077
046B
062A
05B3
04B6
0483
04EA
050E
04B5
046C
0494
04E3
04DF
048B
0450
046F
04C3
0501
0504
04DC
04B8
04B8
04CF
04D6
04CD
04D2
04E5
04DD
04B3
0497
049D
048C
044C
043F
04C1
0532
0413
00B3
FC7F
F9F2
FA04
FB43
FBB7
FB1E
FAA8
FB0F
FBBA
FBD3
FB6D
FB39
FB6D
FB9D
FB77
FB39
FB2C
FB33
FB12
FAF1
FB18
FB65
FB6B
FB0F
FAB9
FACB
FB26
FB60
FB46
FB20
FB47
FBA2
FBA6
FB10
FA92
FB70
FE36
01E3
04A2
0572
04F5
0486
04B4
04FA
04DB
049F
04C2
0522
0530
04CD
046B
046A
04A6
04C7
04B6
04A0
049E
04A2
04AA
04D1
0514
0538
050E
04C0
04A2
04C2
04DD
04AD
044F
043E
04D9
05AE
0564
02EC
FEE3
FB65
FA20
FABF
FB94
FB8F
FB19
FB05
FB4B
FB4C
FAF2
FAD6
FB43
FBB3
FBA5
FB55
FB32
FB28
FAED
FAB4
FAEC
FB7A
FBBD
FB6B
FAF9
FAE8
FB21
FB44
FB53
FB7E
FB82
FB00
FA9D
FBD8
FF32
0319
055F
0581
04CD
048A
04BE
04D3
04B5
04B8
04DB
04C4
0479
0473
04D3
0511
04CC
0469
0474
04CB
04E9
04C5
04C6
04F9
04F6
049D
046B
04B9
0515
04D8
0445
0447
04F4
04E1
02A7
FEC3
FB56
FA05
FA87
FB5B
FB7C
FB14
FAD1
FAFD
FB55
FB7C
FB5B
FB16
FAE3
FAEA
FB2C
FB7F
FBA9
FB9C
FB7B
FB68
FB5A
FB40
FB26
FB21
FB23
FB14
FB0D
FB49
FBB5
FBC5
FB24
FA90
FB93
FED9
0306
05BD
05FB
04F8
047F
04F1
0557
050B
048E
049C
0511
0538
04E5
04A2
04C3
04EC
04BE
0471
046E
04A6
04BD
049A
0469
043C
041B
0436
04B0
0532
0530
04C3
04B7
0545
0529
02DA
FEBB
FB2E
FA0C
FABB
FB59
FB1A
FAB4
FACF
FB18
FB09
FAD5
FAEF
FB2E
FB19
FACF
FAF0
FB7D
FBAB
FB2B
FAC8
FB3D
FC06
FC2B
FBAE
FB62
FB80
FB5E
FABC
FA75
FB28
FBE7
FB64
FA4C
FB17
FEE7
039B
0608
0587
0446
0446
053B
05AB
0531
04B6
04E5
0550
0557
0511
04EB
04E9
04C9
049B
0499
04A7
0479
0430
0440
04B6
050D
04EE
04B3
04CD
04FC
04B7
0439
0466
0543
054B
02FB
FEE2
FB53
FA08
FA93
FB50
FB57
FB04
FAE2
FAE6
FACF
FAB9
FAE3
FB23
FB20
FAE6
FAD3
FAFE
FB18
FAF8
FAE9
FB2D
FB80
FB71
FB1C
FB01
FB33
FB2E
FABD
FA7A
FAEE
FB96
FB7D
FAEB
FB98
FEAC
02F8
05F1
0659
055B
04CE
051D
0567
0525
04CC
04DD
051E
0513
04C9
04AD
04CF
04DA
04C0
04DD
053E
0566
0505
048D
0498
0512
056C
056C
054E
051F
04A5
0415
0435
052A
0581
036E
FF2D
FB40
F9D2
FA86
FB5E
FB45
FACA
FAAB
FABD
FA8B
FA50
FA8F
FB1B
FB42
FAEF
FACD
FB2B
FB6E
FB1E
FAB4
FAD1
FB2A
FB00
FA72
FA62
FB14
FBAC
FB73
FAEE
FB09
FB8A
FB77
FAF6
FBAE
FE9B
026B
04D2
0525
04AF
04B4
0514
052B
050E
0543
05AC
0598
04ED
0474
04BA
053F
0541
04D8
04AD
04E7
0515
0509
0518
0564
0580
0518
0498
0492
04D2
04A5
0419
041B
04F0
0535
033B
FF47
FBAB
FA58
FAFA
FBBD
FB90
FAF6
FACC
FB0C
FB23
FAF3
FAE1
FB11
FB21
FAD9
FA98
FACB
FB40
FB67
FB1D
FAD2
FADD
FB0F
FB1A
FB07
FB05
FB0A
FAFA
FB03
FB57
FBAC
FB7A
FB0E
FBC2
FE8A
0271
053D
05C7
0510
04B4
04FB
0510
0499
0441
049D
0546
057B
0533
04F6
04F3
04D5
0485
046E
04B9
04F2
04CC
04A9
04EF
053E
050B
0498
04A6
0530
0558
04D0
0488
0531
058F
038F
FF2D
FB15
F9B6
FA96
FB64
FB08
FA6C
FA8E
FB0B
FB0D
FAB9
FAD6
FB68
FB9C
FB29
FACF
FB28
FBB6
FBB6
FB4E
FB2B
FB58
FB50
FAFC
FAE3
FB39
FB72
FB2B
FADF
FB21
FB78
FB00
FA2B
FADF
FE2E
029F
058E
05F9
0528
04BA
04EE
051D
050C
0517
0551
054C
04DF
048A
04AD
04F1
04D1
0475
0468
04B9
04EE
04C9
0498
0496
0485
0436
041A
04A9
0570
0575
04B2
0458
0508
056D
038B
FF64
FB66
F9DC
FA87
FB60
FB3F
FAD7
FB1C
FBBB
FBC1
FB23
FAC0
FB0A
FB77
FB63
FAF2
FAAE
FAB5
FAC0
FAC7
FB0C
FB82
FBBB
FB92
FB70
FB96
FBA9
FB55
FAF5
FB0B
FB4B
FB03
FA8A
FB75
FEBC
030D
05DA
060B
04FA
047D
04D4
050A
04B7
046C
0498
04DF
04C9
0484
0482
04C3
04F1
050B
0551
059A
0561
04B2
044E
049F
0503
04C9
044E
046C
0504
0510
044B
03DA
0491
0533
0393
FF7C
FB6F
F9E1
FA99
FB86
FB7D
FB1C
FB35
FB7F
FB57
FAE1
FAC6
FB13
FB32
FAF7
FAE6
FB35
FB53
FAE0
FA76
FAD7
FBB0
FBFE
FB81
FB02
FB14
FB4E
FB2B
FB05
FB72
FC03
FBB2
FAC7
FB34
FE49
02B5
05BA
061E
051C
0477
048E
04B4
04A0
04BA
0527
056A
0532
04DF
04DB
04FA
04EC
04E0
0523
0565
0516
0459
0402
0470
04FE
04F5
0498
04A1
0501
04F6
0472
046F
054C
0594
0372
FF2E
FB4A
F9E9
FAAF
FBA8
FBAA
FB2B
FAF4
FB03
FAF4
FADB
FB00
FB36
FB13
FAB3
FA9D
FAEE
FB1F
FAE0
FAAC
FB0F
FBB7
FBD3
FB4A
FAEB
FB3A
FBAB
FB8C
FB18
FB08
FB4C
FB24
FAA5
FB47
FE33
0270
0585
0617
0528
048A
04C6
0519
04F9
04B9
04BE
04E0
04D9
04CF
0506
054A
0535
04E7
04E8
0541
0551
04CC
0443
044C
04A2
04AD
0485
04B8
0534
0538
04A0
046B
0537
05BC
03E9
FFA9
FB81
F9DE
FA84
FB68
FB61
FB05
FB17
FB51
FB1E
FAB8
FABF
FB1B
FB20
FABA
FAA2
FB24
FB8A
FB39
FAB9
FADF
FB7A
FBA6
FB37
FAF2
FB44
FB8F
FB39
FABF
FAF5
FB8C
FB67
FAA1
FB11
FE11
026D
0578
05F2
0501
0468
049C
04FD
051D
0525
052C
0504
04BE
04CD
0544
0587
052A
04A7
04B2
0526
0541
04D0
0474
04A2
04F2
04D1
0478
0485
04E0
04D3
0451
0450
053C
05B5
03D6
FFAD
FB9B
F9E3
FA69
FB54
FB6A
FB12
FB1A
FB69
FB61
FAF9
FABD
FAE3
FB09
FAEC
FACD
FAF1
FB20
FAFD
FAB1
FABD
FB33
FB9B
FBA3
FB87
FB82
FB66
FB12
FAF1
FB62
FBE1
FB8E
FAB4
FB18
FE0E
0288
05D5
066C
054B
045F
045B
04A3
04BB
04DC
0529
0543
04EC
0493
04B7
0519
051A
04C7
04CC
054C
0589
0506
0456
0444
04A2
04B2
0469
0474
04FB
0537
04B7
0448
04BB
052C
039C
FFA3
FB7B
F9A5
FA35
FB33
FB44
FADC
FAEB
FB5E
FB7F
FB32
FAFF
FB1A
FB1C
FAD7
FABD
FB20
FB8F
FB7A
FB14
FAFC
FB4F
FB9B
FBA3
FB96
FB86
FB35
FAB5
FAA2
FB4B
FBEC
FB88
FAA3
FB2D
FE3F
027D
0565
05F3
054C
04EF
0516
0516
04B8
0478
04A9
0506
053A
054F
055C
0529
049C
0429
0455
04E8
0522
04BF
0450
045F
04AE
04AC
0467
0475
04F0
0539
04F4
04B3
0500
051A
0380
FFE7
FC0D
FA14
FA47
FB1B
FB30
FAAF
FA7D
FAC7
FAF4
FAC0
FAA4
FB06
FB90
FBAC
FB56
FB10
FB1D
FB41
FB42
FB40
FB61
FB75
FB4A
FB11
FB1C
FB60
FB84
FB68
FB3E
FB16
FACC
FA9C
FB74
FE0D
01BF
04C0
05E1
0592
0513
04FB
050E
0511
0527
055B
0561
050D
04B4
04BA
04F0
04DF
048E
0479
04C0
04E2
0491
0443
047A
04EE
04FD
04B1
04AC
0513
0544
04E8
04AD
0531
057E
03B8
FF98
FB5C
F98D
FA4C
FB86
FB95
FACF
FA6D
FAC6
FB2B
FB20
FAE7
FAE1
FAF7
FAF0
FAF2
FB33
FB83
FB81
FB42
FB3E
FB93
FBD1
FB98
FB2A
FB14
FB61
FB7A
FAEC
FA2D
FA61
FC56
FFBB
0341
0585
0602
0560
04C7
04D4
0539
055A
0516
04D5
04E6
051E
052B
0504
04E2
04DD
04D0
04A4
047D
0480
0498
04A0
04A3
04BC
04C6
0485
042F
0466
0547
05AE
0413
0054
FC52
FA4A
FA95
FB79
FB4C
FA45
F9D9
FAAB
FBBC
FBD7
FB0E
FA6C
FA87
FAF3
FB21
FB21
FB42
FB6A
FB49
FB01
FB0E
FB6E
FB7B
FAF2
FA8B
FB17
FC27
FC65
FB68
FA9C
FBE2
FF65
0345
0576
05A4
050D
04E6
0540
0578
0538
04D2
04C7
0526
057F
0563
04E5
0480
0488
04D8
0510
0505
04D5
04AB
0498
04AA
04E6
051B
04EE
0463
041F
049D
0523
0418
00D5
FCD0
FA58
FA3C
FB25
FB62
FAC5
FA62
FAC8
FB4E
FB28
FA90
FA51
FAA3
FB02
FB13
FB13
FB4A
FB7F
FB5B
FB08
FB0C
FB75
FBAF
FB56
FADE
FB0A
FBBC
FBF1
FB24
FA65
FB85
FF0E
0357
05F7
0608
04D8
0443
04C4
0567
0550
04CA
049D
04EF
053A
052C
050E
0529
0538
04D6
0439
0409
0475
04E9
04DC
048E
048C
04C8
04BA
0454
044B
0508
059C
046A
00FB
FCDD
FA46
FA03
FAF1
FB73
FB0A
FA6E
FA65
FAE4
FB55
FB5F
FB2A
FB00
FAE8
FAD0
FACC
FB01
FB4D
FB64
FB43
FB44
FB96
FBDE
FBAA
FB29
FB08
FB74
FBAF
FB17
FA71
FB7C
FEE4
0316
05A5
05B8
04B4
0468
051A
05B1
0567
04B4
0478
04CF
051D
0506
04D9
04F3
052C
051F
04CD
0494
04A1
04AA
0471
0432
0457
04C3
04DB
046B
041B
0493
053A
0474
016A
FD52
FA74
F9F0
FACF
FB64
FB20
FABD
FAE1
FB45
FB4F
FB02
FADB
FB08
FB38
FB32
FB1F
FB29
FB27
FAEF
FAC7
FB19
FBC3
FC14
FBA9
FB0B
FB06
FB94
FBD0
FB33
FA86
FB51
FE40
023C
053D
061D
0577
04CE
04E9
054E
0539
04B0
0469
04C1
053D
053D
04D8
04A5
04D6
04FC
04CB
0490
04A9
04DE
04C1
046B
045E
04A2
04A0
041A
03DD
04B5
05E1
055B
021A
FD98
FA7A
F9E7
FABB
FB39
FAF0
FAA7
FAF0
FB6D
FB7B
FB14
FAB5
FAAB
FAD1
FAEF
FB02
FB15
FB19
FB0E
FB1F
FB6D
FBC6
FBCA
FB68
FB14
FB47
FBD0
FBE2
FB16
FA40
FAF5
FDEE
020D
052F
0617
0566
04B0
04CB
0543
0553
04EE
04A2
04BC
04F6
04FE
04E8
04F8
0526
0529
04EC
04AF
04A5
04AA
0486
045A
0479
04D7
04F1
0487
042B
0491
0561
0519
0290
FE83
FB20
F9F3
FA83
FB2A
FB09
FAA0
FAB1
FB1F
FB4B
FB13
FAEC
FB17
FB42
FB1B
FAE3
FB07
FB68
FB86
FB47
FB2B
FB7A
FBC1
FB74
FADF
FAD1
FB73
FBE7
FB6C
FA9B
FB05
FD88
0145
0463
05BA
0599
051A
04F6
0518
0512
04C2
0477
0481
04CC
04FD
04ED
04D1
04DA
04F3
04E8
04C2
04AF
04B5
04AA
048C
0499
04DA
04E3
0460
03D5
042D
0545
0579
0336
FEFD
FB2C
F9B0
FA40
FB1C
FB2E
FADD
FAF1
FB62
FB93
FB5B
FB25
FB31
FB3F
FB13
FAEA
FB17
FB69
FB61
FAEC
FAA0
FAF8
FBA1
FBE2
FB93
FB4E
FB88
FBD7
FB82
FABC
FAD9
FD01
00C4
0445
05EA
05BC
0506
04CE
0507
0518
04D6
04A0
04B7
04E9
04EC
04CD
04CD
04E9
04E7
04BA
04AA
04E3
051A
04EF
0481
0453
048F
04BA
046B
040B
046E
0575
05A7
0389
FF75
FB9F
FA00
FA7C
FB53
FB3F
FAA2
FA90
FB33
FBAB
FB60
FAC9
FAB3
FB21
FB65
FB2F
FAF2
FB22
FB78
FB6F
FB13
FAF4
FB43
FB88
FB65
FB2C
FB5B
FBB0
FB6A
FA94
FA85
FC92
005A
03E6
0587
0552
04A7
0491
04F9
053C
0520
04F0
04E3
04D6
04A6
0485
04B9
0520
0546
04F5
0485
0478
04CA
04FA
04BE
0477
049D
0500
04FC
0487
0468
0512
0580
03FF
0040
FC24
FA03
FA46
FB3F
FB57
FAB7
FA8C
FB2F
FBC8
FB9D
FB08
FAD4
FB19
FB42
FB0B
FAE1
FB28
FB92
FB8F
FB2A
FAF3
FB2B
FB63
FB33
FAE0
FAF3
FB54
FB4B
FAA3
FA68
FC0D
FFB5
03AD
05EC
05F5
050F
04A8
04F1
0521
04C6
045A
047D
0513
056E
053A
04CE
0493
0482
0466
0458
0499
0504
0520
04CA
0487
04CA
053D
052A
0493
0461
0511
0597
0434
008B
FC6C
FA28
FA4B
FB53
FB9C
FB14
FAC5
FB2E
FB9C
FB49
FA7E
FA32
FABB
FB6C
FB8E
FB42
FB29
FB6A
FB8F
FB4E
FAFD
FB07
FB4B
FB5A
FB36
FB4A
FB9A
FB8E
FAE6
FA99
FC11
FF77
032B
0542
055D
04B9
0494
04F6
0526
04DE
0496
04BE
0525
0550
0524
04EB
04DB
04D2
04A8
0482
04A1
04F0
050A
04C2
0470
047B
04BD
04B1
0447
0425
04C3
055D
0460
012B
FD25
FA97
FA69
FB67
FBD0
FB3D
FA9D
FAAE
FB1B
FB31
FAEB
FAD2
FB12
FB45
FB27
FB0D
FB4D
FBA3
FB8A
FB13
FAE2
FB45
FBBA
FBAD
FB53
FB59
FBCA
FBD8
FB18
FA80
FBA7
FEED
02CA
053F
05B5
0538
04FB
0526
0524
04BE
046A
0490
04F3
0510
04D7
04B0
04D0
04F3
04D4
04A3
04BB
0505
0507
049D
0447
047F
04F2
04E1
0440
03F7
04AC
0585
04AF
0164
FD0E
FA19
F9A4
FAB4
FB8B
FB72
FB06
FB01
FB58
FB85
FB57
FB12
FAF1
FAE8
FAE8
FB11
FB65
FB8F
FB47
FAD7
FAE3
FB85
FC06
FBC8
FB35
FB3E
FBF0
FC26
FB1F
F9F8
FADD
FE89
0317
05C8
05BF
048C
041E
04BA
054A
0518
0499
048E
04F3
0534
0517
04EF
04FD
050D
04E3
04B3
04D4
051F
050C
0476
03F3
0412
0493
04B5
044C
041A
04B4
0568
04A1
01B2
FDDA
FB31
FAA1
FB3D
FB8E
FB2B
FAC5
FAF0
FB5E
FB6A
FB04
FAAF
FABC
FAE9
FAE4
FAC4
FAD2
FB07
FB1A
FB0A
FB29
FB8B
FBB8
FB4D
FABB
FAE5
FBDF
FC8D
FBFA
FADA
FB29
FE01
0220
0509
057E
048B
0411
04B2
0581
057E
04CF
045B
048B
04F7
0521
0514
0522
054E
0553
0522
0501
0513
0514
04CA
0476
0484
04D4
04C7
0434
03DC
0477
056A
04FE
0235
FE23
FB08
FA22
FAB4
FB3C
FB26
FAF4
FB1D
FB5A
FB2C
FAB2
FA7B
FAC1
FB1D
FB18
FAC5
FA8F
FAAE
FAF5
FB28
FB44
FB58
FB5C
FB42
FB2B
FB4A
FB8E
FB96
FB23
FAAB
FB39
FD89
0125
0480
062D
0602
051A
04A8
04E4
052F
050C
04B5
04A6
04ED
052C
0527
0509
050C
0525
052B
0525
0531
0538
0505
04AA
0488
04C3
04F8
04D9
04BB
0527
05B7
0506
0222
FDFF
FADD
FA1A
FAF0
FB91
FB25
FA5E
FA40
FAE3
FB8E
FBB2
FB66
FB10
FAE7
FAE0
FAE4
FAE7
FAE3
FAE2
FAEF
FAFD
FAEC
FACB
FAE2
FB43
FB7D
FB23
FA9E
FB28
FD95
012F
042F
0563
0530
04CF
04F2
0559
0584
0554
04FE
04BA
04A5
04CA
0511
053C
051E
04E0
04CD
04EF
0509
0507
0516
0536
051A
04AC
047A
0509
05C1
0518
0235
FE31
FB3C
FA7B
FB1D
FB95
FB4E
FAD0
FAAF
FAD7
FAEF
FAE1
FADB
FAF9
FB2B
FB55
FB5D
FB2E
FAE3
FAD3
FB2A
FB7E
FB3A
FA7E
FA31
FAC7
FB78
FB36
FA62
FACD
FDA1
01C7
04DA
059A
04F1
0473
04A0
04EB
04F1
04F4
0531
0565
0541
04EB
04C3
04DB
04F1
04E7
04DB
04D8
04BB
0494
04AB
04FC
0512
04BE
0498
0533
05E5
04FF
01BB
FD87
FAD0
FA91
FB88
FBEC
FB5C
FAC2
FACF
FB3A
FB5E
FB19
FABE
FA97
FAA9
FAD2
FAEC
FADF
FAC5
FAE9
FB63
FBC0
FB83
FAEA
FAC9
FB52
FB98
FAE0
FA16
FB2C
FEBC
02F6
055F
0566
049D
048F
051B
0542
04C8
045E
047C
04D6
0503
050B
0526
053C
051D
04E5
04D2
04C6
047E
0430
046E
052D
058E
0511
047F
04D8
0591
04BF
016C
FD23
FA78
FA4C
FB29
FB51
FAB4
FA68
FADF
FB78
FB8C
FB3C
FB02
FB00
FB0B
FB13
FB2F
FB59
FB72
FB71
FB61
FB24
FAB0
FA72
FAF6
FBE5
FC0D
FAED
F9EC
FB27
FEF7
033B
0580
056F
04AB
0496
0508
053B
051E
0524
0551
053D
04DA
048C
0480
0468
0420
0412
0496
053C
0552
04EA
04C1
0509
0514
0491
0455
051E
05E6
049D
00B6
FC4A
FA02
FA4F
FB55
FB6A
FACA
FA9C
FB23
FB9A
FB77
FB0A
FAD9
FAFA
FB3B
FB7D
FBA6
FB8B
FB30
FAF2
FB16
FB4E
FB1F
FAB8
FACD
FB6B
FBA2
FAE9
FA5D
FBCF
FF81
0387
05B4
05BA
0502
04BB
04D2
04BE
0484
047E
04A8
04B9
04BC
04F1
053F
0535
04C2
0463
047C
04C1
04B6
0479
048A
04E8
0508
04D0
04E5
0583
0593
03A9
FFF5
FC63
FAAF
FABB
FB27
FB21
FAF7
FB16
FB42
FB22
FAEE
FB0D
FB5F
FB6B
FB2B
FB0A
FB33
FB4C
FB1C
FAFB
FB46
FBAD
FBA3
FB44
FB33
FB78
FB49
FA6C
FA33
FC37
0034
03E9
0567
04F5
044E
0477
04F4
0504
04C3
04BE
04FE
051A
04F5
04DC
04EE
04E8
04A4
045F
045B
047B
0486
0488
04A0
049B
0442
0403
04A1
05DD
060D
03B9
FF82
FBC7
FA4F
FAB6
FB5C
FB56
FB02
FAF8
FB2D
FB4E
FB55
FB5F
FB4B
FB03
FAD6
FB22
FBAD
FBDF
FB9C
FB71
FBBB
FC05
FBC1
FB3B
FB30
FB8F
FB6D
FAA1
FA98
FCD4
00CC
0437
0575
051D
04CD
0522
0566
050B
047E
0463
04A1
04BB
04A4
04A8
04C5
04B2
0471
0462
049A
04A9
044D
03F3
041B
0485
048F
0454
04A1
0570
0542
02BE
FEA2
FB4F
FA4B
FADD
FB50
FB03
FAA0
FABD
FB17
FB43
FB5F
FBA2
FBCC
FB8B
FB21
FB17
FB6B
FB95
FB62
FB3C
FB6F
FBA4
FB7D
FB50
FB9D
FBF9
FB6F
FA44
FA67
FD57
01FC
0579
062E
0528
0478
04D1
0557
0544
04DF
04B4
04B7
049B
047D
049B
04CA
04B5
0480
049B
04F6
04FB
047F
041F
0462
04D9
04CB
0471
04B5
0575
0508
022C
FDF5
FAE8
FA4C
FB0F
FB79
FB23
FAD6
FB01
FB33
FB13
FAF6
FB3A
FB95
FB8F
FB48
FB34
FB57
FB4E
FB14
FB0F
FB59
FB82
FB4A
FB2E
FB9D
FBFF
FB6C
FA62
FAD4
FDE5
022A
04FE
055E
04A6
048B
0527
0575
0510
0499
049C
04CC
04B6
047E
047B
0494
0482
046C
04A9
050F
0516
04B0
046C
0497
04B5
0460
042E
04E9
05E6
0525
01B3
FD3D
FA7F
FA5F
FB55
FB94
FAF9
FA8D
FAD5
FB57
FB91
FB98
FBA2
FB94
FB64
FB61
FBAC
FBCF
FB63
FAD5
FAE6
FB83
FBCB
FB5A
FAEB
FB28
FB7D
FAF5
FA25
FB12
FEA5
030F
058B
056F
0485
048C
054A
057F
04DC
0446
045A
04A8
0495
0449
043E
0475
049A
04AD
04E6
051C
04F2
0487
0474
04DE
051A
04BB
046F
050A
05D7
04E1
0159
FD00
FA6E
FA4E
FB14
FB38
FAD4
FAD4
FB64
FBD3
FBBF
FB7E
FB62
FB46
FB12
FB1C
FB88
FBCC
FB68
FACC
FAD0
FB6F
FBBF
FB4F
FAD3
FB02
FB55
FAE1
FA31
FB38
FED5
0346
05D6
05C7
04B9
0469
04E0
0520
04C8
0462
0465
04A4
04D5
04FA
050C
04CD
0446
040B
047A
0515
0526
04C0
0491
04C4
04C9
0471
048A
0590
0644
049B
0069
FC1D
FA40
FACA
FBAB
FB8A
FAF4
FAF4
FB75
FBA7
FB5D
FB2A
FB54
FB71
FB3C
FB17
FB4A
FB6D
FB1A
FAB7
FAEF
FB96
FBD6
FB77
FB32
FB71
FB82
FABD
FA23
FBA4
FF96
03CC
05CA
0567
0473
0452
04BC
04D7
0494
0477
049C
04AF
04A5
04CE
0523
0528
04BC
046F
04A5
04E8
04AE
044A
0473
04FE
04FC
0447
040C
050F
05F8
047A
0047
FBEB
FA16
FAC6
FBCF
FBB4
FAF6
FAB9
FB1D
FB6C
FB53
FB22
FB13
FB03
FAF3
FB2F
FBAD
FBD7
FB5E
FAD0
FADD
FB55
FB87
FB5D
FB63
FBA8
FB63
FA5C
FA02
FC21
0074
0468
05CD
0519
046C
04DD
05A0
059C
04EC
0468
046D
04A5
04C9
04E9
04FD
04CF
047E
048B
050C
0555
04E8
044C
0455
04E2
050B
049D
0485
0541
058C
0390
FF6A
FB82
F9FE
FA89
FB38
FB07
FA9B
FACA
FB5D
FB9C
FB6D
FB47
FB57
FB55
FB23
FB0B
FB2B
FB31
FAFE
FAF1
FB41
FB72
FB0D
FA88
FAC0
FB8F
FBC2
FAE9
FA8A
FC96
00D2
04B3
061B
0577
04B7
04D2
0528
04FC
0489
0465
0492
04AF
04B1
04D7
050D
04F7
04AA
04B4
0538
058E
053D
04C2
04CF
0523
04FC
0473
0486
0565
0579
0315
FECF
FB42
FA36
FADC
FB4E
FAFC
FACB
FB45
FBC6
FB9C
FB0E
FAD4
FB00
FB1A
FB03
FB15
FB5A
FB5B
FAF9
FAC8
FB27
FB88
FB4A
FAD0
FAF2
FB89
FB76
FA85
FA64
FCD4
012F
04BC
05A9
04DA
045E
04DA
0559
0525
04B6
04BC
050D
051D
04E9
04E2
0513
050A
04A4
045F
0492
04EB
0501
04FB
0523
0539
04DC
046A
04A7
055A
04F9
0258
FE61
FB5E
FA8E
FB0D
FB52
FB08
FADB
FB0F
FB28
FADF
FAA0
FAD9
FB4E
FB7C
FB5E
FB4F
FB57
FB20
FAAF
FA88
FAE4
FB40
FB24
FAE1
FB05
FB57
FB2B
FABE
FB7E
FE5E
024C
0504
056F
049E
043E
04B7
0541
0550
0522
0511
0503
04CD
04A6
04D2
0526
0536
04FA
04D4
04F2
050A
04E4
04C6
04F3
052D
0518
04F0
052B
0560
0435
00EE
FCCF
FA39
FA44
FBAA
FC58
FBAF
FACB
FAC3
FB62
FBAD
FB40
FAA1
FA73
FAB6
FB04
FB25
FB29
FB1F
FAFA
FAD2
FAEE
FB63
FBCD
FB9F
FADD
FA68
FB68
FE40
01FE
04F6
060D
0583
0490
043C
0497
0504
050F
04DD
04CF
04FA
0521
0516
04EB
04CB
04CE
04F3
052B
0547
04FE
044F
03C9
0424
0545
05DD
0472
00F6
FD1C
FADD
FAB4
FB76
FBCE
FB87
FB3D
FB45
FB4A
FAFD
FAA7
FABD
FB21
FB3D
FAD9
FA77
FAA1
FB1F
FB46
FAEB
FAB6
FB38
FC05
FC15
FB29
FA72
FB8F
FED8
02D0
0563
05B5
04AB
03D7
0403
04C0
053A
0531
0504
0504
0510
04E9
04B0
04B7
0501
052C
0507
04E1
0513
0556
050F
0450
0402
04B7
057D
048D
014A
FD3C
FAAA
FA63
FB35
FB90
FB26
FABC
FAD8
FB21
FB18
FAD4
FAC4
FB01
FB37
FB3E
FB53
FB99
FBB4
FB3D
FA7C
FA4F
FB19
FC13
FC0E
FAEE
FA27
FB6E
FEF1
02F2
055A
058C
04B4
0451
04BF
0540
0529
04B1
047D
04C3
051C
052D
0517
051B
051C
04CE
0455
043F
04C6
054C
0510
0442
03F7
04BB
057A
0462
00EE
FCC5
FA40
FA28
FB40
FBDC
FB98
FB44
FB76
FBCB
FBA2
FB15
FAC9
FAF5
FB15
FABC
FA4E
FA7C
FB3D
FBBD
FB79
FAF6
FB0B
FBA2
FBC1
FB03
FA8B
FBFA
FF86
0372
05B4
05D7
0510
04A6
04B9
04A4
0431
03E6
0439
04E3
053D
0518
04EA
0510
0550
0535
04C8
0492
04D4
0514
04C0
041B
0414
04F3
058B
042F
0096
FC79
FA09
F9E3
FAC8
FB3C
FB03
FAE5
FB57
FBE1
FBE0
FB67
FB0F
FB1D
FB3C
FB1D
FAF2
FB12
FB56
FB46
FAD9
FAB6
FB58
FC33
FC2C
FB0F
FA46
FB9F
FF4E
0372
05D1
05E4
0505
04B4
0517
054E
04E2
045B
045F
04C4
04DE
0484
044A
049E
0521
052F
04D1
04AC
04FB
0524
0499
03DB
03FE
0518
05A6
03FB
0038
FC65
FA7E
FAA7
FB67
FB76
FAEA
FA9F
FAEC
FB4C
FB38
FAE0
FAD6
FB39
FB8E
FB6F
FB14
FAF8
FB27
FB37
FAFF
FAEB
FB61
FBF2
FBC5
FAD6
FA83
FC46
FFFD
03BA
0590
0552
0467
0423
049B
0518
0531
0520
0527
0531
0513
04EA
04F0
0511
04F9
049A
0465
04BA
0555
057C
04E6
0433
043E
04F9
0522
0366
FFD6
FC1C
FA15
FA33
FB48
FBDF
FB93
FB07
FADB
FB00
FB10
FAF9
FAFD
FB2C
FB40
FB15
FAF8
FB33
FB83
FB5B
FABC
FA5B
FAC0
FB75
FB89
FAED
FAEB
FCDD
0089
0419
05CD
0590
04BA
0480
04E8
0536
0506
04AC
0495
04B9
04C5
04A1
048D
04AD
04D5
04D0
04C0
04E8
0532
0531
04C2
046C
04C9
0583
0544
0301
FF42
FBE3
FA67
FAAB
FB52
FB48
FAB5
FA68
FABF
FB4A
FB7C
FB52
FB37
FB5F
FB90
FB82
FB4A
FB30
FB49
FB5D
FB4B
FB42
FB6A
FB7D
FB0F
FA64
FAA0
FCC9
007F
0400
05B1
0588
04D3
04B6
0528
056F
053C
04EB
04DA
04EC
04D1
048D
0466
0470
0473
044F
0443
0486
04DC
04CF
0464
043E
04D6
05A6
055A
030C
FF53
FBE9
FA41
FA5D
FB11
FB47
FAE8
FA96
FAB9
FB09
FB0F
FAD6
FAD3
FB35
FBA5
FBC3
FBA8
FBA3
FBAC
FB72
FB03
FAF5
FB96
FC36
FBD4
FAA7
FA68
FCA2
00C6
0478
05D7
0538
0469
049D
0567
05BE
0561
04F2
04F5
0538
0542
0500
04BD
04A1
048D
0466
0457
0486
04BA
0492
041F
03FD
0497
0561
050E
02CA
FF3E
FC20
FAB5
FACB
FB28
FAF7
FA72
FA4C
FAAF
FB1A
FB16
FAC7
FA9F
FAC5
FB02
FB2F
FB64
FBAE
FBD4
FBA5
FB5C
FB62
FBB4
FBBE
FB20
FA72
FAF1
FD4C
00CA
03DC
056A
059B
0554
0538
0542
052C
04FC
04FC
0542
0580
0560
04FD
04C0
04D3
04E3
049B
042F
042A
04A3
0502
04C7
045C
049F
057F
0584
033D
FF15
FB47
F9C5
FA65
FB67
FB80
FAFB
FAC9
FB16
FB39
FACF
FA53
FA6E
FB08
FB72
FB4E
FAF9
FAF7
FB41
FB69
FB46
FB23
FB3C
FB4C
FAF4
FA82
FB02
FD4C
00F6
0467
061F
05F2
04FF
047B
04A9
0504
051C
050B
0517
0530
0513
04C9
04AC
04DD
0508
04E3
04A9
04CF
053F
0558
04E0
0485
0509
05E8
0572
0297
FE5C
FB1A
FA33
FAE4
FB67
FAF8
FA51
FA66
FB1E
FB96
FB58
FADB
FAC9
FB22
FB62
FB4B
FB30
FB5D
FB90
FB48
FA91
FA24
FA7B
FB1A
FB1B
FA8D
FAD2
FD37
0148
04E2
0634
0578
047B
048C
054C
0596
0512
0480
048D
04F7
0515
04CE
049D
04BE
04CD
047A
0427
0473
0539
0597
0522
0499
04F7
05E7
05AC
02FB
FEA5
FB0C
F9DE
FAA3
FB90
FB83
FAD7
FA7F
FAC9
FB40
FB71
FB6C
FB6A
FB64
FB34
FAFF
FB1C
FB90
FBDF
FBA1
FB18
FAED
FB43
FB6F
FADB
FA18
FAA5
FD65
016C
04A2
05B5
0533
04A7
04DD
054F
0533
04AB
047B
04E7
0543
04EB
0435
0408
049F
052A
04DF
0417
03D9
0479
0528
0515
0497
04A4
053E
04FD
029A
FEAC
FB58
FA35
FAD7
FB95
FB76
FAEC
FAD2
FB34
FB70
FB3A
FB05
FB46
FBBA
FBC6
FB5C
FB1A
FB6E
FBEF
FBE6
FB4E
FAE6
FB23
FB80
FB40
FABE
FB66
FE1F
01F1
04BF
0563
04B1
0451
04D9
0574
0547
0496
0451
04BD
0531
050A
0483
0443
0462
0465
0419
03FD
0483
053F
054A
048F
040F
0498
0565
04A8
0198
FD8E
FAD5
FA65
FB33
FBA3
FB47
FAE2
FB14
FB85
FB8B
FB21
FAE9
FB3D
FBBF
FBE5
FBAF
FB90
FBB6
FBC6
FB6F
FAFB
FB03
FB99
FC07
FBB2
FB11
FB89
FE0E
01EC
052C
0649
057D
044F
03F7
0464
04C7
04BF
049A
04AE
04CC
04A5
045D
045B
04A2
04B9
046F
0439
0481
04E7
04AE
03E9
03AE
04A2
05AF
04D4
016C
FD29
FA81
FA4A
FB43
FBC8
FB79
FB14
FB29
FB76
FB80
FB4A
FB39
FB74
FBB0
FBAA
FB7F
FB77
FB98
FB9C
FB5E
FB1D
FB33
FB87
FB8C
FB03
FAAA
FBCB
FEDA
02A1
0522
0573
048A
041A
04BD
0593
0590
04C8
042A
0445
04B9
04DD
048C
042B
040B
0428
0469
04C7
0527
0534
04C4
043A
043B
04D5
0523
0402
013E
FDE6
FB7F
FABC
FB14
FB78
FB58
FAEF
FAB9
FAD4
FB04
FB1A
FB27
FB45
FB60
FB62
FB70
FBB3
FBF7
FBC8
FB1A
FA9B
FAF1
FBD0
FC21
FB63
FA9A
FB79
FE89
0264
04F8
0574
04C5
0457
04A3
0518
0520
04DD
04D9
0536
057F
0547
04B8
0454
044B
0457
0440
043B
0490
0507
0517
04B5
048C
050B
0565
041C
00C8
FCE7
FA90
FA75
FB77
FC1C
FBEB
FB5C
FADF
FA87
FA6A
FAB7
FB4B
FB97
FB5C
FB18
FB5F
FBEE
FBF3
FB4A
FACE
FB2A
FBC0
FB75
FA7E
FAA3
FD42
017C
04DB
05D4
0512
044F
0461
04D2
04F9
04DD
04E6
0524
0546
0523
04E2
04AC
047D
0459
046D
04AF
04BD
0458
03FE
047B
05AA
0605
03FF
FFE7
FBFA
FA44
FAAE
FB74
FB59
FACB
FACC
FB61
FBA3
FB29
FA9F
FABB
FB39
FB58
FB0A
FAFB
FB66
FBAA
FB4D
FAD1
FAF1
FB5C
FB23
FA75
FB0B
FE2A
02A1
05AF
05F9
04D4
0458
04ED
0565
050A
0489
04B4
053C
0547
04CB
0487
04CC
0506
04C5
047D
04BD
0530
051B
04AB
04D5
05A1
0576
02D4
FE7C
FB04
FA20
FAF7
FB90
FB41
FAF4
FB51
FBB7
FB52
FA80
FA5C
FB20
FBCD
FB93
FADC
FA97
FAE5
FB22
FB0A
FB0A
FB4E
FB3D
FA89
FA51
FC3E
004D
044B
05F7
0559
045D
0459
04CE
04B9
043C
044A
0501
0564
04E0
0436
046A
0542
05A3
0530
04BB
04EC
0542
04F8
046B
0496
0536
0481
014B
FCEB
FA16
FA00
FB4C
FBFA
FB96
FB1B
FB2E
FB6E
FB5D
FB2F
FB41
FB62
FB25
FABA
FAB6
FB1E
FB44
FAD9
FA8C
FB08
FBCA
FBB5
FAE5
FB19
FDBD
01E7
050A
05A8
04BA
042E
04A4
052C
04F4
0460
044D
04C8
0523
0503
04CA
04E0
0512
0505
04D5
04DA
04FE
04D1
0463
046B
051F
0550
036B
FF83
FBBA
FA2F
FAC9
FB9F
FB5D
FA99
FA94
FB5C
FBD4
FB64
FABC
FAC6
FB57
FB91
FB34
FAE3
FB15
FB6A
FB62
FB30
FB4B
FB79
FB1B
FA84
FB3C
FE50
02A6
05BF
0645
053F
048E
04C9
051B
04DE
047F
04A4
0518
0529
04BC
046E
0496
04D5
04BB
0482
0497
04D9
04CE
0493
04D2
0585
0555
02EC
FED2
FB44
F9F8
FA7C
FB1F
FB0C
FAD7
FB28
FBA0
FB7F
FAE1
FA98
FB00
FB87
FB94
FB53
FB43
FB64
FB5A
FB30
FB4C
FB99
FB5E
FA7B
FA42
FC49
004E
040A
0577
04E1
0427
0461
04F4
04F1
048A
0491
0519
055A
04EE
046C
0476
04CB
04CA
0480
0488
04ED
04FD
0473
0427
04E4
05CD
04E1
015E
FD04
FA70
FA71
FB8F
FC12
FBBB
FB56
FB43
FB27
FAD4
FABA
FB29
FBAE
FBA3
FB2A
FAF9
FB4B
FB8D
FB4E
FB01
FB46
FBCA
FB93
FAA3
FA94
FCF5
0135
04D9
05FE
0521
0435
044B
04CD
04D7
0480
0478
04D9
0508
04B7
0460
0485
04E8
04F8
04AD
0488
04B2
04BD
047F
0488
0534
0592
0405
0045
FC33
FA19
FA5C
FB5D
FB94
FB1D
FAFB
FB75
FBD8
FBA6
FB40
FB34
FB63
FB50
FAFD
FAE9
FB39
FB77
FB50
FB1B
FB3D
FB60
FAF4
FA6F
FB57
FE87
02C7
05B7
062B
0525
0468
0489
04D4
04AE
045C
0459
0492
04A3
0494
04BD
0517
0529
04CE
048B
04CD
0534
0519
04AD
04C6
056A
0525
0293
FE56
FAD8
F9D1
FAA1
FB66
FB47
FAF6
FB33
FBA4
FB8F
FB11
FAF1
FB61
FBB3
FB69
FAF2
FAF3
FB43
FB3B
FAD2
FAB2
FB15
FB46
FAD2
FAB8
FC8F
005E
0417
05AD
053A
0487
04B6
0538
0520
049E
049A
052E
057C
04FD
044D
0440
04B6
04EB
04B6
04AB
050F
054C
04F2
0494
04F6
0581
0479
011D
FCFB
FA7C
FA5E
FB38
FB77
FB0C
FADB
FB2B
FB5F
FB1A
FAD0
FAFF
FB5D
FB62
FB24
FB2D
FB7A
FB6D
FADD
FA90
FB1D
FBD5
FB8A
FA78
FA96
FD5E
01C7
0523
05E8
0510
0482
04DA
053F
04FF
0480
0473
04CE
0501
04E4
04D4
04F3
04EE
049B
0466
04B2
0521
0508
0488
0489
0553
059B
03B4
FFB2
FBBB
F9F3
FA5B
FB33
FB2D
FAA2
FA9A
FB3C
FBC0
FBA4
FB48
FB33
FB4B
FB2A
FAE8
FAFB
FB6C
FBAA
FB5D
FAEE
FAE4
FB00
FAB2
FA5C
FB6E
FEB9
0303
05EB
0655
055B
04C8
0519
0574
0532
04AD
047C
0495
0495
0483
04BA
0521
052E
04C0
046F
04B3
051B
04FF
04A6
04F2
05C7
0584
02C0
FE4C
FAAE
F98E
FA34
FAD5
FABF
FA9D
FAFE
FB75
FB68
FB0B
FAFB
FB48
FB69
FB30
FB0C
FB45
FB6C
FB17
FAB0
FAEA
FB85
FB69
FA5A
F9E7
FBEE
0039
0462
063F
05FC
0560
0573
05A6
052C
0462
043D
04DE
0563
0530
04B4
04A8
0501
0522
04E6
04CB
050F
053D
04FB
04C8
0542
05C9
04B1
013E
FCF0
FA39
F9F8
FAD7
FB26
FABC
FA97
FB19
FB8A
FB47
FABC
FAAF
FB19
FB42
FAE6
FA90
FAB6
FB0F
FB1B
FAF6
FB10
FB42
FAF5
FA5E
FAE7
FDAA
01CB
04FD
05D5
0513
0477
04C2
0554
0572
053A
0526
053B
0524
04E4
04D4
050D
053D
052F
051F
0543
0558
0505
0498
04C4
057D
0577
0363
FF95
FBFC
FA56
FA9B
FB5E
FB75
FAF2
FA8D
FA9E
FADB
FAF6
FAFE
FB1C
FB3A
FB26
FAE7
FAB5
FAAA
FAAF
FABF
FAFB
FB55
FB62
FAE9
FA9B
FBC6
FEEB
02CC
0558
05AC
04D4
046A
04E0
0566
0554
04F9
04F2
052E
0521
04B7
047E
04CD
0541
055B
0528
0504
04EB
04A7
0478
04E1
0591
0514
0257
FE45
FB2F
FA6C
FB12
FB6A
FB01
FAB2
FB03
FB60
FB27
FAB1
FAC2
FB4D
FB86
FB1E
FAB8
FADE
FB30
FB15
FAD1
FB19
FBC2
FBBA
FABF
FA58
FC55
006B
042F
05A0
0523
048E
04CC
0531
04FB
0484
0492
050F
053B
04DE
04A0
04F5
055E
0530
04A8
0493
0508
0534
04AC
043E
04C2
057A
047B
010B
FCE1
FA7D
FA8B
FB7C
FBA7
FB0A
FAB0
FAFE
FB59
FB43
FB14
FB3B
FB7B
FB51
FADD
FABD
FB14
FB54
FB22
FAEA
FB25
FB6D
FB0B
FA5F
FB03
FDF1
0206
04EE
0586
04CF
046C
04CB
0533
0520
04E8
04F4
0508
04B8
043B
0431
04B6
052E
0521
04E0
04F0
052F
0519
04BB
04CC
056A
0560
033F
FF50
FBB4
FA4C
FADB
FB9C
FB79
FAF3
FAF1
FB5A
FB70
FB16
FAF7
FB67
FBCD
FB86
FAE3
FAB5
FB08
FB20
FABB
FA8D
FB19
FBAD
FB5C
FAB7
FB9C
FEE4
02FA
0563
0570
04AA
04A4
0536
054C
04AC
0429
044E
04B2
04C6
04A6
04BB
04FA
0506
04E6
0503
055E
0559
04AF
041D
0483
0568
051A
0289
FEA1
FB7E
FA5E
FAB1
FB18
FAEE
FAA2
FAC5
FB45
FBA5
FBA9
FB7F
FB5E
FB42
FB1A
FAF9
FAFF
FB12
FAFC
FAD3
FAF3
FB59
FB64
FAC0
FA68
FC06
FFE9
0420
0638
05C4
0498
0477
0535
0582
04F5
0469
047A
04AE
0481
0459
04C8
056A
0569
04CF
0489
04F7
0557
0510
04D0
0566
05F4
047A
008F
FC6E
FA8D
FAEE
FB9F
FB69
FAD8
FACE
FB21
FB2A
FAF2
FB04
FB66
FB7E
FB1E
FAD1
FAEC
FB12
FB00
FB0F
FB63
FB55
FA86
FA1F
FBDA
FFBB
0398
0559
051D
0496
04B8
0507
04F4
04D9
0517
0543
04EF
048D
04B9
0522
050D
049F
04A8
053C
0563
04AF
042E
04DA
0593
0414
000B
FC03
FA71
FAFD
FB91
FB3E
FAD1
FAF6
FB2D
FAEA
FA97
FADA
FB64
FB6C
FB00
FAEE
FB58
FB73
FAF7
FAB9
FB35
FB83
FAE6
FA93
FC83
00A8
047C
05D1
0520
0471
04AF
0513
04F6
04D0
0519
054D
04E6
0465
0484
04F1
04E5
0480
0491
0523
0554
04D8
04A1
0540
0557
02FB
FE96
FAFF
FA38
FB35
FBAB
FB0D
FA8F
FAE2
FB53
FB38
FAF4
FB26
FB8B
FB7E
FB15
FAFD
FB49
FB5B
FB11
FB04
FB50
FB26
FA65
FAA2
FD6A
01D8
0524
05B6
04B6
043B
04CB
0553
0519
04A3
0498
04CA
04D1
04D1
0506
051E
04CA
046E
048C
04DE
04D0
049A
04FB
05B0
0517
0212
FDD9
FAF8
FA89
FB45
FB82
FB23
FAF8
FB30
FB4C
FB29
FB1C
FB2B
FB06
FABA
FAC7
FB42
FB8A
FB40
FAF9
FB53
FBB3
FB18
FA25
FB0B
FEB0
0309
0543
04F7
0420
0443
04E6
04FC
04A1
04AA
051F
053A
04CA
048E
04E7
0535
04F2
0498
04B5
04E6
049F
045D
04E4
0589
0463
00C6
FC98
FA70
FABA
FBA1
FBA6
FB2E
FB2F
FB84
FB6A
FAEA
FAB6
FAFA
FB35
FB28
FB1E
FB3D
FB3E
FB0C
FB13
FB79
FB8E
FADC
FA80
FC4E
004D
0417
0575
04CD
042D
0488
0510
04F1
0486
048C
04F0
0519
04F3
04ED
0514
0500
04B4
04B4
04FD
04DA
043D
0437
0540
05BC
038F
FF09
FB13
FA03
FB23
FC07
FBA6
FB0D
FB38
FBA0
FB6A
FAE1
FAD5
FB32
FB3E
FAE6
FAC1
FAFF
FB2C
FB18
FB2A
FB86
FB86
FAE3
FADA
FD18
014B
04EB
05F2
0507
043C
0473
04E1
04CB
0481
0493
04E0
04F5
04C9
04B0
04BD
04C7
04DB
0520
0544
04D2
0435
0476
0572
0540
025D
FDE8
FAB3
FA2F
FB29
FBB1
FB62
FB26
FB6A
FB97
FB4A
FAFF
FB25
FB61
FB45
FB17
FB34
FB51
FB12
FAE2
FB51
FBE1
FB8A
FA98
FB07
FE32
02AD
0589
059D
048E
044E
04D1
04EF
047B
0446
049C
04E4
04C4
04A8
04E1
050B
04C7
0478
04A1
04E3
0487
03F4
044B
0547
04C8
016D
FCDB
FA22
FA45
FB7D
FBCE
FB3C
FAFA
FB5D
FBA3
FB63
FB21
FB43
FB68
FB35
FB0B
FB42
FB7C
FB53
FB2A
FB79
FBC7
FB58
FACC
FBF2
FF7B
03A0
05CF
057F
0473
044A
04CD
04FB
04BC
04A3
04C6
04C4
049C
04A1
04CB
04BE
047F
0487
04E1
04F2
047C
0449
04FA
0575
03C0
FFB9
FBC8
FA3B
FAC5
FB6E
FB46
FB01
FB40
FB90
FB5D
FAF7
FAFC
FB46
FB40
FAFF
FB21
FB9E
FBAA
FB22
FAED
FB71
FBAE
FAEA
FA7C
FC7C
00CA
04B3
05EB
050D
045F
04D8
056A
0521
0485
047B
04D8
04F2
04D3
04E9
050F
04D4
046A
0467
04B5
04A9
0442
046D
0569
0599
0327
FEA9
FB02
FA25
FB0F
FB92
FB16
FA9E
FAC9
FB1F
FB2C
FB2D
FB60
FB74
FB24
FAD8
FB10
FB7A
FB6E
FB20
FB58
FBE9
FBAA
FA94
FAA6
FD8E
021B
0549
05AB
04AD
0453
04DA
052C
04E5
04B7
04FE
052A
04DD
049D
04D5
050C
04CC
048B
04D6
0524
04AC
03EF
0436
0559
0532
0226
FD92
FA8E
FA5C
FB54
FB7C
FAEC
FAD4
FB4F
FB74
FAFF
FAA7
FADB
FB2D
FB31
FB22
FB47
FB55
FB09
FAE2
FB6C
FC0A
FB9C
FA9C
FB40
FEB5
0328
05AC
0587
048A
0469
04F5
0525
04DA
04C0
050C
053F
0521
0512
0534
0519
04AB
048D
04F5
051C
047D
03FD
049D
0576
044A
006C
FC13
FA06
FA8A
FB86
FB6D
FACC
FABC
FB17
FB17
FAC3
FABD
FB08
FB1A
FAE2
FAE2
FB35
FB54
FB12
FB0E
FBA3
FC01
FB57
FAA1
FC06
FFFC
042A
05FB
0577
04A9
04CE
0547
0535
04D5
04DC
053E
055C
0514
04E0
04F3
04F3
04C1
04B8
04DF
04AE
041F
041D
050A
0576
037B
FF4B
FB6C
FA07
FAB7
FB79
FB41
FABB
FAB6
FAF5
FAED
FAC7
FAF3
FB48
FB52
FB20
FB0D
FB14
FB00
FB09
FB8B
FC1A
FBBB
FA86
FA5A
FCF9
0191
052F
05F1
04DF
042C
0491
052D
0552
0544
0552
0546
04F4
04AD
04C0
04ED
04E0
04CF
050A
052B
0496
03CD
041F
0571
058F
02AB
FDF8
FA92
FA11
FB24
FBB4
FB52
FAEE
FAFD
FAFC
FAB1
FAA7
FB21
FB7D
FB45
FAF7
FB24
FB6A
FB34
FAE3
FB37
FBD8
FB9F
FAA3
FAE8
FE04
02AE
05CE
05FA
04CA
0462
04E9
0537
04F5
04D4
0517
052C
04CD
0486
04C2
0519
04FF
04B1
04BB
04F1
04BA
0454
04A2
0553
0480
0109
FC93
F9F5
FA0A
FB21
FB77
FB16
FAFC
FB4B
FB4E
FADD
FAAB
FB12
FB79
FB5B
FB14
FB1B
FB39
FB23
FB2F
FBA5
FBDB
FB25
FA70
FBC3
FFAF
0413
0637
05C8
04CC
04C9
0539
050E
0487
0487
0507
053E
04F9
04C4
04D6
04CF
048D
0485
04E2
0503
0482
042D
04E0
059F
0420
FFE1
FB67
F98B
FA49
FB5A
FB4D
FAC9
FADB
FB52
FB63
FB0B
FAF2
FB37
FB4E
FB15
FB18
FB81
FBB2
FB63
FB3B
FB96
FBAA
FADE
FA6D
FC55
0093
049E
0619
055E
0495
04DB
055F
0535
04C4
04C8
050B
04F1
04A5
04B5
04FE
04EE
048F
047B
04C4
04CC
046D
0478
0542
0564
0311
FEB7
FB11
FA1C
FAF5
FB7D
FB14
FAB2
FAE4
FB1B
FAE0
FAA4
FAEC
FB67
FB75
FB2B
FB21
FB61
FB6A
FB3B
FB5F
FBB6
FB5A
FA5A
FA90
FD81
020A
0548
05D5
0500
04B8
0536
0569
04FC
04BC
0517
0566
051C
04AE
04A9
04BF
047E
0446
049C
050D
04D0
0440
0486
0587
0544
022C
FD89
FA68
FA1F
FB11
FB39
FA9E
FA79
FAF8
FB30
FACF
FA8B
FADE
FB52
FB60
FB44
FB6C
FBA2
FB71
FB19
FB37
FB8F
FB3F
FA8D
FB4E
FE9E
02FD
05B7
05EC
0518
04DD
0537
0544
04E0
04B3
04FA
0534
0513
04EC
0500
04FB
04A9
0475
04A9
04D2
0490
0470
0504
0577
040F
0067
FC66
FA4F
FA5D
FAF4
FAF1
FAC1
FB0B
FB6D
FB43
FAD5
FADB
FB42
FB54
FAEF
FAAF
FAE4
FB24
FB16
FB18
FB7B
FBB3
FB2D
FAC0
FC3B
FFFC
03F4
05D3
0588
04D4
04E3
0545
0535
04D6
04C3
050A
0535
0519
0501
0508
04F8
04D2
04EC
053A
052B
049F
0461
04DE
04FE
0329
FF6C
FBC9
FA23
FA61
FB09
FB32
FB1D
FB22
FB05
FA9D
FA62
FAB3
FB20
FB15
FACA
FADF
FB47
FB57
FAEF
FABA
FB17
FB5C
FAFC
FAEF
FCE3
00E6
04C4
0658
05D3
0507
0500
0536
0502
04BB
04FE
058C
05A4
0531
04DB
04F5
0504
04B0
0478
04E6
0585
056F
04BB
0488
0544
0598
03C1
FFCA
FBD1
F9EA
FA24
FAF2
FB24
FAE3
FAD8
FB0D
FB09
FAAF
FA6F
FAA0
FB09
FB3B
FB32
FB39
FB58
FB3D
FACF
FA8D
FADC
FB52
FB3A
FADB
FBA5
FE96
02AC
059A
061A
0522
048B
04EB
055D
0529
04BF
04DA
0555
0575
0515
04CA
04E7
0507
04CF
0499
04E1
0553
0530
0493
047B
0528
0527
02D6
FEA7
FB0B
F9E1
FA95
FB31
FAD5
FA56
FA9E
FB4E
FB70
FAEB
FA93
FAE7
FB70
FB8B
FB47
FB1D
FB24
FB13
FAEB
FB0B
FB76
FB83
FADC
FA7B
FC00
FFB6
03CE
0604
05E6
0505
04F5
05A2
05E8
0550
049D
049A
050A
052A
04CF
0484
04A2
04D7
04CB
04AE
04D0
04FA
04C7
0470
049F
0527
0493
01B7
FD78
FA50
F9BA
FABF
FB60
FAEF
FA65
FAA0
FB33
FB49
FAED
FAD4
FB26
FB4D
FB05
FADD
FB4B
FBD0
FBAB
FB11
FAEC
FB69
FBA1
FB1A
FB0A
FD19
011A
04C6
061D
0578
04B9
04E5
0559
053D
04CC
04C6
052E
0555
04FE
04B0
04D0
04F6
04A4
042D
0443
04D8
0517
04B0
0465
04DD
053C
03CF
0033
FC3D
FA2B
FA5C
FB43
FB72
FAFE
FAC2
FAEF
FAFC
FAAC
FA7A
FAC7
FB38
FB48
FB1A
FB36
FB9C
FBAF
FB33
FACD
FB13
FB86
FB3E
FA8D
FB2B
FE39
028A
0594
060F
0510
0470
04BA
0529
052D
051F
0561
0598
0548
04B6
0498
04F6
051C
04AF
0444
047A
04FC
0503
04A2
04BD
0573
0557
02F3
FECD
FB36
F9E7
FA70
FB26
FB26
FADB
FAD6
FAF3
FAD7
FAAC
FAD5
FB30
FB3E
FAF1
FAD3
FB30
FB96
FB7B
FB19
FB1D
FB82
FB77
FAAC
FA4C
FBFD
FFD2
03D7
05EB
05CB
04F1
04BC
0522
0553
0504
04AE
04B6
04EA
04F1
04DD
04EF
0517
0503
04B9
04A1
04D9
04F1
0499
044D
04BB
0571
04CB
01C3
FD78
FA62
F9D3
FACE
FB7A
FB37
FAD3
FAFD
FB60
FB5E
FB0C
FAF8
FB32
FB3F
FAF7
FAD0
FB1C
FB6E
FB46
FAEB
FB03
FB76
FB6D
FAC2
FAC8
FCFD
0107
04B2
0622
059B
04C0
0496
04CB
04C9
04A6
04CB
0521
052D
04DE
04A7
04CF
0500
04DD
049C
04B1
0505
050E
04BB
04B1
0541
0579
03DA
002F
FC33
FA08
FA2A
FB3A
FBB0
FB52
FAE8
FAF7
FB34
FB2C
FAF1
FAE0
FB14
FB54
FB70
FB6C
FB4D
FB0D
FAD7
FAFC
FB6F
FB89
FADA
FA2C
FB20
FE6E
02B6
059E
0614
0525
0489
04D1
0542
0534
04DD
04BC
04D5
04D0
04A1
0488
048F
0480
0461
0490
051A
0565
04F8
0458
0488
0576
0585
0339
FF1E
FB76
F9F8
FA4C
FAEB
FAF6
FABF
FACC
FB04
FB15
FB12
FB41
FB8B
FB90
FB57
FB52
FBAB
FBE5
FB8C
FAF9
FAE6
FB55
FB6E
FAC8
FA6B
FBE5
FF69
034B
0598
05E3
0548
04F1
0507
0516
04F0
04CB
04C8
04C6
04B7
04BF
04E2
04D9
047D
0424
0442
04B8
04E5
0490
0461
04F9
05B2
04E5
01BE
FD86
FA99
FA19
FB00
FB8B
FB29
FAAB
FAD1
FB53
FB7A
FB33
FB05
FB2E
FB59
FB49
FB46
FB99
FBEF
FBBF
FB2F
FAF8
FB4E
FB74
FAF6
FAD8
FCBB
00AD
048D
062B
058E
0498
049E
052A
052D
04AB
047B
04DA
0519
04C9
046C
0494
04F0
04D7
046A
0462
04D8
0505
0489
0434
04CD
057A
044E
00BA
FC95
FA37
FA0F
FAB2
FAEC
FAE7
FB2B
FB81
FB5A
FADC
FAC4
FB41
FBA6
FB73
FB1A
FB38
FB93
FB7A
FAF4
FACC
FB49
FB99
FB02
FA4E
FB43
FE86
0295
0537
05B2
0527
04F8
0555
058F
0548
04DE
04CB
04FE
050F
04D2
0487
0472
0488
04A2
04BD
04E2
04F2
04D4
04C5
051C
0591
0506
0289
FEA3
FB4A
FA1B
FAC3
FB86
FB41
FA74
FA36
FAB1
FB20
FB06
FAC1
FAD4
FB28
FB57
FB59
FB74
FB98
FB6A
FAFE
FAE7
FB47
FB64
FAC5
FA69
FC03
FFD1
03DA
05DA
0594
04B8
04AC
052C
054A
04F3
04DA
053A
058A
055F
0508
04F2
04F8
04BC
0465
0474
04E6
0513
04B3
0472
04F8
059B
04BA
01A3
FDA6
FAE1
FA38
FAC7
FB39
FB2B
FB12
FB38
FB54
FB18
FAB4
FA89
FAA4
FAC9
FAE0
FB0C
FB4C
FB61
FB2E
FAFB
FB18
FB46
FB01
FA76
FAD9
FD33
00F8
043E
0590
0541
04B9
04C7
050C
04F9
04B2
04B9
0507
0527
04FF
04F9
0545
056B
050F
049D
04BB
0542
055E
04DC
0499
052C
058E
03FA
003A
FC52
FA78
FAC9
FB91
FB82
FAEB
FAB1
FAED
FB0B
FAE1
FADD
FB2D
FB5F
FB1D
FACD
FAF3
FB4E
FB2F
FAA2
FA7D
FB1D
FBA7
FB2F
FA65
FB31
FE70
029C
053D
057A
04AA
046A
04E0
0528
04EE
04C8
0522
0581
0546
04A6
0461
04AD
04F9
04E4
04C7
0510
0566
052C
049B
049D
054C
0537
02E6
FEDE
FB70
FA50
FAE8
FB6D
FB1E
FAC0
FB0E
FB8E
FB65
FAB4
FA6D
FAF1
FB90
FB97
FB3C
FB23
FB57
FB56
FAFF
FAD0
FB01
FB0C
FA9A
FA8D
FC4E
FFF3
03B0
058F
0566
04AD
049E
0508
0520
04C5
0486
04B2
04FE
051A
051C
0523
04FC
0482
0420
0462
0511
0555
04E6
049D
0539
05E4
04C0
012A
FCE6
FA73
FA7A
FB69
FB9A
FB0D
FACD
FB35
FB9B
FB74
FB11
FAEF
FAF6
FAD5
FAC6
FB45
FC0C
FC27
FB48
FA6C
FA92
FB49
FB48
FA87
FAC2
FD70
01A6
04D7
0599
04E9
048E
04F0
052D
04CA
0464
049B
051C
0536
04EC
04D3
050B
0504
047B
0409
0453
0506
0542
04EA
04CB
053F
0540
036E
FFEB
FC7F
FACD
FAC3
FB18
FB02
FAD0
FAFE
FB4F
FB3D
FADB
FABF
FB20
FB81
FB71
FB2F
FB35
FB6F
FB5C
FAF8
FAE9
FB74
FBDD
FB5F
FAA3
FB71
FE91
0285
04F7
0536
04A8
04C9
057D
05AC
0514
048F
04B8
0513
04F5
048F
0485
04CD
04CB
0468
045C
04FD
057E
0503
0414
0413
0516
053A
02CA
FE8A
FB20
FA33
FAE6
FB5B
FAF5
FA8B
FAC7
FB45
FB5F
FB28
FB20
FB51
FB57
FB2A
FB2E
FB7F
FB9F
FB35
FAB2
FAC9
FB59
FB83
FB03
FAF4
FCBC
0048
03D8
05B7
05C4
052A
04E4
04ED
04D5
0496
048D
04D9
0523
0520
04EC
04CB
04C1
04A6
048A
049E
04D1
04D4
04A2
04B2
053C
0571
03FD
009B
FCD2
FA9C
FA6F
FB0A
FB26
FACF
FAD0
FB40
FB6A
FAF7
FA88
FAC8
FB65
FB89
FB1D
FAE7
FB52
FBBD
FB7B
FAF0
FB03
FBA9
FBD3
FB20
FAED
FCEF
00F7
04C4
0657
05E4
051F
050F
053F
04FC
0483
0495
0538
059D
053A
0488
045E
04CC
0517
04C6
0444
0446
04CC
0522
04DE
0476
049D
0518
04A1
0239
FE7A
FB3B
F9E1
FA34
FAE6
FB11
FADC
FAD0
FAFE
FB0B
FAE3
FADF
FB32
FB8B
FB7E
FB27
FB0A
FB55
FB9E
FB74
FB08
FAEE
FB4D
FB93
FB36
FAB0
FB51
FDEB
01B9
04D8
05EF
055A
049D
04C1
0570
05B3
0546
04C8
04C3
04F3
04D0
0470
0469
04D8
0516
049F
03F2
03FF
04D2
0565
050A
0471
04B0
057A
0508
0221
FDD4
FA9F
F9F1
FADF
FB7B
FAFC
FA36
FA36
FAF0
FB8A
FB87
FB44
FB46
FB81
FB7E
FB26
FAEE
FB30
FB9B
FB97
FB23
FAE3
FB33
FB85
FB1D
FA68
FAFD
FDEE
023E
0587
0654
056C
04AE
04ED
056E
0548
04A1
044B
048B
04D4
04B8
0486
04BA
0525
0520
048A
0414
0456
04FB
051F
0493
042E
04B0
0575
04D2
01DE
FDB9
FAA0
F9D3
FA8F
FB33
FB09
FAB0
FAE5
FB6D
FB86
FB10
FAB9
FB00
FB81
FB92
FB3A
FB1C
FB71
FBAB
FB4D
FAC5
FAEC
FBBB
FC21
FB65
FA71
FB1D
FE31
0259
0557
060C
0544
0496
04C9
0563
058F
0528
04B5
04AE
04F0
0508
04CF
048D
0482
0490
0480
046F
04A8
0509
050F
0498
044F
04D2
0582
04BD
01A6
FD79
FA8C
FA02
FAD5
FB47
FAD3
FA52
FA85
FB19
FB4E
FB0E
FAEE
FB40
FBA6
FBA6
FB5D
FB44
FB70
FB75
FB19
FABE
FAEB
FB78
FB9C
FAF6
FA5F
FB59
FE75
027C
0563
0628
058E
0507
0527
0563
0523
04A3
0483
04D4
04FB
049D
0425
042A
0497
04D7
04B3
0497
04E3
0544
0526
049D
046B
04F6
056E
046E
0172
FD96
FAAF
F9C9
FA68
FB3C
FB65
FB11
FAF0
FB41
FB94
FB76
FB13
FAFC
FB5D
FBBA
FB98
FB27
FAFA
FB31
FB56
FB22
FAF0
FB20
FB5B
FB0C
FA96
FB6C
FE75
029B
0589
05FF
04F9
0451
04A7
051D
04E3
0459
0459
04F1
0552
04FE
0477
047E
0502
0540
04DE
046B
0490
0518
0537
04B2
044D
04B7
054E
0478
0176
FD87
FADD
FA70
FB32
FB84
FB03
FA99
FAF5
FB95
FB93
FAF7
FAA4
FB0F
FB98
FB78
FAE3
FAC2
FB58
FBDC
FB8D
FAD6
FABE
FB70
FBE1
FB41
FA64
FB1F
FE3D
0263
054A
05E2
0511
046C
049F
0523
053F
04E7
0498
04A2
04DE
0505
050E
0511
0508
04CE
0470
0442
0479
04D1
04D7
0492
049D
0547
05C2
049E
0154
FD3C
FA86
FA2D
FB1F
FB99
FB0E
FA72
FAB5
FB83
FBC9
FB2F
FA80
FA89
FB1B
FB6A
FB37
FB07
FB3C
FB7A
FB41
FACD
FACF
FB56
FB8D
FAF4
FA71
FBA5
FEFE
02F3
056A
05BC
050C
04C6
0525
0568
0517
049E
049D
0510
055E
0528
04B9
048E
04B2
04C4
049B
048E
04EF
056D
0561
04BF
0458
04C8
054E
0440
00ED
FCC7
FA31
FA1B
FB38
FBB0
FB1E
FA8D
FAC3
FB4C
FB4E
FACB
FA87
FADF
FB55
FB62
FB2F
FB37
FB6D
FB57
FAE7
FAB3
FB24
FBBA
FB96
FABC
FA70
FC0E
FF8E
0358
059D
05D8
0504
0482
04D0
0555
0551
04D6
0495
04E7
0556
054A
04DF
04AF
04EC
051C
04DD
048A
04AC
050F
04FB
0466
0440
050A
05A3
043E
0094
FC8F
FA6A
FA77
FB2E
FB31
FAA2
FA6C
FAD3
FB42
FB40
FB02
FAF2
FB1B
FB38
FB28
FB08
FAF4
FADF
FAC4
FACD
FB28
FBB4
FBFD
FB9E
FACB
FA7A
FBD3
FF14
02FC
05A1
061A
0545
04B6
0507
058B
057C
0504
04CF
04F5
04F2
0493
045B
04B9
0542
0540
04C0
0485
04E7
0545
04EF
0445
0454
0546
05BA
0413
0055
FC5E
FA2E
FA2A
FB0E
FB68
FAEA
FA64
FA91
FB3E
FBA0
FB5E
FAF2
FAF5
FB55
FB7F
FB39
FAF5
FB1F
FB6D
FB53
FAEA
FADC
FB47
FB5E
FAA2
FA26
FBBE
FFB9
040C
0632
05C5
049D
0481
054E
05B5
052A
0473
0463
04CC
04F2
04A5
0465
048D
04D7
04D6
04A3
04AA
04FA
0520
04DA
0491
04E2
059D
0592
039B
FFED
FC36
FA34
FA36
FB09
FB61
FB0A
FAB5
FADE
FB3D
FB54
FB2C
FB32
FB7A
FB9F
FB66
FB29
FB54
FBB2
FBA8
FB1A
FAB2
FAF8
FB7C
FB50
FA76
FA50
FC4F
0038
0416
05FB
05BC
04C1
046D
04D8
052A
04E1
0464
045C
04C9
0514
04E0
0485
0487
04D5
04E3
047B
041B
044B
04D8
051A
04E9
04DF
054F
0557
0396
FFE7
FC02
F9F6
FA32
FB48
FBAC
FB3C
FAE8
FB38
FBAF
FBA1
FB27
FAE4
FB1D
FB68
FB59
FB1E
FB29
FB78
FB96
FB4A
FB00
FB28
FB7D
FB4D
FA9F
FAA2
FC92
0038
03CE
059E
0591
04EF
04CB
050F
050E
04A6
0461
049B
04FC
0502
04C1
04BE
051F
055D
04FD
044B
0409
0473
04EF
04E4
0499
04D1
0589
0580
0367
FF86
FBD1
FA29
FA97
FB7D
FB73
FAA1
FA2C
FAAA
FB81
FBCE
FB7C
FB27
FB2B
FB3C
FB07
FAC8
FAF0
FB68
FBA2
FB64
FB1F
FB4C
FB9B
FB51
FA82
FA76
FC75
003E
03F9
05E4
05D4
0509
04B9
0502
0545
0522
04D1
04AC
04AE
04A3
0497
04C4
0524
054C
04F7
047F
047F
0500
0556
0503
0485
04C3
0598
0583
032B
FF1B
FB86
FA1E
FA86
FB16
FAE2
FA7E
FAC6
FB8A
FBD9
FB5F
FACD
FADB
FB51
FB6F
FB0A
FAC2
FB0F
FB88
FB72
FACF
FA72
FADB
FB75
FB52
FA92
FAAD
FCFA
0107
04B1
061E
0570
046A
046B
052A
0572
04D1
0417
0432
04FD
058B
0564
04FC
04E7
0504
04DE
0482
047D
04FE
0571
0551
04F9
0525
059E
0506
0253
FE4F
FB16
FA13
FAC4
FB94
FB98
FB2B
FB06
FB42
FB70
FB54
FB26
FB18
FB03
FAB6
FA66
FA86
FB1F
FBA1
FB83
FAFA
FAC5
FB2C
FB7F
FAF3
F9FA
FA42
FD05
0174
0528
065F
0590
0495
0490
0502
04F6
046D
0438
04A6
0515
04E9
047C
049C
0554
05C6
0560
04B4
04AE
053D
0568
04BD
0420
04A8
05E1
05D4
0320
FEB2
FB12
F9F0
FAAE
FB71
FB39
FA9C
FA9A
FB3F
FBB7
FB7D
FAFC
FAE0
FB2E
FB56
FB18
FAD7
FAF6
FB36
FB17
FAAD
FA9D
FB1C
FB72
FAE2
FA03
FA87
FD66
0192
04CE
05D3
054E
04C4
04E7
053C
0526
04B9
0479
049A
04D7
04F3
04FA
050D
0518
04F4
04AF
048F
04B9
04FA
0503
04DD
04ED
0566
05BF
04E5
023E
FE85
FB6E
FA39
FAA1
FB4B
FB43
FAC7
FA98
FAE9
FB40
FB45
FB2E
FB47
FB6C
FB53
FB1F
FB38
FB93
FB91
FAE7
FA3C
FA65
FB30
FB83
FADA
FA42
FB58
FE72
0215
0470
04FD
049C
045C
048C
04E3
0520
053C
0542
0524
04E0
049F
049E
04E3
0521
0508
04A7
046E
04B1
052A
0530
0499
0425
049E
0590
054F
02B6
FEA0
FB47
FA26
FAC0
FB85
FB91
FB2B
FAE6
FADA
FADD
FAF9
FB42
FB88
FB7F
FB3B
FB19
FB39
FB5B
FB44
FB16
FB11
FB32
FB4F
FB68
FB84
FB5D
FAB7
FA30
FB20
FE2F
022D
04F8
0582
04B0
041B
045E
04E6
0519
0501
04F3
04FB
0500
050E
0522
0503
0491
0427
043C
04B8
050B
04EC
04B7
04C6
04E0
04B3
0497
051E
05CB
0511
020F
FDFE
FB22
FA7F
FB1E
FB88
FB5E
FB25
FB1D
FAF7
FA99
FA6C
FAB8
FB25
FB48
FB42
FB68
FB9F
FB8B
FB3A
FB1B
FB45
FB47
FAEE
FAB1
FAF3
FB2F
FAB5
FA25
FB3E
FEBB
02EF
055D
055A
047C
046E
0525
0583
0523
04B1
04C4
0518
052D
0501
04DC
04BF
0490
047F
04C0
0518
0519
04D4
04C8
0510
052A
04DC
04CE
058D
0623
04B2
00D0
FC84
FA4A
FA76
FB4A
FB51
FAD4
FAC9
FB3E
FB71
FB20
FAD7
FAFD
FB3D
FB31
FB0E
FB29
FB4D
FB16
FAB8
FAC2
FB3B
FB82
FB4B
FB08
FB17
FB03
FA57
F9F5
FB8B
FF6A
039B
05CD
05B8
04F5
04C7
04F4
04D1
0484
04A8
052B
0557
04F3
049A
04C8
0528
053B
0521
0531
053B
04DD
045C
0476
0538
05B2
054C
04BA
04EB
0541
03EB
0053
FC54
FA51
FA94
FB64
FB60
FADD
FACF
FB3C
FB6B
FB21
FAE2
FAFF
FB1C
FAE6
FAAC
FAD3
FB24
FB2F
FB06
FB0F
FB3B
FB21
FACA
FAD0
FB58
FB93
FAF2
FA84
FC21
FFFE
03E8
058F
04FB
0423
045F
052E
0578
0521
04D8
04EC
050A
050D
0539
058F
058D
04FA
0471
0494
051D
054E
0506
04CF
04D7
04AC
0434
043B
052F
05CD
041D
0002
FBEB
FA4B
FAF5
FBC7
FB6F
FAA2
FA8F
FB1D
FB5B
FAFE
FAA8
FAC0
FAEC
FAD7
FACF
FB24
FB73
FB3E
FACE
FAD0
FB42
FB69
FAFD
FAA2
FADF
FB31
FAF4
FAE0
FC96
005F
0439
05DC
053B
0443
0461
0524
056B
0507
04B6
04E7
053D
054E
052A
0500
04C5
0482
0488
04EE
0539
0503
04A6
04BE
0527
0523
04A6
049E
0570
05B9
0395
FF40
FB59
FA17
FAED
FBA4
FB31
FA7C
FA8A
FB0A
FB20
FADB
FAF3
FB79
FB9F
FB0E
FA85
FABA
FB4C
FB6A
FB18
FB06
FB64
FBA0
FB6B
FB32
FB48
FB3D
FAC2
FAD4
FCEF
00E8
047F
05B3
04FA
0463
04F8
05D6
05D0
050B
048B
04B7
0512
0527
0518
051B
0510
04E8
04E5
0515
050B
0485
040A
043B
04C3
04BC
0425
0419
0510
0584
036C
FEFD
FAEF
F999
FA85
FB84
FB73
FB04
FB10
FB50
FB1C
FA99
FA7C
FADC
FB1C
FAF3
FAD3
FB0D
FB44
FB1F
FAF9
FB4A
FBCA
FBD6
FB81
FB78
FBC5
FB9C
FACE
FAD4
FD52
01B8
0555
0637
052D
0463
04B2
0533
0511
04B4
04D3
0547
0561
050F
04E1
0516
053C
0506
04C9
04D2
04DD
049C
045F
048D
04D5
04A2
043A
048E
0585
055C
0287
FDF9
FA8E
F9F2
FAF8
FB73
FAE5
FA7D
FAF4
FB96
FB7C
FADB
FA86
FAB6
FAEE
FAE9
FAED
FB23
FB42
FB28
FB2D
FB76
FB88
FB0E
FA9A
FAEB
FB9F
FB92
FAC1
FAF0
FDB3
0224
058B
0655
058A
0508
0534
0529
0496
043E
04AF
0561
0583
0520
04DD
04ED
04ED
04B9
04AC
04EF
0518
04E6
04C3
0506
0538
04C8
0427
0459
052F
04E0
0209
FDB1
FA78
F9C4
FA87
FB05
FAE7
FAFC
FB87
FBD8
FB74
FACF
FA97
FACF
FB0C
FB26
FB48
FB5F
FB31
FAE2
FAED
FB54
FB7C
FB26
FAFA
FB7E
FC0B
FB9E
FAB6
FB4F
FE8A
02ED
05B9
05E5
04E6
048C
04F3
0517
049B
0429
0443
04A0
04D7
04FF
0544
0561
0507
0486
047F
04EB
051D
04CB
0483
04B3
04E8
0498
0436
0495
0542
0477
0137
FCEE
FA3A
FA1B
FB22
FB74
FAE5
FA90
FB05
FBAD
FBCF
FB7B
FB33
FB32
FB54
FB6C
FB68
FB3B
FAF4
FADD
FB2B
FB8C
FB7E
FB22
FB2F
FBC8
FC01
FB2C
FA4C
FB62
FF01
0343
05A0
058B
04A5
0481
050B
054D
0503
04BE
04DE
0515
0505
04C7
049C
0490
0495
04BE
0506
051E
04CB
046F
049D
051D
0511
044D
03EB
04C8
05D5
04D1
0102
FC6F
F9E2
FA00
FB0E
FB58
FAFD
FB05
FB9D
FBF3
FB90
FAF7
FACB
FAFB
FB10
FAF5
FAFD
FB43
FB7B
FB63
FB1C
FAE9
FAE5
FB1E
FB98
FBF9
FBA9
FAAF
FA43
FBE5
FF9F
039F
05D8
05EB
0521
04BF
04DB
04E2
04A3
046B
0472
04A1
04DC
0522
0557
054A
04FE
04C0
04B8
04B2
0483
046C
04B6
050C
04D0
0430
042E
0521
05AB
03FB
0016
FC2D
FA61
FA9E
FB30
FB06
FAA2
FAD4
FB6A
FBA5
FB69
FB41
FB60
FB57
FAE4
FA77
FA92
FB0A
FB4A
FB2C
FB16
FB45
FB7F
FB99
FBC6
FC0A
FBE6
FB27
FACD
FC50
FFD8
03A4
05A9
0594
04C3
047E
04C3
04EA
04C9
04BE
04F1
0523
0520
0504
04F0
04E0
04D0
04DB
04FA
04F0
04A7
0478
04B0
04F3
04AB
0411
041B
04FA
0538
032C
FF24
FB73
FA11
FAB2
FB91
FB9E
FB47
FB3F
FB69
FB4B
FAF6
FAD6
FAF7
FB05
FAF8
FB1E
FB79
FB9B
FB56
FB19
FB4F
FBA1
FB76
FB03
FB0F
FBA4
FBC1
FAF9
FAB0
FCBA
00E3
04BA
061F
0567
0486
0494
04F5
04D1
0466
046C
04E3
052E
0516
04F6
0504
0505
04D2
04A9
04C1
04DE
04BA
0484
0495
04BD
048E
043E
048E
055D
0520
028B
FE7B
FB59
FA89
FB1D
FB5F
FAF0
FAC0
FB4D
FBE1
FBBB
FB2C
FAF2
FB1B
FB23
FAEB
FAD7
FB09
FB2A
FB15
FB1F
FB74
FB9F
FB3E
FAD2
FB25
FBE6
FBE3
FAFD
FAFB
FD86
01CC
0519
05CF
04F6
0487
04FF
0554
04E3
044F
0456
04B7
04CD
04A0
04AF
04FC
050F
04D3
04BE
0500
0525
04D4
046E
0479
04B4
0486
0425
0474
0558
0519
0247
FDD2
FA65
F9A0
FAA5
FB8A
FB85
FB29
FB0D
FB14
FB0A
FB28
FB8E
FBD8
FBAC
FB57
FB4D
FB6A
FB37
FAD0
FAD6
FB63
FBBD
FB64
FAEA
FB1E
FBA5
FB6B
FA92
FAF0
FDE4
0242
055C
05ED
052D
04E7
055A
058D
0514
0496
04A5
04E9
04D0
0473
044B
0460
0465
045A
0489
04E0
04EB
0495
0465
04B4
0505
04C3
0451
049B
0566
04F0
01F6
FD95
FA70
F9F0
FB02
FBB5
FB5C
FAC3
FAAF
FAF2
FB05
FAE4
FAF0
FB41
FB8D
FB9A
FB7B
FB5D
FB5A
FB7E
FBAA
FB9A
FB31
FAD3
FB11
FBD5
FC36
FB98
FACD
FB89
FE70
0224
0499
0520
04B9
0498
04EA
052C
0522
0509
050B
0503
04E1
04DA
0508
0521
04E1
0473
043D
0452
0474
0488
04AA
04BF
046F
03D1
03B1
049A
05A1
04DC
0181
FD31
FA85
FA70
FB86
FBE5
FB48
FAD1
FB31
FBC1
FB93
FACC
FA69
FAE0
FB95
FBB8
FB47
FAEA
FB05
FB5D
FB94
FBA7
FBC2
FBDA
FBBA
FB6D
FB41
FB51
FB4E
FB08
FB0D
FC5C
FF44
02C7
0549
05F6
0554
0488
0439
044C
046E
0491
04C3
04E3
04C0
0473
045F
04AF
0514
051C
04BE
0463
0459
047B
0479
0453
0455
0495
04C0
0490
044C
046E
04C8
0445
01F4
FE4A
FB0E
F9C3
FA4A
FB40
FB8F
FB5C
FB57
FB9C
FBAB
FB4D
FAFC
FB2C
FB96
FB99
FB2C
FAF1
FB43
FBB8
FBC7
FB9D
FBC1
FC23
FC15
FB5F
FAC8
FB0F
FBB5
FB9F
FAE3
FB39
FDF7
0220
052E
05C6
04F3
048C
04FA
0539
04B2
041C
045B
0528
057B
0501
046E
0469
04B5
04BC
047B
0467
049D
04AE
0458
0408
043C
04BE
04E5
0493
0471
04F4
056B
0480
01A9
FDF7
FB3D
FA70
FAF9
FB90
FB88
FB2D
FB0E
FB32
FB32
FAE5
FAAD
FAF2
FB7E
FBB9
FB76
FB2D
FB4A
FB9A
FB9D
FB51
FB34
FB7E
FBC2
FB9B
FB5C
FB8D
FBEE
FBAD
FADB
FB01
FD84
01AB
04FD
05CE
04EB
0453
04C6
054D
0509
0482
04B4
057C
05C2
051A
045F
0475
0511
053E
04C8
0468
0495
04C9
0466
03C3
03BB
0461
04CF
0477
0400
0457
0523
04CF
0250
FE84
FB75
FA64
FADC
FB90
FBBF
FB8B
FB54
FB2A
FAEA
FA9D
FA81
FAB1
FAFB
FB1D
FB16
FB19
FB3A
FB62
FB7F
FBB0
FC0A
FC54
FC2F
FB9F
FB2B
FB3C
FB79
FB39
FAAB
FB23
FDB8
01B9
04F2
05CB
04D1
03E2
0408
04AF
04E5
04B4
04D3
0564
05B3
0548
04A1
0481
04E0
0505
049C
0428
0435
0489
048A
0435
041B
0478
04CA
04A1
0466
04D4
05A2
0559
02D5
FECD
FB60
FA21
FABF
FBBA
FBFD
FB9F
FB36
FAFA
FAC6
FA94
FAA6
FB17
FB95
FBBD
FB96
FB78
FB8D
FBA1
FB83
FB60
FB7A
FBB3
FBA2
FB37
FAF5
FB3C
FB9E
FB55
FA85
FA96
FCD4
00CA
045B
05BC
051A
041B
03FC
048A
04EF
04E7
04DD
0513
053C
0508
04AB
0497
04D6
0500
04D4
0489
046C
0470
045E
044C
0483
04F3
0515
049F
0416
044B
0522
0546
0367
FFC6
FC3B
FA8C
FAD1
FBAF
FBE7
FB74
FB1C
FB46
FB91
FB7E
FB24
FAF9
FB24
FB50
FB34
FAFA
FAF3
FB28
FB56
FB5C
FB57
FB52
FB25
FAD9
FADC
FB7A
FC2D
FBFE
FAE4
FA5F
FC20
000B
0402
05E2
0589
0494
045C
04B9
04C9
0461
042A
048E
051C
0535
04DE
04A4
04CD
050D
0512
04F1
04E8
04E7
04BA
047A
0487
04EE
0536
04FB
0498
04C3
0575
057A
0389
FFC4
FBED
F9DD
F9EE
FAED
FB84
FB68
FB30
FB4E
FB89
FB83
FB4E
FB4A
FB89
FBAC
FB71
FB0D
FAE5
FAFE
FB17
FB19
FB36
FB77
FB80
FB17
FAA3
FABF
FB48
FB60
FAB9
FA76
FC31
0006
040A
0619
05E2
04EC
04A6
050C
053F
04F3
04AE
04DB
0524
0504
0491
045C
049B
04E2
04C4
046D
045B
04AB
04FA
0503
04F9
0516
0523
04C7
0441
0452
0524
0595
0416
0073
FC64
FA07
F9E7
FAC9
FB48
FB32
FB26
FB60
FB6C
FB01
FA8E
FAA9
FB34
FB86
FB59
FB1C
FB42
FB9A
FBA3
FB57
FB23
FB36
FB3A
FAF4
FAC4
FB21
FBB9
FBA5
FAB7
FA3C
FBD5
FF97
03A2
05DC
05D6
04E1
0468
04A5
04F6
04FF
0509
0551
0587
0541
04AE
046B
04AE
04F9
04C6
0446
041C
047B
04E9
04F4
04D3
04FB
0556
0556
04E1
04A4
0511
055C
0408
00B0
FCD4
FA85
FA61
FB37
FB92
FB30
FACC
FAD9
FB00
FADA
FA9A
FAB6
FB26
FB6E
FB5C
FB4F
FB9B
FBF5
FBD4
FB43
FAE2
FB07
FB45
FB18
FABF
FAEC
FB99
FBD3
FB0A
FA44
FB52
FEB8
02D2
0561
05BB
0516
04DB
052B
054B
04F1
049D
04C0
0513
050D
04AC
046A
0485
04B5
04A5
0472
0473
04AB
04C6
04A4
048C
04B8
04E3
04A4
042C
0442
0537
060B
0518
01CB
FD8E
FA9E
F9FE
FAC1
FB55
FB28
FAD7
FAFF
FB6A
FB89
FB57
FB4E
FB97
FBC0
FB6B
FAE9
FAD1
FB34
FB92
FB98
FB84
FBA9
FBD9
FBB3
FB53
FB40
FB90
FB95
FAD2
FA17
FB01
FE2F
0246
0515
05A5
04E9
046B
04AE
0515
0506
04B4
04A1
04D4
04E8
04B4
0485
049B
04BE
0494
0440
043C
04A5
04FC
04D1
046F
046F
04D1
04EE
0480
043C
04D9
05B2
050D
01FF
FDCC
FAD8
FA53
FB43
FBE3
FB88
FAE1
FAB9
FB05
FB41
FB3A
FB35
FB66
FBA4
FBB1
FB93
FB7E
FB87
FB90
FB7E
FB5C
FB39
FB10
FAEC
FAF9
FB54
FBBA
FB9C
FACC
FA1A
FAF0
FDF7
021C
053E
0614
0545
0477
0489
04F8
04FC
04B1
04C6
054B
057F
04EE
0429
0408
0482
04C5
0473
0421
0474
052B
0579
0528
04CD
04D3
04E3
049C
0468
04E6
05A2
0506
021A
FDF2
FAE3
FA37
FB15
FBB9
FB66
FAC3
FAA6
FB08
FB5B
FB5E
FB4F
FB58
FB52
FB26
FB0F
FB48
FB98
FB88
FB0F
FAB7
FAE4
FB4A
FB4F
FAEC
FABF
FB1C
FB77
FB1E
FA75
FAF5
FDA4
01B0
04F6
05FD
053F
0460
0466
04EF
0519
04BD
0476
04AE
0511
0514
04C1
049F
04EA
0532
0503
0493
047B
04DB
0531
0514
04C5
04B1
04C3
04A6
0488
04FB
05CE
058C
02EB
FE9F
FB18
FA0B
FACE
FB77
FB34
FADB
FB41
FBF5
FBFC
FB4A
FAC0
FADC
FB20
FB00
FAC5
FB00
FB82
FB89
FAED
FA77
FAD0
FB8B
FBC0
FB51
FB0F
FB7F
FBF9
FB8E
FA8F
FAA8
FD1B
0133
04BB
05FF
0546
043B
0421
04C7
052F
04EB
0477
046A
04B5
04E5
04DE
04EE
0531
054B
04EE
046D
0455
04AC
04E9
04CE
04BE
0509
0542
04D9
0428
042C
04FF
0524
0301
FEF0
FB41
F9E8
FA9E
FB93
FB9E
FB26
FB05
FB4B
FB65
FB25
FAF2
FB12
FB35
FB01
FAB3
FACF
FB58
FBB5
FB84
FB1F
FB12
FB52
FB63
FB25
FB17
FB84
FBDB
FB56
FA53
FA7A
FD14
015E
04F6
0618
0538
0439
0454
051D
0583
0537
04D2
04D7
0515
0516
04DA
04C2
04F5
0522
0505
04CA
04C0
04DE
04D8
04A8
04A5
04F7
0536
04F2
0474
0484
052C
0526
030D
FF24
FB74
F9DE
FA56
FB40
FB65
FAFB
FAD2
FB0E
FB25
FADF
FAB4
FB02
FB70
FB6F
FB06
FAC1
FAE2
FB1E
FB1D
FAFB
FAFA
FB0F
FB01
FADF
FAFA
FB50
FB62
FAE9
FA7F
FB3B
FD98
00F0
03F3
05A1
05D4
0533
049D
048C
04D8
0507
04E3
04AC
04BC
0509
0545
0550
054F
0552
0531
04E5
04AF
04BE
04DF
04D5
04C0
04E4
0511
04D6
0455
0462
0546
05B1
03D7
FFB0
FB86
F9AD
FA2C
FB2C
FB51
FAED
FAE8
FB45
FB5E
FB0A
FAD4
FB06
FB2E
FAE1
FA71
FA7D
FB03
FB6D
FB62
FB1B
FAEA
FAE3
FAF7
FB27
FB58
FB49
FAF5
FAD1
FB3F
FBD9
FBD5
FB58
FBC4
FE36
01FD
050A
0604
056F
04B8
04A4
04EA
0516
0521
052F
052C
04FF
04D9
04F4
052F
0539
050F
04F5
0507
050C
04DE
04AE
04B7
04DD
04E2
04D0
04DD
04E7
0492
0406
040E
04E8
055E
03BC
FFE9
FBF2
FA10
FA69
FB45
FB42
FAAB
FA76
FAC8
FAFD
FACF
FAAE
FAF0
FB43
FB3B
FB08
FB24
FB8F
FBCF
FBA8
FB64
FB44
FB25
FAF1
FAF0
FB4B
FB9A
FB6D
FB11
FB2F
FBAF
FBB8
FB27
FB68
FDF9
022E
0574
0614
04FF
045C
04E6
059B
058E
0517
04F4
051C
04FF
049B
0479
04C0
04E8
04A6
046E
04AB
0506
04EA
0474
043C
046B
049B
048E
0477
046E
0432
03CD
03F4
04F8
0597
03EA
FFD6
FBBC
FA01
FA8D
FB5C
FB35
FABA
FAE8
FB7D
FB94
FB1C
FAE3
FB3D
FB87
FB40
FAD8
FAF2
FB5E
FB84
FB5D
FB64
FBAF
FBCC
FB93
FB71
FBAC
FBD2
FB79
FB1A
FB71
FC2A
FC16
FB1E
FB13
FDA8
0212
058E
0655
0546
0468
0489
04F1
04F3
04D2
04FC
0531
04FD
048D
0475
04C2
04EF
04B3
045C
0449
0466
0472
0471
0490
04B9
04B2
048F
04A3
04DA
04BE
044A
0432
04CD
050B
0358
FFA8
FBF7
FA49
FA93
FB29
FAF5
FA87
FAC0
FB65
FB93
FB2A
FAEF
FB52
FBCE
FBC3
FB5F
FB39
FB6C
FB85
FB59
FB44
FB70
FB80
FB2F
FAD8
FAEF
FB46
FB6A
FB6A
FBAB
FBFC
FBA2
FAB5
FAD1
FD79
01EE
0582
0668
0575
04B2
04DD
0528
04EC
049A
04C1
050E
04DE
0454
042D
0490
04D4
048D
0435
0462
04DC
050F
04EF
04E0
04F6
04E8
04B4
04B0
04DA
04B9
043B
042B
050D
05BA
0432
0025
FBD6
F9CA
FA30
FB34
FB7D
FB55
FB72
FBA8
FB5F
FAC1
FA96
FB13
FB87
FB72
FB36
FB55
FB9A
FB89
FB40
FB3D
FB84
FB94
FB44
FB01
FB14
FB2C
FAFF
FAED
FB66
FBE6
FB7A
FA80
FAE9
FE08
028E
05A8
05F9
04C8
041B
0471
04D7
04AB
0461
0492
0504
0522
04E4
04BD
04D3
04E0
04BC
0499
049E
04A3
0486
0479
04AF
04F8
04FC
04C6
04AA
04B2
048C
043F
0464
052B
057E
03DB
0032
FC64
FA73
FA89
FB36
FB51
FB11
FB25
FB81
FB8D
FB2E
FAF1
FB2E
FB8F
FB97
FB4C
FB15
FB19
FB30
FB43
FB6C
FB98
FB88
FB42
FB25
FB52
FB64
FB1A
FAEA
FB5A
FBFB
FBC9
FAD1
FAD0
FD53
018C
04D0
057D
049B
043A
04E9
0588
053F
0498
047A
04D6
04F8
04AB
0478
04B2
0500
04F8
04C4
04BA
04CC
04BF
04A2
04A4
04AB
048C
0479
04C5
0531
0510
045D
0413
04D6
0589
0431
0078
FC7A
FA8D
FACD
FB7B
FB61
FAED
FAFC
FB76
FBA6
FB5A
FB11
FB14
FB1D
FAF4
FAE3
FB2F
FB92
FBA0
FB67
FB3C
FB26
FAFA
FADB
FB1D
FB96
FBA9
FB2E
FAE2
FB64
FC17
FBD0
FABC
FAC1
FD5C
0199
04E5
05C6
051D
04A4
04E9
0532
04EF
0488
04A1
0527
0576
0535
04AA
044D
045A
04B2
0500
04F7
04A3
0471
04BA
0538
0546
04BC
043E
046F
04FB
0504
0471
0434
04D8
0545
03BE
0013
FC3F
FA69
FAB8
FB85
FB81
FAF3
FAC6
FB1D
FB53
FB1D
FAE7
FB17
FB67
FB5E
FB04
FAD9
FB1D
FB82
FBA2
FB74
FB38
FB1D
FB31
FB64
FB7A
FB31
FAB7
FAA5
FB4A
FC03
FBE4
FB20
FB53
FDD0
01D4
0506
05DA
0504
044B
0475
04E8
04F7
04CB
04DE
052A
0541
0506
04D2
04E2
0507
04FE
04C3
0473
042A
0426
04A4
055F
0590
04DC
0404
040E
04E3
0550
04B4
03FF
0455
0509
040A
0092
FC7C
FA50
FA7A
FB46
FB4A
FAD7
FAE4
FB69
FB89
FAFC
FA77
FA96
FB10
FB48
FB35
FB39
FB67
FB77
FB53
FB36
FB42
FB59
FB63
FB6B
FB6C
FB44
FB0C
FB2B
FBBA
FC0E
FB77
FA92
FB1B
FE0A
022A
0526
05DC
052C
0490
0494
04D0
04F5
0527
0578
0596
053E
04B6
047B
04A3
04E1
04EF
04C8
047E
0430
0422
0481
04FF
04FE
045E
03DD
0446
0544
05A1
04D5
03D7
03DB
0475
03C9
00CA
FCC9
FA37
FA18
FB30
FBC1
FB66
FAE9
FAD7
FAE9
FAC4
FA9E
FAD9
FB4A
FB6F
FB2A
FAE8
FAFA
FB33
FB4F
FB5F
FB8B
FBB2
FB99
FB4F
FB24
FB3B
FB75
FBB7
FBEB
FBD2
FB36
FAA0
FB60
FE3E
0223
04CD
0527
045C
043E
051C
05CE
058D
04E6
04B8
04FB
050F
04D3
04C7
0514
0536
04D2
0456
0454
04B9
050C
052B
053E
0534
04D4
0458
0452
04C5
04E0
042D
0382
03FA
0509
0488
013F
FCB7
F9C4
F990
FACF
FBA8
FB9C
FB4D
FB28
FB06
FADB
FAEF
FB4B
FB75
FB1D
FAA7
FA99
FAE5
FB1D
FB2C
FB4D
FB75
FB4B
FAD1
FA9A
FB06
FB9D
FBA6
FB2C
FAE1
FAFF
FB0F
FB06
FBE9
FE89
020E
048F
0534
0502
054B
05E9
05BE
0492
039D
03EE
0512
05BE
0577
04E6
04C2
050A
0553
0566
0547
0505
04BD
04A8
04D2
04EA
04AA
045B
048A
051B
0542
04AC
042F
04A0
054A
044B
00DB
FC91
F9F3
F9EB
FB19
FBA9
FB2B
FA6F
FA31
FA70
FAE1
FB56
FB98
FB62
FABE
FA3B
FA62
FB11
FB9E
FB9C
FB33
FAC7
FA89
FA8E
FAE7
FB6D
FBA7
FB57
FAF4
FB26
FBC9
FBF6
FB5F
FB3D
FD1F
00E5
0483
0620
05E6
0555
0544
054F
0505
04D1
0542
05FB
0608
052E
0451
0452
0506
0597
058A
050C
048A
0463
04C4
0571
05C8
0558
0486
0427
046E
04A1
0444
03FC
0499
055E
044E
00B1
FC71
FA3A
FA8D
FB83
FB58
FA4F
F9CE
FA5A
FB24
FB59
FB0C
FAC3
FAA8
FAAA
FADB
FB39
FB68
FB17
FA92
FA71
FAD0
FB3B
FB67
FB83
FBAA
FB8A
FAF6
FA8C
FB12
FC2D
FC86
FBA0
FAFB
FC9E
0094
0497
0664
05EB
04E1
04A6
051B
0572
0565
0540
052A
04FB
04B8
04BC
053A
05D2
05E8
0553
0486
041C
0457
04FC
0584
0575
04C5
0408
03F7
04A7
0560
056E
04F1
0484
0427
02F8
005D
FD24
FAE9
FA61
FAB5
FAC6
FA8A
FAB6
FB73
FBF8
FB9B
FAB8
FA3C
FA8C
FB2F
FB77
FB2D
FA95
FA21
FA3E
FB03
FBE6
FC18
FB65
FA93
FA7C
FB0E
FB8A
FB95
FB81
FB7F
FB32
FA90
FAC5
FD38
0186
0543
0655
052B
0401
0443
0547
05AA
0519
0469
045C
04DB
056F
05D2
05E7
058A
04CB
0429
0428
04B5
0540
055D
051A
04BC
047A
047D
04E1
057D
05CD
055F
0467
03B8
03FF
0508
05D3
054A
02FC
FF7B
FC32
FA84
FAB7
FBAD
FBF9
FB34
FA3E
FA12
FAB2
FB4A
FB38
FAA5
FA23
FA16
FA88
FB46
FBE1
FBD3
FB0E
FA3F
FA38
FAFF
FBC2
FBC7
FB3A
FAD1
FAE2
FB21
FB47
FB7C
FBDD
FBF5
FB34
F9FF
F9CB
FBD1
FFAB
0371
0553
0520
043C
0420
0500
05E5
05E7
052B
0490
04AB
053A
059E
0596
055D
0528
04F4
04CF
04F2
055F
059B
052E
0452
03CE
040D
049A
04CA
0491
046E
0489
0483
0438
0447
052B
060F
0533
01DB
FD88
FABC
FA86
FB97
FBEA
FAF0
F9D8
F9E8
FB06
FBF8
FBD0
FAC3
F9C9
F9AE
FA77
FB77
FBDB
FB53
FA64
F9FF
FA92
FB98
FC25
FBE5
FB5B
FB26
FB4C
FB65
FB58
FB83
FC13
FC82
FC12
FACB
F9D1
FA8E
FD66
0132
040E
04F1
048D
047C
0576
0694
0679
0516
03D7
03F4
050C
05C2
0575
04C7
047E
048D
0498
04C0
054F
05DE
059B
047C
0399
03E2
04E3
055B
04D7
041C
03EE
0418
0420
0444
0509
05F6
0592
0300
FF3C
FC46
FB3D
FB78
FB88
FAC9
F9DF
F9D1
FADF
FC32
FC94
FB94
FA10
F972
FA45
FBA7
FC44
FBB5
FAB7
FA3D
FA89
FB40
FBE8
FC2F
FBEA
FB34
FA96
FAA1
FB49
FBDE
FBDD
FB7C
FB2F
FAFB
FABB
FAEA
FC75
FF74
0286
0417
0428
0435
0537
065D
063E
04DB
03BD
0414
055E
062B
05D5
04ED
0446
0418
0439
049C
0531
0595
055D
04A9
0419
041D
048F
04FB
051D
04F5
0496
041D
03D2
0414
04FD
0603
0632
04CB
01EB
FEA4
FC57
FB8C
FB75
FADF
F9BE
F948
FA52
FBF9
FC78
FB49
F9CA
F992
FA9C
FB8F
FB8A
FB01
FAB9
FAC4
FADA
FB1C
FBCD
FC84
FC64
FB49
FA35
FA32
FB1D
FBE8
FBE4
FB5C
FADD
FA7C
FA1B
FA1D
FB37
FD82
0031
0259
03CC
04F3
05FD
0677
05EB
04A7
03B3
03E3
0501
0611
0645
05A5
04D0
0459
046E
04DE
0549
054C
04C7
0410
03C4
0436
0509
058A
056A
0504
04D3
04E1
04EB
04E5
0517
059D
05F4
0538
02F7
FFD1
FD1F
FBD0
FB93
FB55
FA94
F9F8
FA67
FBA2
FC56
FB9A
FA25
F97E
FA38
FB62
FBDE
FB98
FB3A
FB15
FAFC
FAE5
FB1B
FB9F
FBDC
FB56
FA68
F9F4
FA5B
FB1F
FB9A
FBA5
FB65
FAE6
FA4E
FA2F
FB24
FD0E
FF1F
00C4
023B
03F9
05C3
06B2
063B
04EB
03ED
03F6
04C0
057C
0590
04F3
041C
03AC
0404
04F4
05D2
05F7
054D
045F
03E6
0438
0509
05B4
05BF
053F
04B9
0499
04C8
04D5
049B
047C
04D8
0540
04A6
0285
FFA6
FD64
FC35
FB6F
FA7E
F9DF
FA5A
FBA3
FC56
FB9D
FA47
F9DB
FABF
FBEA
FC46
FBD8
FB51
FB0D
FAF1
FAFC
FB50
FBBD
FBC9
FB4E
FAC5
FAAE
FAF9
FB41
FB6E
FBB1
FBE6
FB81
FA6C
F990
FA01
FBD2
FE0F
FFE4
0169
0320
0502
064D
063E
04F3
0379
02F5
03B6
0508
05DD
05BA
0503
0471
0458
0481
04A3
04AD
0496
0442
03CE
03B3
0444
0520
057F
0521
049E
0495
04DD
04D3
0465
0452
0518
05FF
05A7
0390
00AF
FE51
FCC9
FB89
FA59
F9E0
FAB6
FC40
FD10
FC69
FB16
FA70
FAD7
FB84
FBAD
FB62
FB23
FB17
FB18
FB2B
FB7D
FBF2
FC1E
FBDB
FB87
FB80
FB97
FB6A
FB1B
FB3A
FBD0
FC0E
FB4C
FA16
F9B8
FAD1
FCC2
FE91
000B
01BD
03F8
0610
06D0
05C4
03DE
02C5
0352
04D4
05D7
0596
0498
03E6
03E5
0440
04A1
0502
053E
04F7
0439
03C5
042A
04EF
051C
048C
041C
046B
04E2
0497
03C4
03AB
04D8
062F
0624
0476
0230
002E
FE50
FC41
FA6A
F9AD
FA50
FB86
FC2D
FBE0
FB31
FAE5
FB2E
FB9D
FBBD
FB87
FB4D
FB52
FB8B
FBB9
FBB1
FB7C
FB3E
FB20
FB3F
FB81
FB8C
FB1F
FA90
FA9A
FB7E
FC7E
FC8A
FB77
FA49
FA31
FB73
FD61
FF4E
0130
0341
053E
0657
0604
04BF
03B0
03AC
047E
053E
054A
04D0
0462
0440
044A
0471
04C7
0517
04EC
0440
03BF
03FF
04B2
050D
04E8
04DF
053E
0554
046D
0329
030C
0487
0629
063A
04A0
029D
0102
FF6A
FD47
FAFC
F99B
F9B5
FAC8
FBD3
FC29
FBCC
FB31
FAE3
FB1C
FB93
FBB9
FB5A
FADE
FAC8
FB20
FB82
FBA0
FB7E
FB56
FB5C
FB98
FBCE
FBAB
FB39
FAF7
FB52
FC04
FC43
FBA4
FAB3
FA64
FB10
FC57
FDE4
FFE0
025A
04B0
0600
060C
0564
04C1
0479
0488
04C6
04FF
04FC
04B9
0474
046E
049E
04BF
04AE
0498
04B1
04E1
04E5
0498
041D
03D2
0414
04D9
0575
0520
03F5
031B
0398
050D
05FB
0559
0395
01D2
0079
FEF1
FCC5
FA8E
F96B
F9C5
FAEE
FBD6
FBEC
FB62
FAD8
FAD0
FB42
FBB3
FBC0
FB7F
FB4B
FB4F
FB65
FB62
FB5A
FB79
FBB6
FBD1
FB9F
FB3B
FAE1
FACD
FB2B
FBEC
FC8D
FC6F
FB8E
FAB7
FABE
FBB0
FD0B
FE9E
00B6
034B
057B
063B
058F
0499
045D
04C9
0523
050E
04CA
0499
0470
043F
0435
0476
04C9
04D7
049E
047D
04A3
04C1
047C
040E
0420
04EC
05BC
0594
0461
033C
035B
04BC
060C
05F5
046F
028D
0124
FFEB
FE1A
FBB2
F9C5
F960
FA69
FBB7
FC39
FBD7
FB35
FAE5
FAF1
FB1E
FB44
FB63
FB7A
FB7F
FB6C
FB4E
FB39
FB37
FB51
FB7B
FB8A
FB4A
FAC6
FA6F
FABF
FBA3
FC5B
FC33
FB50
FA97
FAB2
FB72
FC4F
FD52
FF1F
01E9
04C0
0642
05FE
04DF
0427
0440
04B2
04F4
04F8
04F1
04F0
04E5
04D2
04CA
04CD
04C4
04B8
04C9
04FB
0516
04E8
0493
0479
04CD
0554
058F
052B
045F
03D0
0405
04D7
057B
053B
0415
028A
00F2
FF29
FD09
FB04
F9EB
FA18
FAF7
FB9B
FB98
FB37
FAEC
FADD
FAEA
FAF5
FB0C
FB45
FB87
FB86
FB14
FA73
FA34
FAAB
FB83
FBFD
FBAE
FAE9
FA66
FA8B
FB24
FBBA
FBEC
FB93
FADF
FA66
FABB
FBCA
FCF1
FDFB
FF95
0257
056C
0700
063F
047C
03CD
04AC
05AE
0598
04DD
04A6
050B
051B
0478
03F6
0467
056B
05E9
057D
04D0
0491
04A3
0494
0479
04C3
055F
0597
04FC
0414
03D5
0486
057B
05CD
0533
03F2
023B
FFF3
FD47
FB11
FA2A
FA70
FAE2
FAD2
FAA0
FAF2
FB95
FBA8
FAE3
FA27
FA65
FB55
FBD4
FB67
FAC2
FAB2
FB1A
FB64
FB76
FB93
FB96
FB0F
FA20
F9B4
FA6C
FBB5
FC5E
FBFB
FB48
FB11
FB40
FB54
FB67
FC43
FE6F
0180
0461
0616
0651
059A
04E4
04D9
0561
05DB
05CA
053F
04A9
0466
0480
04CB
0515
053B
0533
0511
04F2
04CC
0486
043D
043D
049A
0503
052D
0526
051D
0508
04C5
047A
0475
04B0
04C2
0481
0459
04AE
04EB
03CB
00C3
FCE2
F9FC
F90D
F9AC
FAC2
FB71
FB5A
FAA0
F9DE
F9D5
FAC1
FBEF
FC4F
FB8B
FA76
FA2F
FAE6
FBB8
FBC9
FB35
FAC7
FAEE
FB57
FB7D
FB56
FB34
FB32
FB18
FADD
FAE6
FB6B
FBEE
FBC6
FB15
FAB4
FAFB
FB47
FB1E
FB4E
FD2D
00BA
0437
05E7
05CD
053F
051E
052D
050F
0509
055C
0590
0511
0441
0418
04CB
0577
054C
049E
0457
04B6
0515
04EF
0491
0488
04D0
04F7
04DC
04C4
04CF
04C5
048C
046B
04A4
04F8
04E6
0466
0424
04AF
057F
051B
0281
FE5E
FAAD
F914
F994
FAD2
FB79
FB3B
FAA4
FA54
FA82
FB10
FBB2
FBF9
FB94
FAB6
FA11
FA2D
FAD8
FB6A
FB7D
FB42
FB15
FB12
FB20
FB39
FB60
FB75
FB3D
FACD
FA99
FAF0
FB8C
FBD2
FB94
FB3C
FB2B
FB31
FAF8
FAE0
FBFC
FEEF
02D9
05C9
0684
059B
04A9
0497
0500
052C
0506
04F2
0504
04F3
04B2
04A3
04FF
0568
0566
0515
04F4
0515
0508
04A2
0466
04C1
054C
054D
04B9
0447
0469
04C9
04E0
04C2
04D2
04F9
04C6
0451
0455
050B
0547
0386
FFC7
FBEB
F9F5
FA3B
FB61
FBEC
FB7F
FAC4
FA76
FAB7
FB2A
FB63
FB35
FAC4
FA6B
FA6E
FABF
FB0D
FB1F
FB03
FAF0
FB00
FB1C
FB24
FB21
FB32
FB4F
FB3F
FAF0
FAB1
FADE
FB5B
FBA0
FB68
FB21
FB54
FBC5
FBA7
FAE1
FAC5
FCD4
00CD
0485
0601
0567
047B
047B
0510
054D
0516
0506
0557
058E
0549
04D7
04A9
04B2
04A3
0490
04CB
0534
0541
04D4
0490
04FB
059B
058D
04CC
044D
049A
050B
04D2
0441
044F
0506
0556
04B8
0431
04E1
05F6
051F
0167
FCC8
FA38
FA7A
FBA4
FBAF
FAA4
F9F5
FA60
FB29
FB5B
FB00
FAD4
FB21
FB73
FB61
FB15
FAF3
FB03
FB01
FAD0
FAA5
FAAF
FADA
FAF8
FB01
FB0E
FB1E
FB17
FB08
FB23
FB5D
FB56
FAE9
FAA3
FB26
FC18
FC36
FB00
F9F1
FB47
FF60
03E3
0610
0598
0493
04B8
0590
05AC
04E5
0475
0511
05DF
05B1
04A5
03EB
0430
04EA
054D
054A
054C
0562
0541
04F2
04DB
0517
0536
04E1
0468
045B
04BB
0506
04F9
04DD
04E7
04C8
044C
0408
04BC
05E6
05A4
02BB
FE54
FB1F
FA8A
FB65
FB9A
FAA9
F9DD
FA41
FB3F
FB95
FB0D
FA91
FAC2
FB33
FB3A
FAE6
FAC2
FAE8
FAF8
FACB
FAB5
FAF3
FB3D
FB32
FAEB
FAD3
FB07
FB36
FB2A
FB11
FB1C
FB29
FB14
FB20
FB97
FC18
FBCC
FA9A
F9CB
FB0C
FE99
02BF
0551
05AC
0503
04D0
054C
0597
0527
048D
04AE
0586
061D
05B5
04B4
0422
047A
0533
058B
0551
04E3
04A0
04A3
04DE
052B
054C
0522
04D9
04C6
04F6
0516
04E6
0497
0473
0460
0415
03CB
0430
0542
05AB
03E3
0014
FC53
FAA2
FAFB
FBAA
FB63
FA89
FA3F
FABE
FB27
FAD1
FA35
FA3C
FAFF
FBA9
FB8C
FAE7
FA76
FA8B
FAD8
FAFF
FB03
FB11
FB2D
FB3E
FB4F
FB76
FB91
FB6D
FB28
FB21
FB63
FB84
FB4C
FB2D
FBA6
FC4A
FC16
FAFC
FA8F
FC81
0083
044A
05E4
0592
04F9
0502
0529
04CA
0446
0477
0562
0618
05DC
050A
0494
04DB
0562
0583
0523
04AD
0490
04DC
0545
0569
0516
047D
0415
0439
04D4
0567
057F
0516
0484
040F
03BA
038D
03DB
04CC
05AE
0517
023E
FE1A
FADD
F9FE
FAED
FBD8
FBA6
FACF
FA5F
FAA4
FB10
FB27
FAFB
FAD7
FACF
FACB
FAD1
FAF5
FB23
FB24
FAEF
FABC
FAC3
FAF8
FB30
FB5A
FB75
FB6B
FB38
FB15
FB47
FBB6
FBEA
FBA4
FB43
FB57
FBD7
FC07
FB72
FACF
FB8C
FE4E
020B
04ED
05FB
05BE
0553
052B
04FA
0496
046C
04E3
059B
05CA
053D
04A2
04AF
053E
0596
0557
04D4
0485
047E
0494
04BF
0509
053F
0511
0494
044C
0487
04F1
050A
04CD
0494
0476
043A
03F7
0438
0515
0564
039F
FFC5
FBEA
FA4D
FB0D
FC31
FBFD
FAB6
F9E5
FA4B
FB1F
FB53
FADC
FA7D
FA95
FACB
FAC7
FABC
FAFE
FB62
FB73
FB28
FAF7
FB25
FB65
FB51
FB08
FAF1
FB19
FB26
FAFA
FAF8
FB6D
FBF6
FBF2
FB6E
FB20
FB64
FBB1
FB81
FB77
FCEA
0033
03DB
05F1
05F4
0514
04A8
04DD
0515
0508
050A
054B
0576
053B
04D8
04C7
050D
0538
0507
04C6
04C8
04ED
04DD
04A5
04A7
04F6
0525
04E2
047F
048E
050F
0569
0534
04B6
0464
0438
03FD
03EA
046D
0526
04AF
0206
FE06
FAEC
FA24
FAF4
FB8E
FB20
FA5F
FA3B
FAAC
FB09
FB0F
FB0C
FB2E
FB36
FAFD
FAD3
FB0E
FB6E
FB67
FAEC
FA91
FAC3
FB3D
FB6D
FB36
FAF1
FADC
FADA
FADA
FB10
FB87
FBD4
FB97
FB2A
FB50
FC18
FC87
FBDF
FAF6
FBAA
FEC3
02C9
055F
05A7
04DC
049D
0528
058D
0538
04AD
04AE
052E
057B
0537
04B8
0479
048D
04BD
04ED
051B
051F
04CF
045E
044F
04D1
0568
057C
0517
04C9
04E2
050C
04DA
0465
0414
03FE
03E7
03D5
0432
04FF
0534
038A
0005
FC4E
FA44
FA46
FB1F
FB85
FB49
FAFD
FAF1
FAE2
FA9B
FA63
FA97
FB18
FB64
FB3F
FAF8
FAF3
FB30
FB65
FB69
FB56
FB49
FB39
FB1F
FB1A
FB39
FB4B
FB1B
FACE
FACD
FB3A
FBB7
FBE0
FBCB
FBCC
FBD5
FB7F
FAE5
FB1B
FD3B
00FC
0486
0618
05AD
04BE
0492
0517
0573
0549
0508
051C
054E
052B
04BF
0488
04C6
051E
051A
04C1
048A
04B9
0517
053C
0508
04B2
0480
0497
04E7
0536
053A
04D9
0460
043C
0475
0493
0445
03FA
0459
0517
04BC
021E
FDFC
FAAB
F9D2
FAD6
FBB6
FB58
FA70
FA34
FABD
FB21
FADE
FA78
FA9E
FB27
FB5C
FB01
FA9C
FAAE
FB12
FB53
FB53
FB50
FB61
FB52
FB0B
FACB
FAD1
FAFE
FB18
FB2B
FB6E
FBC6
FBCB
FB65
FB07
FB13
FB38
FB01
FAE2
FC25
FF5A
0336
0595
05A9
04B5
0468
0509
0594
056B
0513
0541
05B3
059F
04ED
046D
04B0
053F
0543
04AF
043F
046F
04EB
051F
04FE
04D9
04D4
04CD
04CE
050D
056E
056E
04DB
0449
046D
0511
054D
04CB
044D
0475
0479
02D5
FF5C
FBE5
FA6F
FAF1
FB9F
FB31
FA3A
FA00
FAB0
FB50
FB32
FAC2
FAB1
FAF0
FAFE
FAD0
FAE3
FB5C
FBBE
FB9A
FB31
FB0C
FB2F
FB28
FAD7
FAA4
FAD9
FB2C
FB39
FB2D
FB6E
FBD2
FBC1
FB2B
FAD9
FB4C
FBD1
FB5C
FA53
FAA2
FD91
01F0
051A
05BD
04F7
04A7
053D
05BC
057A
0504
0526
05B5
05E1
0566
04D0
04A0
04AE
0494
0461
046C
04B7
04EB
04E7
04F4
053A
055C
04FA
0455
0418
0474
04E4
04E6
04A2
048A
04AB
04B0
0492
04B4
0525
054B
04B6
03FC
0412
04C0
0461
01B7
FDA9
FA97
F9E5
FAB2
FB34
FAD2
FA61
FA9C
FB24
FB3A
FADB
FAAA
FAEE
FB39
FB19
FABB
FA8E
FAA3
FABC
FAD4
FB1F
FB99
FBE0
FBB9
FB6E
FB6A
FB9E
FBA4
FB61
FB31
FB51
FB78
FB4B
FAEE
FACF
FAFE
FB22
FB1C
FB3F
FBA4
FBBF
FB21
FA8F
FBA6
FF01
0326
05C8
060C
0523
04AD
0507
0569
0549
04FB
04FD
0530
0521
04C2
047E
0493
04C5
04C6
04A2
0496
04AD
04B2
048A
045D
0459
0487
04D3
0524
054F
0520
04A4
0444
0461
04D2
0509
04CD
0486
049F
04D8
049B
03F9
03C8
046E
04EA
03A0
0042
FC7B
FA60
FA6A
FB47
FB8D
FB20
FACD
FAFE
FB4D
FB44
FB01
FAEE
FB22
FB54
FB54
FB41
FB3F
FB3F
FB2D
FB24
FB42
FB6E
FB74
FB51
FB32
FB2B
FB21
FB0C
FB13
FB46
FB6B
FB4A
FB19
FB41
FBAD
FBC9
FB59
FB04
FB78
FC44
FC34
FB08
FA5D
FC1F
0030
0431
05EB
0570
048F
0488
0500
0511
04AF
0485
04D7
0526
04F5
046F
0414
0412
0444
0490
04F4
053E
0528
04BF
0476
0496
04E8
0508
04F5
04F4
050B
04F4
04A8
048F
04DB
050D
049A
03D5
03B9
048C
055D
0533
0476
0469
0533
0534
02D4
FEAE
FB3B
FA3F
FB1F
FBF6
FBCA
FB32
FB09
FB3D
FB38
FAE3
FABD
FB08
FB60
FB55
FB05
FAE2
FB0D
FB3C
FB37
FB16
FB03
FAFA
FAF4
FB0A
FB49
FB77
FB59
FB18
FB23
FB86
FBBF
FB6A
FAE3
FAD5
FB44
FB81
FB34
FAE5
FB23
FB84
FB27
FA52
FABC
FDAF
0221
056C
060A
0500
045B
04D0
0566
0538
04A5
048F
0503
054B
0509
04B1
04BF
0501
0502
04C9
04B9
04E6
04F4
04B6
0475
0480
04AE
04A9
0478
0476
04B8
04F0
04F8
050E
0556
0579
0521
049D
0489
04DD
04DA
0437
03CF
0478
0569
0499
0122
FCBB
FA25
FA50
FB97
FBE9
FB02
FA2F
FA62
FB24
FB85
FB58
FB26
FB3E
FB58
FB2E
FAE9
FAD8
FAFD
FB1E
FB25
FB2E
FB46
FB54
FB47
FB38
FB3D
FB46
FB47
FB56
FB7E
FB85
FB37
FACD
FAD3
FB68
FBEC
FBBF
FB1D
FAE5
FB5E
FBB9
FB3E
FAA6
FBAB
FF01
032B
05CD
0600
04F9
0465
04AC
0509
04ED
04AE
04CD
052D
054D
0510
04D5
04DD
04EE
04C2
047C
0472
04B4
0500
051D
0509
04D5
0487
0441
0442
0492
04D7
04B9
0461
0445
047A
0497
0463
0441
049A
051E
051B
0498
0477
0524
0586
03F4
0042
FC4E
FA2D
FA28
FAE4
FB2B
FAFB
FAE2
FAF7
FAEA
FAB9
FAC7
FB30
FB88
FB73
FB28
FB19
FB4D
FB69
FB41
FB10
FB0E
FB24
FB2E
FB48
FB93
FBD8
FBBB
FB45
FAF0
FB05
FB48
FB60
FB63
FB8D
FBB0
FB5F
FAB7
FA83
FB29
FBE6
FB9E
FA8F
FA80
FCE0
00ED
044C
056A
04E1
0461
04B6
054D
0568
0521
050A
0540
0554
04FF
048D
0466
048F
04BE
04D0
04DB
04ED
04EF
04D9
04CB
04D3
04CA
0499
047A
04AD
0511
0533
04EC
0498
0490
04A4
0473
0427
0453
0503
056F
0503
045C
0495
0585
0566
02C3
FE77
FB0E
FA26
FAF3
FB94
FB48
FAC6
FAC4
FAFC
FAD7
FA6E
FA58
FAB8
FB12
FB15
FB05
FB31
FB62
FB3A
FADC
FABC
FAED
FB10
FAF5
FAF3
FB4C
FBAE
FB98
FB2E
FB10
FB66
FB96
FB39
FAC8
FAF1
FB82
FB9F
FB13
FAB1
FB16
FBA1
FB53
FA90
FB21
FE1D
0248
0538
05CE
0512
049C
04E0
0545
055F
056A
059E
05AF
0550
04C2
048D
04BE
04E7
04CE
04BB
04F7
054F
0563
0534
0518
0529
0517
04B4
0450
045B
04C1
0506
04F2
04D1
04E8
0508
04E1
0491
047D
04A5
049C
044D
0451
0503
057D
0425
0096
FC83
FA37
FA44
FB2E
FB5B
FAC7
FA87
FB0C
FB9B
FB6D
FABD
FA5E
FA99
FAFD
FB23
FB28
FB3F
FB44
FB0C
FACD
FAE0
FB2E
FB46
FB0E
FAF2
FB43
FBA8
FB93
FB14
FAC7
FAF6
FB3D
FB2C
FAE8
FAD7
FAF6
FAFD
FB04
FB66
FBFB
FBF8
FB1C
FAA8
FC51
0026
040F
05DD
057C
04A8
04B2
0544
0565
04F7
04BB
0517
058B
057A
04F6
048B
047B
049F
04CD
0509
0540
0539
04EA
04A1
049F
04BB
04A4
0465
045E
04AD
04FC
04F7
04CB
04DB
0523
053F
0509
04CE
04C6
04AE
0442
03E4
0443
052C
0531
0304
FF20
FB97
FA25
FA97
FB62
FB72
FB04
FADD
FB1B
FB3F
FB01
FABA
FAD5
FB34
FB65
FB3C
FAFF
FAF5
FB18
FB37
FB41
FB3E
FB2F
FB16
FB10
FB36
FB65
FB56
FB07
FAD2
FB01
FB65
FB94
FB7A
FB5E
FB5A
FB2E
FAC2
FA86
FADD
FB5A
FB34
FA94
FAF5
FD97
01BB
050E
0600
0540
04A0
04EB
0562
0528
0479
042B
0480
04F2
0510
04FA
04F7
04F6
04CA
0495
0494
04B5
04B4
0491
0497
04DD
050E
04EA
04B2
04C9
050E
0505
049F
046B
04C9
0551
0563
0511
04F5
052B
051A
0476
03FA
047A
055B
04CB
01CA
FD9E
FAB2
FA27
FAF2
FB67
FB08
FA90
FAA4
FB0E
FB42
FB28
FB13
FB2B
FB44
FB3A
FB28
FB31
FB43
FB3E
FB2C
FB27
FB2D
FB20
FB08
FB0D
FB37
FB51
FB39
FB1F
FB48
FB93
FB94
FB24
FAAD
FA9E
FAD7
FAE8
FACE
FB07
FBB2
FC16
FB8B
FAC0
FB79
FE9D
02D3
05A5
05F9
04F7
046C
04D0
053E
050B
04A0
04B2
052F
056F
0532
04E2
04DF
04FE
04F1
04D1
04E9
0527
052F
04E9
04A1
0494
049F
0494
0497
04D9
0521
0506
0497
0463
04AA
04F5
04C7
0465
0473
04E9
050D
0493
043F
04BF
054A
041E
00AD
FCA4
FA50
FA44
FB20
FB6B
FB1A
FAFC
FB53
FB8F
FB46
FAC9
FA9C
FABD
FACE
FAB2
FAAB
FADD
FB12
FB16
FAFF
FAFF
FB0F
FB09
FAF2
FAF7
FB1C
FB2A
FB07
FAEB
FB16
FB69
FB93
FB7F
FB6B
FB75
FB6C
FB2B
FAFA
FB2E
FB87
FB5A
FA9D
FA7C
FC54
000C
03CE
05B0
057E
04A6
0473
04DD
0516
04DD
04B9
050E
057D
0572
04F7
04A3
04C2
0505
050F
0502
0531
0589
05A2
0553
04EC
04C2
04CA
04C4
04B3
04C9
04FF
050C
04D3
0497
049C
04CD
04EB
04E3
04C3
0481
0422
0415
04D2
05E2
05BA
032B
FF06
FBAE
FAC2
FB82
FBF7
FB44
FA5B
FA60
FB2A
FBAD
FB6E
FAF7
FADB
FAF4
FAD7
FA99
FAA7
FB0C
FB52
FB2E
FADE
FAC3
FAD7
FADA
FAC1
FAC8
FB02
FB31
FB29
FB0F
FB1A
FB38
FB37
FB20
FB2A
FB52
FB55
FB1D
FAF4
FB1E
FB63
FB5D
FB1B
FB21
FB8F
FBBB
FB0F
FA3A
FAE3
FDE0
01FF
04FD
05AE
04EE
0469
04D0
057F
05AB
055F
052B
0543
0559
0534
050A
051C
0548
0539
04ED
04BD
04DC
050E
0508
04DE
04DE
0519
054D
054E
053F
0545
053D
04F6
0494
0473
04A2
04D1
04C0
0498
04A0
04CB
04DA
04D2
04F0
0521
0501
0491
0483
053C
05C7
0476
00D8
FCAA
FA41
FA3B
FB26
FB6B
FAEE
FA8D
FAA8
FACC
FAAB
FA97
FAE8
FB53
FB53
FAF6
FAD0
FB20
FB78
FB5F
FAFC
FACA
FAEA
FB18
FB2E
FB4E
FB86
FB96
FB4B
FAE3
FACF
FB1B
FB6C
FB78
FB5B
FB54
FB5D
FB51
FB41
FB58
FB76
FB43
FAC1
FA81
FAF2
FB9F
FBA2
FAF1
FADF
FCDD
00B2
046A
0631
0605
055A
0545
0587
0569
04F0
04C7
052D
0590
0560
04D9
04A5
04E9
0520
04ED
049C
049C
04CE
04C0
045F
041B
044B
04C1
0515
052F
0536
0532
0501
04AA
0474
0483
04AA
04B3
04B3
04CC
04DC
04AD
0469
0476
04D9
0508
04AD
0449
048F
0521
0486
01C5
FDD2
FAD9
FA18
FACD
FB5A
FB1E
FABB
FAE0
FB51
FB64
FB00
FAB7
FAE9
FB4C
FB6E
FB53
FB5F
FBAD
FBDE
FB9B
FB0E
FAAC
FAAE
FAEE
FB27
FB39
FB28
FB0F
FB10
FB44
FB8B
FB9F
FB67
FB31
FB52
FBAE
FBD3
FB99
FB5C
FB65
FB78
FB42
FB03
FB49
FBFA
FC22
FB3B
FA58
FB57
FEBE
02D7
055A
05AA
050B
04DB
0532
055B
0517
04D7
04EA
0504
04C1
044B
0428
0482
04FA
0524
04FA
04BB
049D
04B0
04E3
0513
0512
04D3
0487
0474
0499
04B4
0496
0471
0490
04E5
050D
04D0
0473
0458
0476
0477
0448
0442
0499
04EF
04C2
044D
0469
0549
05A9
03E8
000B
FC20
FA48
FA9F
FB74
FB6D
FAD4
FAB3
FB35
FB8F
FB49
FAE3
FAFB
FB5F
FB69
FB03
FABA
FAED
FB53
FB80
FB78
FB7D
FB8D
FB71
FB37
FB36
FB81
FBBD
FBA9
FB85
FBA1
FBD0
FBB0
FB5C
FB59
FBC3
FC0B
FBBA
FB28
FAFE
FB3A
FB38
FACD
FAAD
FB56
FC0C
FBB3
FA93
FA84
FCF0
0108
0466
057A
04DF
044A
0496
0541
0585
0551
051B
0518
0510
04D2
0484
046C
048F
04B2
04B1
04A6
04B2
04C1
04AB
0473
044D
0461
04A3
04EC
051B
0516
04D4
0474
043C
045B
04A7
04CA
04B1
04AA
04E7
051F
04ED
047E
046B
04D1
050D
04AE
0447
04B5
0590
0514
0218
FDC5
FAAD
FA29
FB23
FBB5
FB53
FAE0
FB0E
FB7C
FB85
FB31
FB00
FB15
FB15
FADF
FAC8
FB0D
FB60
FB57
FB04
FAD7
FAFC
FB3B
FB60
FB7B
FB9B
FBA0
FB7F
FB73
FBB6
FC08
FBEB
FB53
FAD6
FAF7
FB76
FBB3
FB87
FB5C
FB72
FB72
FB08
FA91
FAB8
FB6B
FBBC
FB27
FAA3
FBDC
FF3A
031C
0553
054A
0456
040E
04B1
055D
056B
051A
04F8
051A
052E
0514
0500
050D
050D
04D8
0495
0487
04AA
04C4
04B7
049A
0482
0470
046C
0496
04E5
0509
04C6
0457
0437
0482
04CC
04B9
047D
047E
04B3
04BF
0493
0499
0501
0551
0507
0480
04A8
0589
05B3
039F
FF9C
FBD3
FA36
FAB1
FB9E
FBB0
FB09
FA8A
FA8D
FAB9
FAB7
FAA7
FAC9
FB16
FB54
FB6D
FB76
FB71
FB50
FB26
FB26
FB5A
FB86
FB7A
FB5E
FB73
FBA9
FBAD
FB64
FB23
FB34
FB63
FB4D
FAFB
FAE2
FB33
FB88
FB7D
FB44
FB4B
FB85
FB73
FB06
FAE1
FB6C
FBFE
FB9E
FAA8
FAE4
FD95
01BB
04E3
05A1
04D3
044A
04BF
0576
0593
0522
04BF
04B4
04D6
04EF
04FB
04EF
04B5
0465
0447
047D
04C7
04D9
04C3
04D0
0510
0535
050A
04C1
04B0
04D7
04EE
04D7
04C8
04E8
0505
04E0
0490
046E
0493
04B8
04A8
0497
04CA
050E
04E6
045A
042B
04DA
0592
04AB
0179
FD63
FABC
FA80
FB86
FBF8
FB4B
FA6E
FA5C
FAF1
FB63
FB50
FB00
FAD3
FACE
FAD4
FAED
FB26
FB55
FB45
FB0B
FAEF
FAFD
FB00
FAE5
FAEA
FB3A
FB92
FB95
FB52
FB2A
FB45
FB5E
FB47
FB3A
FB77
FBC5
FBB3
FB50
FB23
FB5D
FB7D
FB24
FAC3
FB04
FBA3
FB94
FA9A
FA20
FBE1
FFC5
03B0
0598
0574
04D3
04EF
05A0
060F
05DD
0550
04D6
049E
04A8
04DC
0508
0501
04D3
04C1
04E7
0512
050E
04F8
0511
054E
0558
0507
04A1
0485
04AD
04C1
0491
0450
0440
0450
0445
0424
0437
0495
04EC
04E4
049C
0486
04BE
04D6
047F
042A
0496
058D
0590
033B
FF11
FB54
F9E5
FA81
FB5F
FB49
FAA7
FA78
FAE2
FB33
FB04
FAB6
FABE
FAFC
FB0F
FAFB
FB08
FB35
FB3A
FB04
FADD
FAF2
FB06
FAE2
FAC5
FB13
FBA0
FBCA
FB5A
FAD9
FAD4
FB1D
FB37
FB1E
FB40
FBAE
FBF4
FBCB
FB90
FBB3
FBF3
FBBE
FB2F
FB12
FBAB
FC1B
FB8F
FAB7
FB5A
FE48
0239
0501
05AB
0518
04B5
04FE
0573
0586
0543
050B
050C
0523
0511
04C9
047E
0477
04C7
052F
055E
0540
0509
04F7
050E
0524
0513
04E5
04C3
04C3
04D4
04DA
04CD
04B4
049E
048F
0487
048C
04A5
04BC
04AD
0478
0460
048E
04B9
0472
03E6
03DD
04AC
054D
0418
00A6
FC9E
FA39
FA0E
FACD
FB00
FA96
FA68
FAC9
FB32
FB2B
FAE8
FAD8
FB08
FB34
FB45
FB5B
FB67
FB33
FAC9
FA8C
FAAF
FAE1
FACF
FAAC
FAE3
FB67
FBB5
FB89
FB3D
FB3C
FB74
FB89
FB75
FB89
FBD6
FBF8
FBAE
FB4E
FB47
FB69
FB28
FA8D
FA58
FB02
FBE0
FBD7
FAEE
FAAD
FC94
0057
03F0
0598
055C
04AD
04AD
0536
0585
0558
0517
0522
054D
053A
04EE
04C3
04E2
0515
0523
0519
0517
050A
04D5
0492
0483
04B2
04E2
04E3
04CF
04CE
04D1
04AD
0471
045C
0473
0479
045C
045B
049C
04D6
04B6
046F
047F
04DE
04EA
0454
03D0
0441
054B
053B
02CF
FEC9
FB5C
FA05
FA58
FAE0
FACB
FA6D
FA6C
FAD6
FB33
FB37
FB18
FB2B
FB6C
FB94
FB7C
FB49
FB30
FB35
FB37
FB25
FB14
FB16
FB20
FB1C
FB0F
FB13
FB2B
FB47
FB64
FB87
FB9A
FB7A
FB38
FB14
FB22
FB26
FAF4
FACE
FB14
FBAE
FC11
FBF6
FBC6
FBE9
FBFD
FB60
FA8F
FB2B
FE28
0250
053B
05BE
04DA
044C
04A2
0523
0522
04CC
04A6
04C3
04E0
04E2
04E4
04EC
04E8
04E3
04F1
0501
04F0
04CD
04CE
04FB
051D
0508
04DD
04D9
04F7
04FD
04DD
04C9
04E1
04F4
04CF
048C
0461
045A
0461
0470
0486
048E
0479
0460
045D
0467
046C
0488
04DB
052A
04FF
0465
0429
04D8
0587
0477
0122
FD30
FACD
FA7E
FB08
FB36
FB02
FAF0
FB0E
FAFD
FAB1
FA8B
FAB5
FAE6
FAEA
FAFA
FB3B
FB66
FB3C
FAFD
FB0F
FB59
FB72
FB49
FB2F
FB46
FB47
FB01
FAB2
FAB3
FAEE
FB06
FAF0
FB04
FB5A
FB9C
FB9A
FB9C
FBCE
FBDD
FB78
FAED
FAC6
FB02
FB2B
FB12
FAFC
FB16
FB26
FB0E
FB28
FBA2
FBDF
FB3A
FA78
FB71
FED5
02F0
0565
05AA
051E
0500
0539
052B
04E5
04E9
053D
055D
051E
04EC
050A
0525
04EB
04A5
04B1
04DC
04C4
0488
049C
0502
0545
0528
04F1
04ED
04FD
04E1
04AC
04A4
04C9
04D1
04AF
04A7
04C6
04BE
0480
0479
04D6
051F
04ED
0496
04A4
04F1
04EC
048F
0475
04C9
04DF
044F
03E4
0484
0551
0429
006F
FC42
FA3D
FA97
FB72
FB7B
FB14
FB08
FB2F
FAF4
FA79
FA6D
FAEB
FB49
FB21
FADE
FAEA
FB03
FAD3
FAA5
FAE4
FB51
FB59
FB02
FAD9
FB0D
FB34
FB00
FAB7
FABB
FAED
FAEC
FAC1
FAD7
FB40
FB8E
FB81
FB67
FB7A
FB77
FB34
FB0F
FB57
FBB0
FB96
FB38
FB23
FB5E
FB68
FB30
FB56
FC04
FC44
FB51
FA56
FB94
FF85
03CA
05C8
0570
04B1
04BB
0508
04DB
0489
04C3
055D
0593
0533
04DE
04FB
0530
0517
04E8
04F0
04F9
04BB
047B
04A1
0505
0526
04F4
04D3
04E6
04E3
04A6
0484
04C1
050D
04ED
0484
0467
04B4
04EB
04D2
04DA
053F
0573
04FC
044C
0422
0472
049F
0483
0491
04DB
04C7
0429
03F6
04E6
05C8
0466
0063
FC29
FA3D
FA85
FB0B
FAC3
FA65
FAB4
FB3F
FB35
FABC
FAA2
FB18
FB72
FB44
FAF3
FAF4
FB0F
FAE5
FAA8
FABF
FB0C
FB24
FB05
FB09
FB47
FB7D
FB84
FB83
FB8A
FB6B
FB0E
FAB9
FAB9
FAE8
FAEF
FAE1
FB1F
FB8E
FB98
FB1E
FACD
FB1C
FB8B
FB73
FB0D
FB01
FB49
FB48
FAED
FAEE
FB84
FBBF
FAEF
FA45
FBDF
FFF0
0403
05B2
0541
04B4
0507
057A
0544
04D2
04E9
0560
0577
0507
04AE
04C4
04E5
04BB
0496
04D7
0534
052F
04E1
04BD
04D3
04CC
0497
0485
04BF
0504
050B
04E3
04CA
04C9
04C1
04BD
04E4
0516
0500
04B0
0493
04C5
04D9
0499
0474
04C4
0522
0503
049B
0490
04DB
04C7
0438
0421
050D
05AA
03ED
FFCB
FBC7
FA2E
FAA8
FB36
FAE2
FA76
FAC2
FB5D
FB78
FB1C
FAF4
FB2E
FB4F
FB15
FAE5
FB12
FB4D
FB31
FAE6
FACC
FAD2
FAB6
FA96
FAD4
FB61
FBBA
FB95
FB3B
FB14
FB22
FB27
FB1C
FB30
FB5B
FB59
FB1F
FAFB
FB16
FB35
FB2D
FB2F
FB5B
FB6F
FB3C
FB0D
FB3A
FB8B
FB88
FB4D
FB64
FBCB
FBB2
FAD2
FA87
FC94
00C1
0494
05F4
0556
04B6
0504
0580
0557
04D3
04B1
04F5
0510
04D2
04A5
04CF
0501
04ED
04BB
04B0
04B5
04A5
04AA
04F0
0531
0506
048F
0456
0490
04E7
0505
04FF
050B
050D
04CB
0469
0459
04B3
0509
050F
04F5
04F0
04D1
0472
041F
042B
0467
046F
044E
045C
0487
045C
03EA
03F5
04BF
04F4
02E0
FEC7
FB23
FA07
FAE7
FBAA
FB52
FAB0
FAB5
FB1D
FB1D
FAB4
FA96
FB0A
FB89
FB92
FB54
FB3F
FB57
FB67
FB70
FB8D
FB9A
FB67
FB1E
FB15
FB4B
FB6F
FB5E
FB49
FB53
FB55
FB25
FAEF
FAFF
FB45
FB67
FB45
FB23
FB2F
FB48
FB56
FB8A
FBEC
FC27
FBFD
FBAF
FB8D
FB74
FB20
FAD6
FB16
FBA8
FB9F
FACE
FAB5
FD06
0144
04D7
05D9
050E
0486
04FE
057F
0545
04CD
04E1
0557
0569
04E7
0471
0477
04AF
04B4
049E
04B3
04D8
04D1
04B9
04CD
04F5
04EB
04BD
04B3
04CF
04C8
048B
046B
04A7
0500
0508
04C5
04A2
04C5
04E5
04D3
04C3
04DB
04DE
049E
045D
0463
0488
048B
0491
04DB
051E
04D5
0434
0426
04D7
04D3
027F
FE63
FB0C
FA40
FB1E
FB99
FB11
FA93
FADF
FB61
FB44
FAB4
FA81
FADF
FB34
FB15
FAD5
FAE5
FB26
FB37
FB1B
FB1A
FB3D
FB52
FB4E
FB49
FB3C
FB18
FAFA
FB0E
FB3E
FB49
FB1C
FAF5
FB03
FB22
FB1A
FB06
FB20
FB52
FB4E
FB20
FB28
FB6D
FB80
FB3B
FB1B
FB6E
FBB9
FB7B
FB16
FB44
FBC6
FB8B
FA8D
FA9C
FD6B
0209
0577
05FA
04DD
0466
0503
0575
0518
04B4
050A
05A5
05A8
051D
04C9
04F7
0520
04E0
0496
04B3
0502
050B
04D6
04C1
04D1
04BC
047F
046A
049D
04DA
04E5
04D3
04D9
04F5
0503
04FF
0507
051E
0522
050D
0500
04F9
04D8
04B0
04BE
04EA
04D0
0473
0464
04D4
0518
049E
040C
047E
059E
0556
0233
FD8A
FA5C
FA04
FB03
FB48
FAB1
FA77
FB02
FB73
FB2B
FAAF
FAC2
FB48
FB99
FB81
FB60
FB6D
FB6A
FB31
FB0D
FB32
FB58
FB38
FB0B
FB2B
FB75
FB8A
FB68
FB5B
FB6B
FB53
FB02
FAC6
FADB
FB0A
FAFE
FAC4
FAB0
FAD6
FAF1
FAE3
FAE5
FB0C
FB27
FB29
FB56
FBAD
FBC3
FB7A
FB67
FBE5
FC37
FB73
FA43
FACD
FE39
02D6
05A8
05A7
0494
046C
0519
0552
04D1
0488
04FA
057B
0552
04C4
048B
04C3
04E6
04B6
0491
04C3
0501
04EE
04A7
0482
047D
0463
043A
043A
0464
0490
04B8
04F0
0520
051C
04F5
04F5
0534
0568
0547
04F5
04CD
04D9
04CF
049C
047C
0482
0472
044A
0461
04BE
04D7
0476
0456
0523
0600
0500
016D
FD0F
FA7B
FA5B
FB21
FB47
FAF0
FAF2
FB40
FB26
FA97
FA4F
FAA8
FB1D
FB2A
FB06
FB2B
FB7E
FB78
FB0B
FAC9
FB0D
FB72
FB6E
FB19
FAEC
FB0D
FB38
FB3E
FB30
FB24
FB19
FB1E
FB40
FB5F
FB4A
FB0B
FAE7
FB06
FB34
FB33
FB1F
FB3E
FB7D
FB7B
FB2D
FAFF
FB2C
FB63
FB61
FB66
FBA5
FBAD
FB0A
FA6F
FB73
FEBE
02DF
0586
05DB
050C
04A2
04EA
0543
0558
0558
055E
0545
0511
0503
0525
052F
04FD
04DC
0519
0579
057A
050F
04BA
04D0
0506
04F1
04A2
0479
048D
04A3
0498
0486
0486
0493
04AC
04D4
04F8
04F5
04CF
04BD
04E4
0513
0511
04F9
0512
053A
0509
047D
0428
0455
048E
045D
042B
049E
0539
0460
0133
FD03
FA39
F9E4
FAD3
FB42
FACE
FA55
FA77
FAE5
FB11
FAEC
FACC
FAE0
FB0C
FB21
FB0A
FAD5
FAAB
FAB3
FAF5
FB41
FB57
FB2F
FB04
FB00
FB0E
FB11
FB18
FB30
FB3E
FB27
FB06
FB0B
FB37
FB65
FB80
FB89
FB70
FB29
FAD6
FAC0
FAFB
FB44
FB5C
FB6F
FBB7
FBFC
FBCA
FB4D
FB3B
FBBA
FBE2
FB06
FA2D
FB53
FF07
035A
05C6
05CC
0515
051F
05A8
05A8
0512
04CA
0535
05AD
0588
04FF
04BB
04E0
04FD
04D1
04A7
04CF
0517
0522
04F3
04DD
04F8
0508
04E5
04BB
04B9
04CD
04C2
049B
048F
04BE
04FD
0510
04F1
04CE
04BC
04A8
0488
047A
0490
049D
0473
0441
0472
0500
04F7
0329
FF91
FBD0
F9DA
FA13
FB15
FB62
FAF1
FABB
FB2B
FB96
FB4D
FAA1
FA6A
FAD5
FB3A
FB26
FAF2
FB18
FB6C
FB6E
FB1D
FAF8
FB34
FB71
FB58
FB27
FB49
FBA4
FBBA
FB6C
FB30
FB5D
FBB1
FBC2
FBA2
FBA5
FBCA
FBC2
FB7E
FB49
FB46
FB3A
FB06
FB05
FB7F
FBF5
FBA6
FADC
FB25
FDA4
0180
048E
0589
0522
04D3
0522
0577
054F
04F6
04F0
052F
053F
0500
04C7
04CF
04EA
04DF
04C7
04DE
0513
0511
04B9
0453
043A
0469
048F
0482
0468
0472
0493
04A2
049D
04A5
04C1
04CF
04BF
04AB
04A5
048F
044C
040E
0426
0481
04A1
0458
0440
04ED
05B5
04EC
01C1
FD93
FACB
FA6C
FB3D
FB7E
FAEB
FA84
FACE
FB1D
FAC7
FA3C
FA54
FB05
FB73
FB38
FAEC
FB31
FBBE
FBDD
FB81
FB4F
FB92
FBD0
FB94
FB2F
FB35
FB99
FBCD
FB98
FB58
FB51
FB4C
FB0D
FADC
FB24
FBB1
FBE5
FB9E
FB6F
FBBA
FC09
FBCA
FB4C
FB5E
FBFD
FC24
FB53
FABD
FC31
FFD9
03AF
0587
053A
046E
0475
050E
0544
04EB
04AF
04F5
0550
0531
04BA
0485
04C5
050B
04F2
04AB
04A3
04DC
04F5
04C2
0488
048F
04BB
04C9
04BE
04D1
04FC
04F6
04A8
0465
047C
04BD
04C1
048C
0483
04BF
04D5
0486
043C
046E
04DD
04DB
0470
046E
0511
050D
02CC
FE9B
FADD
F99D
FA78
FB67
FB3C
FA9C
FA9C
FB2F
FB7B
FB34
FAED
FB19
FB66
FB5A
FB15
FB13
FB5E
FB80
FB3F
FAE2
FABF
FAC8
FACD
FADD
FB28
FB89
FB9E
FB52
FB08
FB1F
FB6F
FB91
FB73
FB58
FB5A
FB45
FB03
FAE0
FB20
FB86
FB99
FB59
FB4F
FBB5
FBF9
FB7E
FAC6
FB5D
FE2F
0241
055E
0637
0574
04B9
04D3
053D
0537
04D3
04AE
04FE
0554
0546
04FB
04D4
04DC
04D8
04B9
04B9
04F6
0538
0540
0523
0520
053B
053B
0512
04F1
04F3
04E3
0496
0442
043F
0488
04C3
04C4
04B9
04C4
04B2
045C
0414
044B
04D4
0500
04A9
048C
052E
05AA
0458
00D4
FCD1
FA85
FA77
FB48
FB83
FB16
FAD0
FB05
FB43
FB21
FACE
FAA5
FAA6
FA9A
FA8B
FAB5
FB1A
FB70
FB7B
FB5B
FB45
FB35
FB09
FAD5
FAD2
FAFD
FB16
FAFA
FADF
FB04
FB50
FB70
FB4B
FB22
FB2E
FB51
FB54
FB4E
FB7F
FBD5
FBE9
FB94
FB49
FB7A
FBD3
FB85
FA8A
FA3E
FC29
001A
03FB
05BD
055A
047C
0476
0508
0540
04EF
04BE
050C
0561
0534
04C0
04A5
04FB
053B
0511
04D0
04DF
0518
0519
04EB
04F3
053F
0566
0524
04CD
04D5
051D
0526
04D0
0489
04A0
04D8
04D8
04BE
04D7
0505
04E6
0485
046C
04CF
0521
04DF
047E
04E3
05D5
05A3
02EA
FE80
FAED
F9E6
FAC1
FB93
FB64
FAD2
FAC3
FB29
FB4C
FAF7
FAB2
FAEE
FB66
FB91
FB5D
FB37
FB5F
FB97
FB8D
FB50
FB2C
FB34
FB33
FB0C
FAEB
FB01
FB2E
FB2C
FAF2
FAC4
FAD2
FB02
FB24
FB2D
FB26
FB06
FAD5
FAC5
FAFE
FB48
FB3E
FAE1
FABA
FB1B
FB7E
FB36
FAB4
FB87
FE96
02AF
0576
05C7
04C0
043D
04C9
0579
057D
0524
0524
057C
0594
0533
04CA
04BA
04D5
04BA
0472
0450
046B
0487
047C
0473
048F
04AB
049A
0480
049F
04EC
051B
0512
0506
0518
0515
04D8
04AA
04EB
056D
058A
0506
0478
0480
04DE
04D2
0452
0442
0511
059F
042A
0076
FC74
FA63
FA93
FB70
FB86
FAED
FA9D
FAE4
FB2C
FAFD
FAA3
FA9B
FADA
FAFB
FAEF
FB0A
FB6A
FBAF
FB89
FB31
FB1D
FB5B
FB92
FB91
FB8C
FBA4
FBA4
FB61
FB28
FB63
FBEF
FC2F
FBDF
FB75
FB75
FBB0
FB98
FB29
FAFC
FB50
FB93
FB38
FAA8
FABF
FB6C
FBA5
FB02
FAD0
FCC4
00B5
045E
05B7
0505
042E
0459
04F8
0511
04B3
04A2
050C
054E
0505
04A0
04AE
04FF
04F9
0489
043D
046A
04B6
04AE
0470
045F
0474
044E
03EE
03E0
046B
050B
050F
048D
043A
0469
04A7
047E
042C
0431
047A
047F
042F
041B
048E
04F7
04C6
046E
04D6
05BC
056D
02A5
FE62
FB22
FA56
FB1D
FBAD
FB69
FB0B
FB2F
FB7D
FB68
FB19
FB1F
FB83
FBBA
FB78
FB20
FB25
FB6B
FB81
FB63
FB70
FBCA
FC0C
FBE1
FB86
FB70
FBA3
FBB6
FB79
FB3B
FB4C
FB7E
FB72
FB2E
FB0E
FB30
FB46
FB23
FB11
FB5C
FBC0
FBBC
FB64
FB61
FBE2
FC18
FB59
FA7D
FB69
FED8
0322
05BE
05D6
04D5
046C
04BF
04E1
0476
0424
046B
04E2
04E8
049D
049A
04F0
04FE
0473
03DD
03E7
046D
04C2
04AC
0496
04C8
04F8
04CC
047C
047E
04C9
04E5
04B1
049B
04E9
0537
050C
04A1
0492
04EB
0515
04C4
047D
04C4
0533
04FE
044A
0431
051B
059F
03DB
FFD0
FBBF
F9E9
FA5E
FB5B
FB7D
FAF7
FAB7
FAFF
FB55
FB6E
FB8A
FBDE
FC1B
FBDA
FB48
FAFA
FB2E
FB84
FB8D
FB56
FB35
FB48
FB56
FB41
FB35
FB58
FB89
FB8E
FB79
FB85
FBB4
FBC3
FB99
FB7A
FB9A
FBBD
FB87
FB12
FAD8
FB02
FB23
FAE7
FAB3
FB16
FBC6
FBD0
FB18
FB08
FD28
0115
0495
05D4
0531
0476
04AA
0540
0555
04F4
04C0
04E3
04EF
04B1
0488
04BE
0507
04EB
0478
042A
0439
0456
0441
042E
0465
04C4
04EE
04D7
04CA
04E5
04F2
04D0
04BC
04F4
053E
0529
04BC
0482
04C3
0512
04E4
045D
0427
046F
04A8
046A
0428
0485
0513
045D
0192
FDC0
FB01
FA62
FB08
FB73
FB25
FAC6
FAE6
FB43
FB54
FB17
FAF5
FB13
FB25
FAFC
FAD8
FB07
FB66
FB8B
FB60
FB35
FB40
FB52
FB31
FAFE
FAFC
FB26
FB36
FB1C
FB1A
FB52
FB82
FB5C
FB0C
FAFA
FB30
FB45
FB07
FAD6
FB15
FB8F
FBBC
FB94
FB8D
FBCA
FBC1
FB21
FACD
FC3D
FFB5
038C
05AF
05AA
04CE
0486
04EA
0534
0500
04B3
04BB
04F7
0507
04E4
04D7
04F5
0501
04D6
04A4
04A8
04D1
04E3
04D3
04D0
04F2
0515
0516
050B
051E
053D
052E
04E8
04A9
049D
04AF
04BA
04CE
0505
052E
04F8
047A
043F
0492
04F8
04CB
0433
040E
049E
04B6
02DB
FF28
FB96
FA0D
FA8F
FB8D
FBC7
FB58
FB01
FB05
FB13
FAFE
FAFC
FB28
FB3F
FB07
FAB3
FA9C
FAC6
FAF5
FB14
FB48
FB89
FB95
FB54
FB16
FB30
FB81
FB9F
FB73
FB4D
FB5E
FB69
FB3A
FB0F
FB32
FB6A
FB3F
FACE
FAD9
FBB4
FC85
FC36
FB13
FAF2
FD42
0149
04B7
05F5
0578
04CE
04D0
051B
0517
04DA
04E0
053A
0578
054A
04EC
04C8
04F2
0524
052E
051F
0510
04F5
04C4
0496
048D
049C
049D
0492
04A1
04CC
04DC
04AF
0478
0474
0489
0468
041F
0418
0471
04B0
0473
0427
048B
054C
04D2
01F4
FDAF
FA7E
F9D4
FAC6
FB6D
FB1B
FAA9
FADA
FB51
FB4A
FACE
FA8F
FAD9
FB31
FB1C
FAC9
FAA3
FAB1
FAAE
FA97
FAA9
FAED
FB1E
FB16
FB0B
FB2D
FB51
FB3C
FB16
FB33
FB80
FB89
FB2F
FAF7
FB4B
FBCE
FBDB
FB80
FB6D
FBD3
FBF5
FB3E
FA89
FB8E
FEE4
0303
05A7
05FE
0527
04AA
04F0
055B
0558
0501
04C7
04D6
050A
0534
054B
0558
0561
056F
0585
058C
0569
0523
04EF
04EC
04FD
04F2
04C9
04AB
04AA
04A3
047E
046A
0497
04DE
04D8
0474
042A
045E
04BD
04A1
0411
03EB
04A8
0546
0407
0074
FC45
F9D4
F9D6
FAF6
FB93
FB54
FAEA
FACC
FAC8
FAA5
FA89
FAA6
FACC
FABC
FA98
FAB1
FAF9
FB11
FAE4
FAD1
FB0E
FB3D
FAF9
FA89
FA8B
FB0F
FB76
FB52
FB02
FB11
FB5C
FB53
FAEC
FACA
FB33
FB90
FB58
FAFC
FB4D
FC11
FC18
FB0B
FA71
FC39
004A
0452
062A
05E5
0532
0531
0591
059A
0543
04FB
04E0
04C0
04A2
04CC
0536
0563
0510
04AA
04BA
0523
0549
04FA
04B1
04D6
051F
0506
049D
0471
04B7
04FC
04DD
04A1
04C3
0523
0531
04D3
0498
04D7
050E
04AC
0420
0471
058A
05AF
033F
FED1
FAEA
F97A
FA13
FAE0
FAD8
FA74
FA75
FAC2
FAD1
FA9F
FAA0
FAEA
FB0D
FAC9
FA8C
FAD1
FB63
FB9F
FB5F
FB1F
FB35
FB53
FB15
FAB4
FABC
FB38
FB94
FB71
FB1C
FB06
FB1C
FB09
FAE6
FB1A
FB93
FBAB
FB23
FAAD
FAFA
FB97
FB72
FAAE
FB0E
FDF9
026B
05A7
0621
04FB
045C
04ED
059C
057A
04EC
04CA
0515
0528
04DB
04C1
0527
0587
0550
04C2
048F
04E1
0532
0524
04F8
0505
0528
050D
04C9
04BD
04F2
04FF
04BE
0493
04CC
050D
04D5
0458
0442
04A1
04BA
042D
03C7
0473
057F
04DC
017C
FCF3
FA09
F9E2
FB15
FBA3
FB24
FA9F
FAD4
FB57
FB70
FB26
FB02
FB2E
FB4A
FB17
FAD8
FADF
FB12
FB1E
FAF6
FADB
FAF4
FB22
FB39
FB3B
FB32
FB14
FAEE
FAFB
FB58
FBB4
FB91
FAF4
FA7D
FAA9
FB31
FB74
FB60
FB75
FBDE
FBF8
FB4D
FABC
FBF1
FF6B
0385
05E8
05E3
04D9
046F
04D4
051E
04D1
0472
048E
04F0
050B
04DB
04D7
0527
055F
0529
04C5
04AB
04E4
0516
0515
0506
0501
04E9
04B9
04AB
04DA
04F5
04A6
0430
0432
04C5
053E
0514
049C
0479
04A6
0491
043B
0463
0545
0598
03B2
FFAE
FBBE
F9FB
FA53
FB13
FB14
FAB2
FAB3
FB07
FB17
FADF
FAF3
FB7E
FBDD
FB79
FAA8
FA43
FA94
FB22
FB6E
FB74
FB60
FB30
FADC
FAA1
FAC2
FB12
FB20
FAE1
FAD3
FB45
FBD6
FBF6
FBA8
FB6B
FB6B
FB56
FB0E
FB14
FBC0
FC66
FBFC
FAB6
FA69
FCAD
00DD
0482
05D4
0553
04BD
04F0
0555
052F
04BF
04BB
0531
057D
053F
04E0
04E8
053D
0555
0501
049B
047F
0496
04A8
04B5
04DF
050B
04FF
04C1
04A2
04C3
04E8
04DA
04BF
04D8
04FF
04D7
0476
045D
04AB
04C2
0428
037E
03D4
04FB
0515
0290
FE3A
FAB9
F9D2
FAC0
FB88
FB4F
FAD8
FAF0
FB53
FB52
FAF6
FAD3
FB0A
FB14
FAAC
FA53
FA91
FB26
FB65
FB2C
FAFB
FB23
FB5B
FB43
FB00
FAED
FB02
FAF3
FACD
FAF7
FB76
FBB6
FB5B
FAE6
FB0E
FBA9
FBDC
FB65
FB07
FB66
FBEB
FB94
FAB9
FB29
FE0D
023D
0548
05FF
0559
04E4
0506
0521
04E5
04BD
04FB
0542
051E
04C4
04C5
0527
0558
0500
0482
046C
04BD
0500
04FD
04E7
04EC
04EA
04C1
04A3
04C3
04F2
04D4
0476
0454
04A5
0504
04FB
04B3
04AC
04E7
04DF
046F
044B
04FD
05AA
0493
011B
FCE0
FA4C
FA2A
FB1C
FB75
FAFA
FA96
FACE
FB27
FB18
FAD6
FAE3
FB32
FB45
FB00
FADD
FB28
FB7E
FB63
FAFD
FAE1
FB34
FB80
FB5E
FB06
FAE3
FAFB
FB0A
FB09
FB31
FB77
FB7A
FB1F
FADC
FB14
FB72
FB67
FB1E
FB46
FBE8
FC08
FB13
FA40
FB9B
FF84
03D4
05FB
05A0
0492
0468
04F2
0529
04CF
0493
04D1
0515
04EC
049D
04AE
0506
051D
04CE
048C
04A8
04E2
04D9
04A0
048E
04B0
04C1
04B3
04CC
0520
054F
0510
04B1
04B5
0504
0508
0493
0438
0474
04E3
04CC
044B
044D
0509
052A
0320
FF2E
FB85
FA17
FAAC
FB83
FB76
FAF9
FB00
FB96
FBEF
FB9B
FB0A
FAD4
FAFA
FB15
FB08
FB13
FB56
FB93
FB8C
FB5A
FB40
FB47
FB4A
FB42
FB51
FB71
FB6E
FB39
FB18
FB46
FB8F
FB85
FB27
FAE9
FB13
FB5F
FB74
FB76
FBB4
FBF2
FB8F
FAB8
FAD7
FD3E
015C
04E5
0610
054D
0470
0487
0508
050D
049D
046D
04B7
04FD
04DE
04A1
04B0
04EE
04F3
04B8
04A0
04D7
0519
0515
04DD
04AC
0488
045B
043D
0461
04B1
04CF
04A2
0484
04B8
04F4
04D1
0474
0463
04AD
04BD
044C
0400
0495
0573
04DC
01DF
FDB5
FAB6
FA07
FABF
FB4F
FB2C
FAE8
FB04
FB4F
FB60
FB39
FB21
FB24
FB10
FAD4
FAA2
FA9D
FAB5
FACF
FAF7
FB35
FB69
FB6F
FB59
FB54
FB60
FB4A
FB0B
FAED
FB28
FB81
FB93
FB60
FB51
FB94
FBC3
FB77
FAFA
FB00
FBA0
FC05
FB89
FAEC
FBD7
FEFF
0305
05A5
05E7
04DA
0431
0480
051A
0544
050C
04E7
04F3
04F8
04E7
04FA
0545
057C
055C
0507
04D6
04DE
04ED
04E4
04E3
04FB
0509
04EE
04D0
04D9
04E6
04B4
0460
045F
04CD
0528
04F8
0481
0468
04B9
04D8
0485
0468
050B
0594
044B
00B9
FC99
FA3C
FA30
FB04
FB3E
FAD8
FAA9
FAF2
FB28
FAF1
FAAC
FAC6
FB15
FB28
FAFD
FAEB
FB01
FAF6
FABC
FAAD
FAFE
FB50
FB30
FACA
FAB8
FB1C
FB6A
FB3C
FAF0
FB14
FB87
FBA3
FB43
FB03
FB52
FBBF
FB95
FAF9
FAC3
FB3D
FB9D
FB3E
FAEA
FC40
FFAB
038A
05B9
05B1
04C7
0477
04EF
0561
054E
0508
0501
052C
0533
050A
04F6
0518
053D
052F
04FE
04D9
04C7
04AC
0491
04A1
04E4
051C
0515
04F3
04F8
051F
0520
04E1
04A0
0491
048E
046A
0468
04EB
058D
04F6
022F
FE0B
FAC0
F9D7
FABD
FBA8
FB90
FAF6
FAC6
FB13
FB47
FB22
FB07
FB3F
FB7F
FB64
FB0C
FAE4
FB01
FB13
FAF9
FAFA
FB4C
FBA3
FB8A
FB08
FA97
FA86
FAAC
FAD1
FB0A
FB6A
FBA5
FB6B
FB00
FB08
FB9B
FBF4
FB7E
FAEE
FBCB
FEAD
025D
04F6
05BF
058A
0566
057A
0550
04D0
047D
04B9
0542
0588
0561
0515
04E9
04D9
04CD
04CF
04E5
04EC
04BF
0481
0481
04D0
0520
0523
04EA
04C2
04C3
04C4
04B3
04BF
0501
052E
04F2
048C
04A8
055C
0589
03CA
0015
FC2D
FA1C
FA4F
FB67
FBD5
FB55
FAB3
FA8D
FABA
FAD0
FAC8
FADC
FB08
FB10
FAE9
FADD
FB16
FB5D
FB63
FB37
FB27
FB4D
FB6B
FB50
FB16
FAF7
FAF8
FAFF
FB16
FB54
FB8B
FB69
FB07
FAF9
FB8D
FC19
FBAB
FA7C
FA3B
FC6A
007E
0427
0592
0521
0493
04EF
059D
059D
04EB
0463
0487
04F5
0518
04F2
04E6
050C
0516
04E0
04B1
04CB
0507
0511
04E5
04C9
04D7
04DF
04CB
04D6
0527
056F
0544
04C9
0488
04A5
049D
0422
03D9
048E
05B9
056F
0271
FDEA
FA90
F9EA
FAF9
FBB6
FB66
FAE8
FB13
FB8D
FB8B
FB16
FAE7
FB42
FB96
FB61
FAF3
FAE9
FB44
FB72
FB2F
FAE7
FB05
FB52
FB4F
FAF9
FAC1
FADD
FB06
FAF9
FAE4
FB0A
FB3D
FB1E
FACD
FAD4
FB4D
FB86
FAFF
FA86
FBAF
FEFA
02EE
056B
05BF
0513
04D0
0526
054D
04E6
0475
0488
04EE
0517
04EC
04DC
051A
0544
04F5
046A
0437
0486
04DF
04D3
0488
046D
049E
04D8
04EE
04FD
0511
0503
04C5
04A1
04D1
0505
04C3
0449
0479
0586
0611
0450
0041
FC22
FA4A
FAD5
FBE2
FBE0
FB12
FAA6
FAF9
FB65
FB62
FB31
FB35
FB45
FB0F
FAC7
FAE0
FB45
FB5B
FAEA
FA87
FAC9
FB69
FBA9
FB62
FB2F
FB66
FB90
FB33
FAB6
FAE2
FBA4
FC05
FB7F
FACC
FAE0
FB77
FB78
FAC2
FADA
FD36
0137
048D
059C
04F7
0451
0478
04DB
04C6
0464
0450
04A3
04EA
04DE
04BB
04C7
04DE
04C2
0488
0481
04B1
04C5
0496
0473
04B7
053A
0576
053F
04F8
0500
052D
0517
04C5
04A7
04DD
04F6
04A4
045E
04C8
056C
04B8
01B1
FD76
FA77
FA03
FB16
FBBA
FB43
FAA3
FACE
FB77
FBAF
FB3A
FAC4
FAD2
FB24
FB4B
FB5B
FBA2
FC01
FBFD
FB82
FB13
FB1E
FB6D
FB89
FB64
FB4D
FB50
FB1E
FAB4
FA94
FB0B
FB97
FB82
FAF2
FAC7
FB51
FBB7
FB37
FA98
FBAB
FF13
032F
05A7
05CD
04FE
04C1
0533
0577
052B
04D1
04E7
0530
0526
04C8
0490
04B9
04F7
04F9
04D0
04BB
04BA
049B
045D
043D
0458
047F
0482
047F
04B0
04FB
0508
04C4
048A
04A0
04C2
0489
0425
0449
0516
0563
03B1
FFF8
FC18
FA32
FA97
FBAF
FBDC
FB0E
FA5E
FA7C
FAF6
FB11
FAC6
FA9C
FAD1
FB11
FB11
FB00
FB29
FB73
FB81
FB44
FB1D
FB4D
FB9E
FBB0
FB75
FB34
FB19
FB18
FB29
FB60
FBAA
FBB7
FB67
FB19
FB35
FB7C
FB4B
FAB7
FB04
FD67
0161
04D8
0612
0560
047C
0489
0527
0566
051B
04DE
0508
054F
0559
053E
0541
0548
0509
049B
0473
04C1
0523
051D
04BD
0470
0468
047A
0486
04AF
04FA
0516
04C4
045B
0465
04D0
04EC
0472
041B
04A9
057B
04C9
01A6
FD6D
FA95
FA3D
FB40
FBC9
FB56
FABE
FAB8
FAF8
FAE5
FA8D
FA76
FAC2
FB06
FAF5
FACC
FAE0
FB11
FB07
FAD4
FAE1
FB48
FB92
FB5F
FAF6
FAE7
FB41
FB83
FB6A
FB4D
FB8D
FBE7
FBD4
FB69
FB49
FBA3
FBBE
FB0E
FA7A
FBC2
FF6A
03A8
05FE
05B7
046E
040B
04C4
056B
0540
04C8
04D8
0562
05AA
055B
04E9
04D4
0503
050F
04E6
04CF
04EE
0518
052E
0547
056B
0562
050C
04B7
04CE
052B
0534
04B0
042C
043E
04A8
04B6
045C
045F
0504
0524
0334
FF50
FB8A
F9EE
FA73
FB60
FB6D
FAEC
FAD5
FB4A
FB94
FB44
FAC6
FAB5
FB0A
FB51
FB54
FB41
FB40
FB3A
FB1B
FAFE
FAFA
FAF8
FAE8
FAED
FB20
FB3D
FAF7
FA83
FA88
FB35
FBD1
FB95
FAC8
FA83
FB32
FBE3
FB85
FA9A
FB08
FDF2
0235
0565
0633
0570
04C1
04DA
0536
052E
04D8
04AD
04CF
04F2
04DD
04B7
04C0
04FA
0533
0542
0524
04E9
04A7
0484
049A
04D5
04F9
04EC
04D7
04ED
051A
0517
04DF
04CD
0518
0564
0527
0485
0452
04F0
0560
03FF
006F
FC6B
FA3E
FA7B
FB97
FBCE
FAFE
FA5F
FAB9
FB81
FBBA
FB40
FABC
FAA7
FAC9
FAC3
FAA6
FAB7
FAF4
FB1F
FB28
FB3A
FB57
FB45
FAF8
FAC6
FAF7
FB48
FB43
FAFA
FAF8
FB69
FBB4
FB55
FAC3
FAEA
FBCD
FC4E
FBC2
FB3F
FCA0
0037
0410
05E2
0566
044F
0428
04D5
0549
0517
04CC
04EC
0540
0547
0500
04D4
04F0
0515
050A
04EF
04F6
050E
0509
04F5
0506
0534
0534
04EA
04A4
04B4
04F0
04EA
0496
0462
0489
04A1
0438
03A6
03C5
0498
04B8
02A9
FEC4
FB42
FA15
FAF8
FBF4
FBAD
FAA6
FA34
FAB8
FB5C
FB60
FB03
FAF2
FB3F
FB60
FB12
FAB8
FAC0
FB05
FB1B
FAF5
FAED
FB2C
FB6C
FB62
FB28
FB04
FB06
FB10
FB29
FB6E
FBB6
FBB0
FB6F
FB7E
FC0B
FC5C
FBAA
FA8E
FAF1
FE00
027B
05B0
062C
0507
0451
04BD
0559
053A
04AC
0485
04E6
0533
050F
04CE
04D9
0512
0523
0511
0519
052D
0502
04A1
0478
04BF
050E
04E8
0479
045B
04AA
04D0
046F
0406
0446
04F3
051F
0488
0417
048B
0512
03E5
007F
FC93
FA69
FA89
FB7D
FBBB
FB31
FAC8
FAF0
FB39
FB30
FB01
FB06
FB26
FB04
FAA5
FA81
FAD8
FB4D
FB62
FB1F
FAF1
FB0D
FB35
FB2C
FB16
FB2F
FB5D
FB4E
FB06
FAF1
FB47
FBAA
FB98
FB30
FB0B
FB5B
FB95
FB50
FB3A
FCA2
FFD9
0374
0591
05B4
0512
0500
0587
05C7
054E
04A1
046A
04AB
04F1
0509
0525
055D
0573
0537
04E3
04D1
0502
0521
04F8
04AD
047A
0475
0499
04E4
0537
0546
04E9
046A
044A
04A2
04F7
04E8
04B6
04DA
050E
043F
01C4
FE5C
FBA9
FA9E
FABB
FAEB
FAC4
FAA8
FAE2
FB20
FAFC
FAA1
FA96
FAF3
FB3F
FB1B
FAC3
FAB3
FAFF
FB4E
FB65
FB66
FB74
FB68
FB1C
FAC9
FACA
FB10
FB29
FAEF
FAD0
FB2B
FBAF
FBC3
FB6B
FB49
FBA3
FBD1
FB37
FA84
FB61
FE86
0296
0553
05D2
0521
04CC
0535
05A1
057B
050D
04E5
0506
0505
04BF
0490
04BE
0504
04F3
0493
0463
04AC
051E
0532
04DF
049F
04C7
050E
04FD
049D
0467
0494
04CA
04B5
0497
04E8
0557
04B7
0231
FE76
FB56
FA17
FA6B
FB13
FB3D
FB09
FAE5
FAE9
FAEE
FAEA
FB00
FB2D
FB47
FB3C
FB3A
FB69
FBA4
FBA0
FB58
FB20
FB3B
FB87
FBA9
FB7F
FB41
FB34
FB4D
FB48
FB1B
FB12
FB64
FBB9
FB7C
FAC9
FAC8
FCB3
006A
0430
0625
05F3
04E3
045A
0493
04EC
04FB
04FC
0532
056D
055A
0515
04FF
051E
0507
0486
0416
0454
051D
05A0
0554
04A1
044D
047E
04AC
0483
0461
04BC
0544
0532
046C
03E3
045D
051D
0450
0122
FCF8
FA38
F9EE
FAF2
FB77
FAFA
FA5E
FA77
FB0E
FB68
FB50
FB23
FB23
FB1D
FAE7
FAB9
FADF
FB35
FB4C
FB08
FAC9
FAE1
FB23
FB31
FB11
FB2A
FB94
FBDD
FB9D
FB1E
FB0F
FB89
FBC1
FB13
FA33
FADE
FDFB
0253
057C
062B
0547
04A5
0503
059B
0587
04EE
049D
04D5
0517
0505
04EA
051E
0560
0539
04C3
049F
0502
0559
0511
0476
0451
04D1
0545
0517
04A5
04AE
0529
0540
0485
03BB
03F5
050A
0557
035A
FF71
FBB7
FA09
FA5D
FB28
FB30
FAAC
FA8A
FB0E
FB84
FB48
FAA2
FA54
FA96
FAEE
FB03
FB11
FB5B
FB95
FB52
FAC6
FAA2
FB22
FBA4
FB83
FAFA
FAC4
FB0A
FB32
FAE3
FAAA
FB23
FBE0
FBCF
FAD2
FA5B
FC06
FFBB
038E
0591
058C
04CB
0489
04DD
0522
04FF
04C3
04DA
053A
057D
0562
0516
04E3
04DC
04E2
04F5
0528
055F
0550
04EA
0485
047C
04AA
04A7
046C
047C
0519
05AC
055E
0458
03D6
04AA
05DB
055C
0242
FDF3
FAE1
FA32
FAEC
FB62
FB04
FA97
FADC
FB89
FBC7
FB54
FAC0
FA9C
FACD
FAE0
FAC0
FAC5
FB14
FB5A
FB46
FB07
FB04
FB35
FB2F
FADF
FABF
FB1E
FB8D
FB6A
FADE
FAC6
FB75
FC16
FBAF
FAA6
FAB2
FD0A
00ED
0441
0595
0541
04A2
049E
0501
0522
04CB
046D
0480
04EC
0531
0509
04B5
049E
04D8
0519
0525
050B
04F2
04DD
04C1
04C3
0500
053C
0519
04AB
0482
04E2
0540
0500
0471
048B
0570
05BF
03DC
FFF0
FC0B
FA2D
FA6B
FB50
FBA0
FB5D
FB24
FB2C
FB30
FAFF
FAD5
FAF9
FB51
FB7F
FB53
FB05
FAE8
FB08
FB2A
FB20
FAFB
FAEC
FAFE
FB10
FB16
FB32
FB6C
FB7D
FB27
FAB5
FAC6
FB65
FBC0
FB2B
FA64
FB33
FE79
02D5
05C3
0615
04F7
0464
04F0
0590
0540
0453
03E1
0452
0503
0534
04F3
04D4
0517
0564
055F
0524
04FC
04EC
04CA
04AB
04D5
053F
056B
050E
0492
049C
0519
0548
04D0
0470
0501
05EE
0561
0251
FDFB
FAD6
FA1C
FAD1
FB3E
FAD7
FA5C
FA82
FB11
FB69
FB63
FB50
FB55
FB39
FAE3
FAA2
FACC
FB3D
FB7C
FB4E
FAFF
FAFC
FB43
FB67
FB2D
FAE4
FAF3
FB3D
FB3B
FACB
FA7F
FAE3
FB90
FB84
FA9E
FA53
FC56
007E
048F
065D
05E8
04F2
04E0
0576
05B2
0548
04D6
04E0
052B
0533
04E5
0497
0483
049F
04D9
052D
057B
057C
051C
04A4
0477
049D
04C3
04B1
0497
04CB
0539
055C
04E7
0459
0484
0571
05D8
042B
004E
FC1A
F9CF
F9F9
FB1E
FB81
FAE2
FA46
FA69
FAEC
FB18
FADE
FAC0
FAF4
FB1E
FAF3
FAB7
FAD7
FB3E
FB75
FB50
FB2A
FB4E
FB7D
FB4D
FAD1
FAA0
FB0B
FBA4
FBBE
FB55
FB11
FB4D
FB7F
FB04
FA65
FB35
FE5C
02AB
05BC
0644
0541
04A5
0529
05E0
05CA
0520
04D1
052F
05A3
059F
0543
04F7
04CF
049C
046C
0483
04D1
04E8
0494
0445
0485
0528
0573
050E
047D
046B
04C8
04DF
0465
0403
0489
0594
057F
0302
FECD
FB25
F9CA
FA61
FB2A
FB0A
FA7B
FA78
FAFF
FB31
FAA8
FA11
FA26
FAB7
FB06
FAE9
FAE6
FB4A
FBAB
FB92
FB3A
FB3D
FB9D
FBBC
FB4D
FADD
FB0B
FB98
FBBF
FB51
FAFF
FB55
FBD9
FBA2
FABC
FA8C
FC84
006D
044D
0629
05CF
04C2
047B
0508
056F
0526
04BD
04FA
05BB
0627
05D3
053C
04F5
04E5
04A8
0455
045D
04C6
0506
04CD
0486
04BB
0532
0538
04B3
045D
04B1
051E
04D2
0409
03E0
04BD
0562
0414
0095
FC9B
FA3C
FA06
FACF
FB31
FAE9
FAA9
FAEE
FB5B
FB4A
FAB4
FA3E
FA69
FAF3
FB3E
FB27
FB11
FB35
FB51
FB2C
FB08
FB31
FB6B
FB35
FAA1
FA67
FAF2
FBAA
FBB9
FB3D
FB31
FBF3
FC86
FBDC
FA97
FAC4
FDA8
0227
05AF
06A4
05AA
049E
049A
0535
0580
054C
0527
0569
05B0
0574
04D7
0487
04D4
0541
052B
04A8
0458
0480
04BF
04C2
04C0
04FE
0535
04FA
047D
0465
04D5
0519
04A9
041E
0476
0573
055D
02DD
FEB5
FB25
F9BE
FA20
FAD9
FAFE
FABF
FAB3
FAFD
FB36
FB06
FA9E
FA7B
FACE
FB43
FB69
FB38
FB11
FB32
FB60
FB4A
FB15
FB28
FB7A
FB93
FB52
FB2E
FB70
FBA0
FB36
FAA3
FAE4
FBF3
FC75
FB7F
FA54
FB64
FF5F
040D
068D
0647
050E
04AB
0525
0571
051E
04BB
04D5
0538
0550
04F4
048B
0479
04B8
04FA
0509
04EB
04C7
04AF
0494
0469
0450
046E
04A8
04B6
0493
048B
04B9
04CB
0485
0453
04C4
056E
04CC
01D4
FD88
FA50
F9A0
FA98
FB56
FB16
FAA0
FAC5
FB41
FB52
FAE6
FAA3
FAEC
FB56
FB4E
FAF3
FAE8
FB64
FBEB
FBF8
FBA8
FB79
FB8B
FB88
FB3E
FB05
FB3E
FBA7
FB99
FB09
FACD
FB7E
FC60
FC2A
FAEF
FA9B
FCEB
0130
04C5
05CA
04EE
043F
04C0
05AF
05F7
0599
0545
0541
0538
04F3
04A6
0488
0483
0469
044E
0462
04A9
04E6
04E7
04B5
0481
0470
0489
04B7
04D7
04D2
04B1
0481
043B
03F9
041D
04C8
051C
03A7
0018
FC1F
FA02
FA46
FB4A
FB57
FA90
FA4B
FAF5
FB8F
FB47
FAAF
FAC6
FB74
FBC9
FB6C
FB00
FB0D
FB3C
FB0B
FAB9
FAEF
FBA6
FC11
FBB6
FB20
FB0F
FB72
FBA9
FB7B
FB4C
FB67
FB85
FB4A
FAEB
FB2A
FCAF
FF6D
028F
04F5
05E2
0583
04C8
0493
04F4
054C
0531
04E9
04DB
04FA
04F8
04DC
04F6
0549
0568
050D
0483
0448
0464
047D
0478
0497
04ED
050B
049F
0417
042A
04D0
0530
04CB
0443
047E
051F
0487
01B0
FDAA
FAC4
FA3C
FB1D
FB99
FB09
FA47
FA46
FAED
FB74
FB79
FB41
FB1F
FB09
FAE2
FAD4
FB13
FB71
FB83
FB33
FAE4
FAF9
FB5F
FBBA
FBCF
FBA8
FB69
FB3E
FB44
FB5D
FB3D
FAE5
FB08
FC8D
FF87
02CD
04F7
05A3
0589
0563
053F
04F2
04B6
04D7
0523
0526
04DB
04B4
04E6
0516
04E3
0484
0471
04AE
04CE
04AC
0498
04C0
04D4
04A6
048D
04D6
051D
04E3
047C
04B8
056B
04FB
0224
FDD3
FA93
F9EA
FAEB
FBA8
FB61
FACF
FAB3
FAF9
FB33
FB44
FB48
FB37
FB03
FAD4
FADD
FAFE
FAF3
FAD3
FB01
FB7E
FBC6
FB8B
FB2F
FB1F
FB27
FAE6
FAA3
FB02
FBD3
FBF4
FAEC
FA27
FBB7
FFC3
03F8
05EC
058E
04B3
04B1
052B
0533
04B8
0468
049B
04F9
051F
051C
0524
0526
0503
04DD
04E2
04F0
04C9
0481
046A
049D
04D9
04F0
04F9
0503
04CD
0444
03FB
0493
058C
053F
0297
FE89
FB54
FA4C
FAC2
FB33
FAF9
FA96
FA9B
FAF3
FB38
FB49
FB3B
FB0E
FACA
FAAE
FAE5
FB32
FB33
FAFB
FAFC
FB5B
FBA3
FB72
FB1E
FB32
FB8C
FB85
FB09
FAD8
FB52
FBAA
FB12
FA5D
FB87
FF3A
0388
05C9
057A
047F
0497
056E
059F
04D9
042B
0469
0526
0577
052B
04D2
04DA
0523
055C
0566
053B
04D8
046E
0455
0499
04D6
04C7
04A5
04B7
04C6
047E
0434
0498
056B
0522
0282
FE63
FB23
FA29
FAA5
FAFC
FABF
FAA7
FB13
FB80
FB73
FB30
FB25
FB33
FB00
FAB8
FAD3
FB36
FB36
FABB
FA8A
FB21
FBCE
FBA8
FAF0
FAB6
FB44
FBBD
FB7E
FB18
FB47
FB9C
FB32
FA94
FBB5
FF61
03B0
05E7
058C
0493
04B5
0591
05C8
050C
044F
044A
04A5
04C8
04B9
04CB
04F3
04F6
04E7
04FA
0517
0507
04EF
0511
0539
04E6
042E
03E2
047B
0543
053F
049F
0483
0513
04C3
0235
FE39
FB22
FA36
FAA3
FAF3
FAC5
FAAC
FAED
FB2A
FB2F
FB46
FB8D
FB98
FB26
FAB6
FADF
FB55
FB51
FAC0
FA72
FAEE
FBA4
FBB9
FB3A
FAF6
FB44
FBA3
FBA1
FB81
FB8E
FB66
FAB0
FA4A
FBD5
FFAD
03F2
0636
05EF
04BD
045E
04E6
054D
0514
04B2
04A9
04D5
04D7
04B9
04C4
04F5
0504
04DA
04B3
04B8
04CA
04D1
04EB
0515
0504
048D
040D
03FA
043F
0466
0470
04DE
0596
0545
02A6
FE5E
FAD1
F9B7
FA79
FB46
FB45
FB00
FB05
FB1A
FAEC
FACC
FB25
FBA2
FB8B
FAF4
FAB7
FB2B
FB94
FB4E
FAC5
FABF
FB2E
FB6A
FB58
FB81
FC00
FC27
FB8D
FAE3
FAF8
FB63
FB2A
FAAC
FBBC
FF32
0355
059D
058E
04D8
04E8
0564
0553
04BD
047A
04C7
0508
04E7
04DA
0531
0572
051D
0492
0480
04D3
04EC
04A1
0462
046B
0471
044C
0462
04EB
054F
04E4
042F
0464
056F
056E
02CF
FE7C
FB0D
FA07
FAA1
FB38
FB31
FB05
FB19
FB3E
FB40
FB3F
FB4C
FB2A
FAC8
FA8D
FAD2
FB47
FB5C
FB16
FAF9
FB34
FB61
FB36
FB06
FB3D
FBA3
FBA0
FB2A
FAE5
FB1F
FB45
FAD1
FA83
FBE6
FF66
036A
05C2
05D1
04E0
0471
04B9
04F4
04B6
0461
0469
04B0
04D8
04DA
04F6
052B
052E
04EA
04AB
04B1
04DA
04EA
04E6
04EF
04EF
04C1
048C
049B
04DC
04E7
04B5
04D0
0557
0524
02CD
FEA8
FB05
F9DA
FABA
FBA5
FB75
FAC7
FA9B
FAEF
FB2C
FB34
FB5D
FB96
FB61
FAC9
FA93
FB1B
FBB7
FBAE
FB45
FB2E
FB62
FB4C
FAE0
FABD
FB1D
FB66
FB27
FAEC
FB58
FBE0
FB75
FA94
FB53
FEB9
0304
057C
0584
04D0
04DF
0569
0579
0512
04EC
0516
04EF
045B
0420
04AD
0559
0566
0508
04DD
04D6
0485
0423
045A
051C
057F
0503
045B
045C
04BC
049A
0417
044C
0554
0573
0311
FEFD
FBBC
FAC1
FB2F
FB67
FAF4
FA85
FA99
FAEB
FB1D
FB3C
FB64
FB5B
FAF4
FA82
FA7D
FADC
FB34
FB50
FB4E
FB3D
FB07
FACD
FAF0
FB7F
FBEF
FBB8
FB2C
FB18
FB96
FBBD
FAF5
FA3D
FB5D
FECA
02C4
0511
053B
04AD
04CC
057E
05C7
054D
04B6
049F
04E5
050C
0503
050C
052A
0518
04D0
04AB
04D7
050E
0515
0512
052E
0529
04C7
0459
046E
04E6
0505
049A
0475
0518
0557
0359
FF2D
FB49
F9EC
FAAA
FB61
FB05
FA7A
FAC5
FB78
FB8A
FAF4
FAA2
FAF7
FB4F
FB21
FACB
FACA
FAEC
FAD3
FAB2
FAE3
FB24
FAFD
FAA6
FABF
FB40
FB65
FAF0
FAB5
FB53
FBEF
FB5C
FA5E
FB57
FF2E
039F
05B0
0513
040C
044C
053A
0578
04F3
04A4
04E5
051B
04EF
04DF
0541
0593
0557
04F3
04FE
0539
0505
048E
049B
053E
0593
050F
0469
048F
0534
0545
04AB
0486
053E
0551
0312
FF0B
FBB6
FAB5
FB46
FBA2
FB32
FAC5
FB03
FB81
FB81
FB00
FA90
FA8C
FAD3
FB22
FB4B
FB25
FAB1
FA4E
FA71
FB06
FB6F
FB4C
FAF1
FAE4
FB12
FB00
FAB7
FAD8
FB88
FBE2
FB21
FA2B
FB08
FE85
02DD
056B
0565
045D
0418
04A2
04F2
04A0
0453
0489
04E1
04D4
0496
04B7
0536
0587
0575
055C
0572
055A
04DC
0470
04A0
0531
056A
0521
04D4
04CB
04B4
046C
0484
0539
055D
034D
FF47
FBBB
FAB0
FB89
FC1E
FB8C
FAE3
FB28
FBD5
FBD2
FB29
FAD8
FB39
FB91
FB4C
FAD6
FABC
FAC6
FA90
FA67
FACF
FB7C
FBA0
FB21
FAC6
FB03
FB54
FB2E
FAF9
FB58
FBD3
FB69
FA84
FB28
FE66
0290
04F8
04FE
0461
04A2
0553
0550
04A5
0456
04AB
04DA
0471
041F
0490
0542
054F
04CE
049D
0506
0564
0537
04CA
049A
049E
0497
04A8
0505
0548
04DB
0429
045F
0594
05EE
0396
FF34
FB83
FA5C
FAEC
FB42
FAC2
FA69
FAE9
FB95
FB82
FAE7
FAAD
FB16
FB83
FB79
FB35
FB1E
FB2B
FB22
FB1F
FB5E
FBB7
FBB7
FB50
FAFD
FB10
FB45
FB4D
FB4B
FB6C
FB56
FAAB
FA1C
FB37
FE9E
02D0
056C
05AD
04F2
04D7
0564
0599
0527
04C2
04ED
053A
0513
04A9
0499
04EE
0512
04C7
0481
04A4
04EC
04E9
04AF
0494
0494
0480
0477
04C1
0525
050E
048A
0479
052D
054C
0312
FECA
FB0C
F9FA
FAF4
FBB8
FB3D
FA80
FA9D
FB45
FB77
FB15
FADB
FB16
FB3E
FB01
FAD2
FB11
FB4F
FAFB
FA68
FA65
FB0B
FB98
FB8C
FB3D
FB2B
FB42
FB2C
FB10
FB56
FBD2
FBEA
FBC3
FC8A
FF0B
025E
04BC
055C
0509
04D4
04F9
051C
0523
0543
056B
0547
04DA
049E
04D0
050E
04F6
04C9
04FF
057D
05AA
054E
04DB
04BE
04DA
04DD
04C9
04CD
04C5
0469
0402
043B
04F1
04B9
024F
FE4F
FAF1
F9D5
FA85
FB58
FB60
FAFF
FAD8
FAE3
FACC
FAAA
FADB
FB4F
FB87
FB4B
FAF6
FAEA
FB07
FAF5
FAB7
FAAA
FAE5
FB0D
FAEA
FAD8
FB53
FC2C
FC8B
FBF1
FAF9
FAF9
FCD5
0030
03AB
05E0
0651
059D
04E1
04D6
054C
0599
0564
0504
04F9
0548
057A
053C
04C0
047B
049F
04F0
0517
04FC
04D1
04D3
050E
0541
0512
047B
0407
044F
0512
050E
0315
FF70
FBE2
FA17
FA32
FAF6
FB45
FB11
FAE9
FAFF
FB0D
FAE9
FAC6
FACE
FAD3
FAA5
FA7B
FAB1
FB35
FB7B
FB32
FABB
FAA4
FAE9
FB06
FACD
FABC
FB40
FBE2
FBBC
FACC
FA71
FC2D
FFF0
03E5
0617
0621
0532
049E
04B9
0501
0503
04D4
04C2
04E9
0523
0546
053D
050C
04CE
04B6
04DC
0517
0518
04DD
04C4
0517
0584
0568
04A4
03FB
044D
055F
05BC
0407
006D
FCA2
FA68
FA20
FAC8
FB30
FB01
FAB2
FAB5
FAF8
FB24
FB13
FAF2
FAED
FB03
FB1B
FB30
FB3B
FB25
FAE9
FABF
FAE7
FB3F
FB52
FAF1
FAA7
FB0D
FBD4
FBE7
FAE3
FA1D
FB84
FF64
03B2
05F2
05AD
0499
0469
051D
059B
055F
04F4
04E8
050A
04E1
0482
046B
04B6
04F8
04ED
04DD
0515
0558
0538
04CE
04A8
04EA
0506
048A
03F1
041C
0507
0560
03C9
005F
FCC2
FA9F
FA50
FAE4
FB41
FB0D
FAA9
FA92
FAD7
FB2D
FB53
FB47
FB2B
FB17
FB0F
FB13
FB1E
FB1A
FAF0
FAB7
FAAE
FAE8
FB1E
FB0D
FAF6
FB50
FBFC
FC1A
FB3B
FA74
FBA2
FF48
0387
05D0
0584
0466
0461
056B
0612
0590
04A6
045D
04B6
04F6
04DB
04D5
0526
0568
0533
04CE
04C5
0509
050E
04AD
046E
04AC
04EE
0491
03E2
03F1
050C
05DF
049D
010A
FCEE
FA71
FA23
FADC
FB36
FADD
FA6F
FA77
FAD9
FB29
FB3F
FB40
FB3F
FB1B
FAC2
FA6D
FA6D
FAC5
FB28
FB54
FB5A
FB64
FB65
FB43
FB31
FB86
FC11
FC09
FB0F
FA2B
FB2A
FEAA
030A
05C9
05F8
04EF
047F
0501
0578
0538
04BB
04B4
0505
050F
04C2
04B7
0537
05B4
0589
04E8
048F
04B7
04E3
04B8
0492
04D8
0531
04DE
03F0
0385
0454
055A
0494
0139
FCE0
FA13
F9E1
FB1B
FBE0
FB8D
FAEC
FAD8
FB32
FB4D
FAFD
FABF
FAEF
FB42
FB34
FAC3
FA6E
FA8B
FAE2
FB17
FB23
FB34
FB3A
FB0D
FADF
FB2C
FBE5
FC39
FB93
FAD2
FBC2
FF17
0340
05C5
05C2
0499
041E
04A1
0522
04F9
04A1
04C1
052B
0536
04CA
0483
04C6
0532
0540
0510
0526
0584
058E
04EE
042D
040F
048A
04D9
0497
045B
04D1
056D
0499
0177
FD3A
FA3C
F9C8
FAEE
FBBD
FB54
FA80
FA64
FB0A
FB8B
FB5E
FAF0
FADF
FB1F
FB2F
FAEC
FABA
FAD7
FB00
FAEE
FADE
FB35
FBC2
FBEA
FB94
FB68
FBC7
FBFB
FB2C
F9F7
FA60
FD99
024C
05AD
064A
0544
04A4
0511
059D
0572
04E3
04AE
04E0
04E9
0496
045E
04A4
0520
0547
0514
04F5
0514
0518
04BD
0454
0455
04AA
04B6
043D
03E4
0466
055C
0534
02BF
FEB2
FB33
F9E3
FA6D
FB31
FB1D
FA8F
FA6D
FADC
FB38
FB1F
FAEB
FB0E
FB5B
FB5A
FB0F
FAF6
FB33
FB44
FACE
FA50
FA8A
FB5D
FBD6
FB78
FAF6
FB2D
FBCD
FBC3
FAFD
FB0C
FD68
016C
04B9
05AA
04EC
045B
04CA
0577
0575
04E5
0491
04C7
0517
0521
0511
0531
055C
0530
04BB
047A
04B8
0528
0551
052B
050E
0510
04E0
045C
0404
0471
054A
0523
02DF
FF0F
FBB1
FA56
FABE
FB66
FB4E
FACE
FAB8
FB22
FB60
FB11
FAA0
FA96
FAD8
FAED
FAC7
FAD4
FB43
FB9D
FB6B
FAF0
FACE
FB19
FB39
FAE4
FAAC
FB30
FBF7
FBE2
FADA
FA7A
FC7E
0095
0466
05E7
054A
0461
046B
0502
0530
04DC
04BC
0530
05B6
05AD
0526
04B6
04A2
04AC
049E
04A6
04EC
052A
04F8
0479
044A
04A7
050C
04EC
0490
04C1
0573
0550
0310
FF24
FBA5
FA4E
FAE3
FBBC
FBB3
FB10
FAB5
FADF
FB0F
FAEE
FABF
FADB
FB24
FB43
FB35
FB44
FB7E
FB83
FB1D
FAAB
FABC
FB46
FBA4
FB6B
FAFE
FAF9
FB44
FB28
FA83
FA78
FC6F
0052
0433
0603
058B
0472
044D
0516
05AC
056E
04E3
04C3
04F5
04E0
046D
0430
0487
0500
04F7
047D
043E
0490
0510
0548
0553
0570
056C
04E7
043A
0457
0565
05EF
042E
0031
FC29
FA46
FA91
FB4B
FB26
FA78
FA44
FAB9
FB22
FB11
FAE6
FB18
FB76
FB7C
FB25
FAF5
FB31
FB7F
FB74
FB2C
FB17
FB4C
FB67
FB32
FB00
FB2F
FB76
FB2A
FA4D
FA0F
FBCC
FF85
0388
05E1
0607
051D
0497
04DB
0549
0549
04FA
04D1
04EA
0501
04F0
04E6
0509
052E
051E
04F5
04F5
050A
04D3
0445
03EA
0436
04CF
04F6
04A0
049E
055C
05C5
0425
0043
FC15
F9FA
FA60
FB9D
FBF7
FB56
FAC5
FAD3
FB0C
FAED
FAB1
FAD6
FB3F
FB4D
FACE
FA54
FA6A
FAE1
FB29
FB2C
FB55
FBC2
FBEF
FB7F
FAF6
FB25
FBE4
FC0B
FB04
FA0E
FB36
FEF5
0351
05C5
05B8
04BB
0478
04F9
0535
04C0
0447
0472
04F7
051C
04D3
04B9
051A
0580
0564
04FA
04DB
051A
0529
04BD
0457
048F
0520
0535
04A3
0447
04CE
0564
0450
00F8
FCE8
FA6D
FA4C
FB37
FB85
FAF8
FA8F
FAF6
FBAB
FBD3
FB61
FB04
FB21
FB53
FB23
FABF
FAB7
FB1B
FB5D
FB1D
FAB8
FABD
FB1D
FB4B
FB11
FAD9
FAF2
FAFD
FA9B
FA76
FBEF
FF6B
035C
058E
0568
0466
0442
0510
0594
0517
0452
044C
04F6
0559
04F9
0468
046E
04F6
054B
0516
04BD
04BB
04FD
0521
0519
0524
054D
0547
04FC
04E0
0541
0576
0435
0100
FD0F
FA62
F9EC
FAD6
FB99
FB8B
FB21
FAF8
FB15
FB21
FB12
FB22
FB5B
FB75
FB4A
FB13
FB10
FB25
FB0E
FADA
FAE4
FB31
FB47
FADB
FA63
FA92
FB40
FB72
FAB3
FA21
FB7D
FF1C
0334
058A
059F
04D9
04AE
0527
055C
04EB
0470
0487
04F4
0505
049A
044C
048E
0512
053B
04F7
04CA
0506
055E
0562
051C
04F5
0508
04FD
04B3
049F
051C
057A
0456
0129
FD3E
FAAA
FA45
FB03
FB59
FAEB
FA89
FACD
FB50
FB65
FB18
FB05
FB5F
FBAB
FB79
FB08
FAE6
FB1E
FB36
FAEF
FAA3
FAB6
FAFB
FAF7
FAA8
FA97
FB0A
FB82
FB61
FAFB
FB9B
FE2D
0202
0532
0650
05A9
04B7
048B
04FB
0544
0519
04D9
04D7
04E0
04A7
0454
0458
04B8
04F7
04CF
049C
04D1
0536
0533
04BC
0484
0502
05A9
05A3
0508
04B6
04D2
041F
017F
FDAF
FAD5
FA41
FB20
FBB1
FB49
FAA8
FA95
FAE2
FAFE
FAE9
FB06
FB5D
FB8D
FB65
FB2B
FB2C
FB5C
FB7C
FB73
FB51
FB24
FB0B
FB3A
FB9A
FB92
FABB
F9EA
FAD2
FE2B
027B
0556
05BF
04E5
0475
04D0
052D
0506
04B6
04B7
04F2
0514
051D
052E
052A
04EA
049E
0490
04A7
0492
0463
0480
04DF
04DB
0435
03D4
049F
05BD
04FD
017A
FD1E
FAB5
FAE1
FBC9
FBA8
FABE
FA56
FAC5
FB3D
FB3E
FB38
FB87
FBB4
FB4D
FAC6
FADE
FB70
FBAC
FB50
FAF6
FB0F
FB44
FB2F
FB1F
FB7F
FBD8
FB62
FAA3
FB6D
FEA4
02BC
053D
057B
04EA
04EF
054E
051F
0470
0429
049A
050C
04EA
0493
049A
04D4
04C9
048C
048D
04CD
04DF
04B9
04C2
0505
04EF
044F
0401
04C3
059B
0477
00CC
FCAF
FA9D
FAC5
FB50
FAFF
FA6C
FA9E
FB5E
FBB1
FB62
FB31
FB80
FBBA
FB57
FAC0
FAA2
FAF0
FB26
FB30
FB61
FBA1
FB79
FAF9
FADE
FB72
FBDB
FB4F
FAAD
FBE1
FF6D
0361
056B
0550
04AA
04A8
04F7
04DE
047D
046F
04C4
0504
050E
0534
057B
0564
04C9
044C
046E
04CD
04C0
046B
0476
04DA
04D6
0440
040D
04E1
058D
0414
0044
FC56
FA89
FAC2
FB3E
FB0B
FAC8
FB2C
FBC6
FBBB
FB13
FA99
FAAD
FAE6
FAE7
FADF
FB04
FB1A
FAF5
FAEE
FB53
FBBC
FB9A
FB2F
FB47
FBDD
FBE2
FADF
FA3B
FBF2
0000
03FF
05B4
0550
04A8
04C8
0531
0525
04CC
04AD
04C7
04C1
04A6
04D1
052F
053F
04E7
04AA
04D1
04E6
0484
0429
047D
052A
0531
0474
0419
04C8
0541
039B
FFCE
FC1C
FA8D
FAD4
FB3E
FB01
FABA
FAF6
FB43
FB11
FAAE
FAC4
FB43
FB7D
FB37
FAF7
FB18
FB40
FB24
FB22
FB94
FC03
FBB7
FAF2
FAB5
FB41
FB9D
FB21
FAEB
FCBE
008E
0423
0584
0512
0491
04D0
0524
04EB
048C
04A9
0511
0520
04D2
04B9
04FD
051C
04CE
0483
0497
04B0
0463
0412
045D
0503
051E
0496
0472
052D
056C
0350
FF1B
FB62
FA41
FB1C
FBCE
FB64
FAC3
FAE1
FB69
FB83
FB22
FAE3
FB01
FB18
FAF9
FAFC
FB4A
FB7D
FB51
FB2C
FB6E
FBB8
FB7C
FB07
FB28
FBCC
FBDA
FAF0
FA94
FCAD
00E5
0497
05B3
04DD
042F
0489
050E
04EE
0487
048F
04E4
04EC
04A7
04A3
04FE
0528
04D8
0485
0498
04BA
047F
043A
047B
04FE
04F4
045F
0445
0501
0524
02F1
FED4
FB59
FA5F
FB20
FB99
FB1F
FAAF
FB0C
FBA3
FB9A
FB19
FAED
FB43
FB87
FB5D
FB1E
FB23
FB3E
FB3B
FB4C
FB93
FBAE
FB4A
FAE0
FB21
FBC3
FBB6
FADD
FAD6
FD3B
0162
04BC
05A5
04FA
0491
04EB
0525
04BC
044A
046C
04D7
04E8
04A8
0499
04CB
04D1
0499
049A
04F6
051D
04B2
0442
0476
04F7
04EA
0460
045B
0510
0504
02A4
FE90
FB45
FA63
FB0E
FB71
FB0A
FAB7
FB01
FB61
FB4C
FB11
FB38
FB9A
FBA3
FB45
FB0F
FB3B
FB5B
FB22
FAEA
FB12
FB55
FB4C
FB2D
FB68
FBB8
FB68
FABA
FB43
FE1A
0227
04F8
0565
04A1
0463
04E2
0528
04D2
0483
04AF
04EA
04B6
045D
047C
0501
0540
04FD
04B5
04C4
04D8
04A9
0486
04C5
0504
04B8
043C
0468
0502
0466
0172
FD54
FA98
FA5E
FB50
FB9C
FB17
FAD9
FB51
FBC6
FB9E
FB39
FB2B
FB51
FB27
FAC2
FABC
FB33
FB8E
FB65
FB16
FB1A
FB4C
FB51
FB52
FB9C
FBD9
FB71
FAD8
FBA4
FEBC
02D4
057E
05C0
04E5
0492
04E6
04F5
0480
0435
0482
04F3
0503
04DF
04F4
0522
04F7
048D
047E
04F0
0544
050A
04A2
0482
0476
0429
0403
04A2
0568
048A
012A
FCDC
FA3C
FA23
FB0B
FB43
FAD8
FAD3
FB56
FB8E
FB21
FABF
FB01
FB7E
FB76
FAFD
FACB
FB18
FB58
FB27
FAE4
FAF8
FB32
FB3C
FB41
FB87
FBB3
FB44
FACE
FBD9
FF0F
0303
0579
05BE
051E
04FE
0552
054E
04DB
0498
04C4
04F7
04E6
04D5
0507
0536
0512
04CF
04DC
0519
0509
04AF
049E
04F1
04F5
0457
03F6
049F
0563
0434
007C
FC4C
FA3E
FAA1
FB7F
FB4A
FA82
FA63
FAFF
FB64
FB30
FAED
FB05
FB25
FAF3
FAB0
FAC5
FB09
FB0B
FAE1
FB06
FB73
FB93
FB42
FB28
FB95
FBC6
FB14
FA81
FBFA
FFDA
03FE
05EE
057B
048A
048E
0523
0547
04F9
04DF
0515
051A
04D9
04D2
0534
057A
0532
04BC
04B1
04F4
04F1
049D
048A
04DB
04F3
0492
0475
051C
056A
039E
FFB2
FBE2
FA59
FADE
FB85
FB3E
FABE
FAEA
FB61
FB45
FAAD
FA70
FAC9
FB13
FAEA
FAC2
FB1A
FBA1
FBAF
FB47
FAFF
FB0A
FB08
FAE2
FB10
FBA3
FBC9
FB0D
FAA2
FC5C
0052
0444
05ED
055F
0485
04A5
0539
0544
04D9
04B4
04FA
0520
04EE
04CC
04FD
052B
04F4
048E
0474
04B2
04EC
04FE
050C
0505
04A9
043C
0486
0587
05B5
036B
FF19
FB43
F9FA
FAC8
FB9B
FB4B
FA94
FA92
FB33
FB95
FB64
FB18
FB14
FB35
FB38
FB2B
FB2D
FB2A
FB0D
FAFC
FB1E
FB43
FB2B
FB0D
FB4D
FBAE
FB6E
FA94
FA92
FCDB
00F3
0493
05EC
055D
049C
04A6
0514
0533
0508
04F3
04F1
04C4
048A
0497
04E8
0518
04FA
04D1
04D4
04E0
04D0
04D0
0501
0508
048D
0412
0482
059B
058D
02E1
FE7E
FB01
FA0B
FAC4
FB4E
FB03
FAAC
FAEC
FB57
FB4F
FB01
FAF5
FB29
FB2A
FAF0
FAE8
FB3A
FB80
FB68
FB31
FB31
FB43
FB17
FADB
FAFF
FB4F
FB17
FA78
FAE7
FD9A
01B9
04EE
05D5
053C
04CC
050C
0545
04F7
0498
04B3
050B
0517
04E0
04D4
0505
0518
04E7
04B3
04A7
04A2
0493
04B3
050C
0526
04B1
044C
04D1
05C2
053C
021F
FDC6
FACC
FA4F
FB11
FB5C
FAF3
FABA
FB11
FB68
FB51
FB2A
FB52
FB7C
FB3B
FAD1
FAC9
FB17
FB35
FB0A
FB09
FB5A
FB7B
FB21
FADC
FB4B
FBE3
FB8B
FA8F
FAED
FDFD
0264
0557
05A1
04AC
045F
04F2
054D
04F1
0482
049B
04E6
04DB
04A3
04B5
0502
051C
04FA
04F5
051B
0510
04B8
047E
049E
04AE
044F
040A
04A0
057D
04D1
01AF
FD90
FAE5
FA84
FB25
FB52
FAFD
FAEC
FB42
FB68
FB21
FAEE
FB2E
FB7E
FB66
FB15
FB01
FB22
FB1B
FAF2
FB02
FB45
FB43
FAE5
FAC8
FB53
FBDB
FB80
FACB
FB88
FE9A
0291
051A
0575
04E0
04B6
04FE
050C
04CC
04BE
04FC
0509
04B0
0474
04C1
0535
0527
04A3
044E
0477
04C8
04EE
0505
052A
051C
04B8
0481
04FB
057B
0465
010B
FCEE
FA70
FA5E
FB52
FB94
FAF2
FA75
FAB9
FB3D
FB4E
FB08
FB09
FB6F
FBB7
FB85
FB26
FB15
FB4D
FB5C
FB16
FADD
FB20
FB9E
FB99
FAD4
FA44
FB62
FE9B
029D
0559
05E3
0523
04A4
04EE
054F
051C
049F
048C
04EF
0521
04C7
0455
045E
04C0
04DF
0496
0471
04CD
0530
04F4
0453
0442
050D
058B
042B
00C2
FCF5
FAB3
FA70
FB0F
FB51
FB09
FAD3
FB0A
FB5B
FB5F
FB2B
FB1D
FB45
FB4B
FB07
FAD4
FB1B
FBA4
FBC3
FB45
FACA
FAFA
FB90
FB99
FAD7
FA7D
FC17
FFBA
039C
05B6
059E
04A7
0446
04B8
0536
0527
04BD
0483
049B
04B6
049C
0474
047D
04AC
04C6
04C8
04E4
0520
0529
04C1
0448
0473
0542
0586
03DA
0042
FC7B
FA69
FA58
FAFB
FB19
FAC6
FAD3
FB70
FBE4
FBA0
FB07
FADE
FB3C
FB82
FB4E
FB06
FB2E
FB9B
FBA8
FB2F
FAD8
FB2A
FBB9
FB9A
FAC2
FA77
FC1E
FFA9
036D
059C
05D0
051A
04B0
04D7
0509
04E2
0495
047C
0491
0496
048A
04B0
0515
0553
0512
0498
0483
04E9
0521
04A8
03FC
041C
0516
0583
03D6
0020
FC3F
FA30
FA41
FB25
FB7E
FB20
FACB
FB03
FB7D
FBA4
FB5C
FB18
FB2C
FB5D
FB41
FAE5
FAC8
FB26
FB96
FB88
FB15
FAE3
FB37
FB7E
FB34
FAFD
FC4B
FF93
035F
0593
0592
04B3
0488
0531
05A5
0546
0495
0454
048B
04BF
04C2
04D2
0502
0504
04AF
045F
047F
04E1
04ED
0480
0438
04B3
058A
0576
0382
000C
FC98
FA9E
FA6C
FB19
FB74
FB1D
FAA3
FAAF
FB2F
FB7D
FB3D
FAD1
FAC7
FB16
FB45
FB2E
FB33
FB8D
FBD7
FB9F
FB2B
FB2C
FB9F
FBB0
FAFB
FA96
FC29
FFDF
03CC
05C4
0584
049A
0472
04F3
052C
04CF
0478
04B0
052E
0552
0508
04C7
04DB
04FA
04C8
046A
0453
049E
04D6
04A1
0453
0497
0558
055F
0366
FFA1
FBEB
FA22
FA6F
FB5D
FB87
FAF4
FA93
FAD5
FB33
FB24
FAE1
FAF7
FB60
FB8A
FB3E
FAF8
FB31
FB9D
FB92
FB0B
FAC7
FB36
FBB7
FB66
FA80
FA82
FCA5
0069
03E5
058C
056F
04D5
04C1
0520
0547
04F3
0491
049F
04FF
0526
04D8
0481
049C
0505
051F
04B7
0454
047A
04E6
04EC
0487
047E
0521
0555
038A
FFBE
FBF4
FA40
FAAC
FB77
FB4C
FA96
FA80
FB3C
FBDA
FBB2
FB39
FB2F
FB84
FB8A
FB12
FAC0
FB15
FBA9
FBB4
FB30
FAE8
FB58
FBE4
FBA2
FAC1
FAB8
FCCE
0097
0427
05CB
0576
0486
043C
04AB
0510
04E6
0470
043A
0463
0498
049B
0492
04B0
04DD
04D6
04A8
04A5
04E3
04F7
0495
0429
046F
053D
0529
02DB
FEC9
FB2C
F9EA
FAC6
FBD7
FBC3
FAFB
FAC2
FB66
FBFA
FBBA
FB11
FAF3
FB80
FBEA
FB9D
FB08
FAF1
FB56
FB84
FB30
FAF4
FB5E
FBF5
FBC6
FAED
FAF3
FD38
0129
0498
05E1
0568
04CB
04E7
0537
04F6
0455
0429
04AD
052E
04FE
045F
041D
0477
04DC
04CA
0483
049B
0503
050E
0474
03EA
044A
0535
0515
02B9
FED4
FB7B
FA30
FA9A
FB40
FB3D
FAE0
FAD4
FB22
FB47
FB0F
FADF
FB17
FB80
FB9A
FB53
FB1E
FB4F
FBA2
FBA5
FB65
FB61
FBC0
FBEA
FB50
FA76
FAD7
FD6B
015B
0490
0596
04EB
043B
048A
055C
05A8
053C
04CC
04E1
0529
0513
04B2
0498
04E9
050F
0497
03F5
03F5
0492
04E4
046A
03E4
0455
055D
053A
02B2
FEB2
FB7B
FA66
FAD2
FB4B
FB37
FB04
FB14
FB28
FAEB
FA99
FAB3
FB35
FB8C
FB5D
FAFE
FB01
FB68
FBB3
FB93
FB5D
FB8A
FBF9
FBFB
FB36
FA60
FADD
FD70
014A
048B
05DC
057E
04CA
04B6
0509
050E
04B0
048D
04FB
0570
0540
0494
0440
049E
0512
04E9
045A
0432
049D
04E1
047F
041A
0495
0588
0533
026C
FE34
FAEE
FA07
FAC5
FB6F
FB39
FABB
FABE
FB32
FB76
FB44
FAF3
FAE2
FB06
FB1E
FB28
FB53
FB95
FB9C
FB40
FAE3
FB0B
FBA5
FBF2
FB65
FA9E
FB24
FDDF
01E8
0519
0602
0528
0443
0465
051D
0565
04FD
0490
04A4
04FA
050A
04D2
04BF
04EF
0502
04C1
048C
04D1
0541
051C
0453
03DE
0482
0575
04D8
01CD
FDAC
FAD8
FA62
FB39
FBA8
FB33
FAB0
FAD8
FB57
FB6D
FB07
FAC8
FB18
FB8D
FB88
FB10
FABD
FAE3
FB23
FB07
FABA
FAD2
FB69
FBCC
FB62
FAC1
FB61
FE1E
020D
0523
060D
0548
0462
0457
04DD
0526
04F6
04B9
04C8
04EC
04CC
047C
0465
04AB
04F9
04FC
04DA
04EA
0521
0515
04B4
0486
04FA
0572
0493
01AB
FDBF
FACF
FA07
FAC9
FB8E
FB7D
FAF7
FAC5
FB13
FB66
FB5F
FB25
FB11
FB34
FB54
FB54
FB57
FB6F
FB6D
FB2A
FADE
FAEF
FB50
FB68
FAD7
FA54
FB4A
FE5B
025F
053F
05E7
0525
0496
04E1
055C
053D
04AC
0469
04B4
0509
04F1
04A9
04AE
04F4
04F6
048A
043A
0483
0517
0535
04C4
0491
0525
05B9
04BC
0196
FD98
FAD8
FA41
FAF0
FB69
FB25
FABC
FAD2
FB42
FB7A
FB4A
FB0F
FB16
FB38
FB30
FB0F
FB23
FB68
FB7B
FB2C
FADE
FB0B
FB7F
FB75
FAB2
FA3A
FB84
FED6
02B9
0537
059C
04E5
0479
04CA
053E
0534
04C8
048B
04BF
0515
0524
04E5
049F
0486
0491
04AF
04EC
0541
0566
0515
048F
047D
051C
058F
046B
0135
FD39
FA8D
FA29
FB21
FBCA
FB78
FAD6
FABB
FB17
FB45
FB07
FAD1
FB05
FB5E
FB62
FB1E
FB13
FB5D
FB77
FB01
FA70
FA90
FB4F
FBAA
FB0C
FA6F
FB88
FECD
02AA
0507
0554
04CB
04C2
0542
0574
04FF
0479
048A
050C
0557
052A
04E5
04E4
0501
04E3
049D
049C
04FC
053F
04EE
045B
0465
0543
05D7
048E
0118
FD12
FAA1
FA74
FB48
FB7F
FAD4
FA54
FAC5
FBA4
FBE1
FB44
FAA2
FAB0
FB26
FB48
FAF6
FAC2
FAFF
FB44
FB20
FAD5
FAFE
FB86
FB8C
FAB0
FA0D
FB5E
FEFE
032D
05A1
05B3
04BB
0461
04F1
0582
0565
04EC
04C4
0501
0523
04EA
04AD
04C6
0503
04FB
04BB
04BC
0520
0559
04EA
0446
046C
057B
0611
0490
00EE
FCFB
FAAD
FA63
FAF9
FB42
FB16
FAEE
FAFD
FAFE
FACB
FAAB
FAE2
FB41
FB5E
FB2B
FB09
FB3B
FB76
FB4A
FACD
FAA2
FB20
FBBC
FB90
FA97
FA15
FB86
FF07
02FE
0570
05B5
04DA
0460
04CC
056D
0574
04E4
0470
048F
0502
053B
0513
04D3
04B2
0494
045F
0454
04B5
0540
055F
0508
04EB
056D
05A0
03FD
004B
FC64
FA80
FADE
FBB9
FB8D
FAB7
FA83
FB2F
FBB2
FB5F
FAD7
FB04
FBAB
FBD4
FB45
FAD5
FB18
FB82
FB5C
FAF1
FAFF
FB62
FB31
FA76
FADA
FDBE
0220
0543
05AC
0494
0422
04D1
056E
0527
049B
04A5
0503
04D5
0416
03B1
0425
04D3
04F7
04BC
04CA
0520
0523
04C1
04BE
055F
0569
034D
FF42
FB7B
F9F4
FA79
FB4D
FB53
FAF8
FAFC
FB3A
FB20
FACA
FAEC
FBA4
FC27
FBDC
FB42
FB2E
FB90
FBA1
FB2B
FAE6
FB3E
FB75
FACA
FA20
FB76
FF58
03B6
05ED
059C
04A7
04AD
0557
0576
04F0
04B2
0510
0546
04C4
0420
042B
04AC
04C6
045C
0433
04A3
04FA
04A6
044F
04E8
05DB
0524
01C3
FD53
FA86
FA4C
FB31
FB74
FAED
FA97
FAE3
FB41
FB28
FAE1
FAF1
FB45
FB62
FB32
FB20
FB62
FB9A
FB74
FB31
FB45
FB8B
FB64
FAC9
FADD
FCEC
00C4
047C
062A
05B2
04A6
0468
04E8
0536
04ED
0493
04AF
0507
0510
04C6
0499
04B7
04D4
04C1
04BC
04E3
04DC
0474
0435
04BA
055D
045D
00E5
FC86
F9EA
FA00
FB30
FB88
FAE9
FA90
FB05
FB84
FB59
FAED
FAFC
FB61
FB6A
FB08
FAEF
FB60
FBAE
FB5A
FAF6
FB42
FBCB
FB7B
FA86
FAD5
FDD5
025B
0596
0614
050C
0484
04EA
0531
04C2
044E
0495
0533
0540
04AD
0453
04AC
052F
0522
04A1
0457
0478
0497
0488
04B7
0539
050D
02F4
FF23
FB86
F9F6
FA66
FB3A
FB44
FADB
FAEA
FB79
FBB8
FB46
FABD
FAD2
FB57
FB96
FB55
FB11
FB2E
FB72
FB76
FB4D
FB3C
FB2B
FADF
FADF
FC58
FFB0
0389
05D1
05D2
04C4
0440
0495
04F3
04D7
0499
04AC
04E4
04E3
04BB
04C1
04E9
04DD
049B
0486
04BB
04CA
0478
0456
04FD
05BA
04D6
0189
FD47
FA7B
FA1C
FB04
FB95
FB70
FB40
FB61
FB79
FB3C
FAFE
FB1E
FB61
FB4A
FAEA
FACD
FB1E
FB68
FB53
FB35
FB7B
FBCC
FB66
FA72
FA79
FCDD
0109
04AB
05EA
051F
041E
0420
04CD
052B
04FD
04CD
04F5
0529
0504
04A9
0482
04A6
04CE
04D1
04C9
04C2
0494
0459
0491
0564
05D1
0454
00A6
FC8E
FA53
FA7F
FB8C
FBD9
FB51
FAE7
FB00
FB14
FABF
FA6B
FAA0
FB25
FB58
FB2B
FB21
FB69
FB8C
FB46
FB0F
FB52
FB8E
FB04
FA37
FADB
FDDE
01F0
04B6
0543
04C0
04A5
0507
051B
04BF
04A5
0516
056E
0521
04A2
04C2
0566
059F
0508
045E
0474
04F8
0500
0482
0479
053F
0584
039B
FFA8
FBE7
FA69
FB06
FBDC
FB9F
FACB
FA83
FAFB
FB6B
FB4E
FAF7
FADF
FAEE
FAD7
FABA
FAF1
FB60
FB7B
FB27
FAFC
FB54
FB89
FAEC
FA43
FB6F
FF11
034B
0585
0539
043B
0445
050F
0546
04AB
0448
04BE
055D
055A
04F8
04FA
0552
054F
04D1
0481
04AE
04C1
0450
0413
04E3
05FF
0559
0209
FDBF
FB0A
FAAB
FB48
FB7D
FB46
FB45
FB77
FB55
FAD8
FA9E
FAEA
FB39
FB0D
FAB6
FACC
FB38
FB60
FB29
FB27
FBA5
FBFE
FB6E
FA5C
FA60
FCA9
0097
0429
05C7
0587
04B3
0460
049F
04E7
04E8
04D2
04E7
0510
0512
04F1
04E7
04F4
04DD
049C
047F
04A6
04C8
04AA
04A8
0528
058D
045D
00F6
FCD2
FA56
FA4C
FB37
FB60
FACA
FAA0
FB39
FBAA
FB41
FA99
FA9F
FB37
FB7D
FB2B
FAF1
FB43
FB9C
FB69
FB04
FB14
FB55
FB03
FA64
FB16
FE1E
0248
051C
0581
04A9
0454
04CF
052F
04F6
04AA
04CF
0523
0520
04DA
04CE
050A
0517
04BE
0469
048B
04E6
04F2
04C3
04F8
0591
055F
032D
FF5A
FBDD
FA69
FAD2
FB8D
FB80
FAFB
FAD4
FB25
FB58
FB1F
FAD9
FAE5
FB15
FB12
FAF3
FB0F
FB52
FB4F
FAF7
FACE
FB1C
FB56
FAED
FA8D
FBC0
FF0A
02E7
0536
0569
04C8
04A5
04FA
0504
04A2
046C
04B2
0506
0506
04EB
050E
0538
0503
04A1
04AD
052E
0569
04F6
0483
04E5
0593
04DD
01E5
FDEA
FB23
FA7B
FAFB
FB4E
FB30
FB27
FB59
FB5C
FB06
FAD3
FB2B
FBAF
FBAF
FB26
FAC1
FADF
FB14
FAE4
FA99
FAC9
FB46
FB36
FA87
FAA3
FD07
0135
04CB
05E4
04FE
0419
0454
0508
052C
04C8
0497
04CC
04EB
04B2
0489
04C4
050B
04EB
04A1
04C7
0545
055C
04D5
0485
0506
0565
03E5
003D
FC56
FA6F
FACB
FBBF
FBCF
FB1F
FAB5
FAF2
FB53
FB66
FB4C
FB3B
FB17
FAC7
FA9F
FAF8
FB8A
FBAC
FB3E
FAEA
FB2E
FB89
FB31
FA89
FB2C
FE1E
0241
0534
05C2
04EE
047A
04DF
053D
04EF
0474
0486
04FC
0518
04BF
049A
04FB
0550
0505
0476
0461
04BD
04CE
046F
0472
0536
0572
0362
FF31
FB47
F9D4
FA83
FB55
FB28
FAAE
FADC
FB6B
FB7A
FAFE
FAC8
FB33
FB9C
FB6C
FB06
FB14
FB70
FB6C
FB06
FAFE
FB96
FBEC
FB4D
FAAB
FBE8
FF82
0399
05D3
05C6
04FE
04D9
0528
0515
04A3
0490
0507
0550
04E9
0456
045C
04D8
0501
04A6
047B
04E9
0549
04DD
0422
0444
051F
04D4
01F2
FD93
FA74
F9FA
FAF1
FB60
FAEB
FAA8
FB20
FB92
FB4E
FAD4
FAF2
FB75
FB7E
FAF4
FAB2
FB32
FBC2
FB97
FB0C
FB11
FB95
FB8D
FABE
FAB6
FD0D
012D
04A5
05C5
0531
04A7
04E0
0537
0507
049E
0492
04D8
04FA
04E1
04E6
0521
0534
04E2
0484
0482
04B8
04B0
046C
0481
0525
0567
03E4
0070
FCA5
FA7F
FA74
FB42
FB7F
FB0C
FABD
FB01
FB5C
FB3D
FAE1
FAE5
FB50
FB8B
FB4F
FB07
FB1D
FB59
FB52
FB2C
FB51
FB8F
FB3E
FA8F
FB01
FDCE
0207
0528
05C2
04E5
0489
0527
05A4
0544
04A3
049C
04F9
04EF
0470
043D
04A2
04FF
04D0
0488
04C8
053F
051A
0475
045E
052B
056D
036E
FF75
FBCC
FA5B
FAC2
FB42
FAF7
FA82
FAAC
FB42
FB89
FB5F
FB3C
FB57
FB60
FB26
FB01
FB40
FB8B
FB53
FAC6
FAB5
FB5B
FBD1
FB4D
FA98
FB93
FEF4
031D
05A0
05BA
04CD
0483
0509
0568
051B
0497
0472
0499
04AD
04A6
04B2
04BF
049D
0478
04AD
051F
052D
04A4
0447
04DC
05BE
0522
021E
FDF9
FB05
FA4F
FAE5
FB4D
FB17
FACF
FAE5
FB2F
FB5D
FB73
FB89
FB82
FB48
FB1F
FB59
FBBE
FBB5
FB21
FAB2
FAFF
FB96
FB73
FA8E
FA62
FC7A
0081
044C
05F8
05A7
04EF
04D9
0510
04E2
0467
0436
0476
04B6
04B1
04A3
04BB
04B4
045D
0420
047E
0521
0533
04B0
049C
0566
05C3
03EB
FFF6
FC20
FA6F
FABB
FB55
FB45
FB04
FB39
FBA6
FBAE
FB59
FB1B
FB1A
FB27
FB3F
FB80
FBBA
FB9B
FB49
FB46
FB96
FB80
FABE
FA80
FC62
003F
03EB
0579
0538
04CA
04FB
053A
04F5
047B
045E
0496
04B4
04A4
04AC
04DB
04ED
04D2
04B9
0495
042A
03CE
044A
0575
059E
0343
FF12
FB7E
FA33
FAA1
FB2D
FB2A
FB0E
FB32
FB48
FB1F
FB12
FB56
FB8C
FB6E
FB53
FB7A
FB76
FAF9
FAAA
FB52
FC55
FC30
FAC6
FA44
FCCA
0185
0546
0615
0515
047D
04DA
052E
04F1
04AA
04C6
04F4
04DC
04A8
0493
0479
0442
0454
04F3
0576
0511
0443
0464
0564
052C
0228
FDA4
FA7D
F9EC
FAAA
FB15
FB0D
FB38
FB84
FB53
FAC2
FAA7
FB31
FB93
FB60
FB3C
FBA1
FBE1
FB50
FA91
FAAB
FB4D
FB3E
FA93
FB2C
FE50
029C
055F
05B5
0527
0526
0553
04D1
0416
0431
050C
058A
053A
04C7
04B9
04C1
0486
0461
04B0
0505
04CF
0481
04FC
05A3
0478
00C5
FC9A
FA9F
FAFB
FBA1
FB35
FA76
FA9C
FB73
FBDA
FB70
FAEA
FAD7
FAF8
FAF9
FB07
FB39
FB36
FAF4
FB06
FB9B
FBD5
FB13
FA78
FBF5
FFC7
03BE
058E
0532
0471
0472
04C5
04C0
04A0
04D0
0504
04D1
048B
04B6
0517
0522
04F1
0511
0560
0517
0434
03EA
04E0
059E
03E2
FFA6
FB94
FA08
FA96
FB48
FB49
FB36
FB78
FB93
FB3F
FB03
FB4E
FBA6
FB63
FAD1
FAB8
FB0C
FB03
FA95
FAB2
FB94
FBFE
FB2B
FA93
FC67
0098
048D
0615
05A1
050A
0510
0503
0484
0441
04B0
0526
04EA
0462
0460
04D0
050A
04F8
050D
053C
04F0
0442
0435
051A
0563
032A
FECB
FAF9
F9BF
FA71
FB14
FAF5
FAD7
FB3B
FB9E
FB83
FB31
FB1D
FB2B
FB08
FAD6
FAF6
FB43
FB44
FB09
FB21
FB84
FB68
FAB6
FAE7
FD69
0190
0501
062E
05B4
051E
050A
0504
04B7
0473
0481
04AA
04BB
04DE
052A
0549
0513
04E7
0505
0504
0485
0425
04BA
05B9
0533
0206
FD93
FA85
F9FE
FABB
FB12
FAD3
FAC3
FB1D
FB6A
FB76
FB76
FB78
FB45
FAF1
FADD
FB16
FB25
FADB
FAC3
FB46
FBAC
FB0B
FA1C
FB04
FEAD
032F
05C7
05CC
04E7
04A3
04E7
04EB
04A6
04A3
04E4
04E9
04A4
0499
04ED
0510
04C4
049A
04EB
0521
04B8
0460
0502
05DB
04CE
0105
FC6F
F9DF
FA00
FB12
FB6B
FB2F
FB3D
FB8E
FB86
FB2B
FB0F
FB49
FB64
FB39
FB1E
FB35
FB2A
FAE8
FAEF
FB72
FBA3
FADA
FA2E
FBBB
FFDB
0425
05FC
0568
0484
04A6
0531
0523
04A1
0473
04BB
04EA
04C1
049F
04AF
04A8
047B
048F
04F0
0507
04A7
049D
055C
05A5
03AD
FF8B
FB9E
FA10
FAA0
FB6E
FB67
FB13
FB1B
FB36
FAF9
FAC1
FB07
FB79
FB7B
FB2E
FB24
FB5F
FB66
FB34
FB49
FB9D
FB63
FA78
FA6D
FCF8
016F
04FD
05C3
04D2
0454
04CF
052A
04CD
046C
04AF
0535
0554
051E
050C
0513
04D1
0474
0486
04E1
04BF
0433
0459
055E
0566
02A2
FE06
FAA1
FA32
FB64
FBE2
FB35
FAA9
FAFF
FB77
FB46
FAD2
FAC9
FAF8
FAD2
FA8D
FAB8
FB33
FB65
FB47
FB5A
FB95
FB4D
FA9C
FB10
FDFF
0267
058C
05EF
04C6
041D
046D
04CD
04B7
0493
04B8
04ED
0502
0524
056C
0586
053C
04EA
04F2
050D
04C3
0471
04D9
0580
0493
012A
FCE7
FA5C
FA42
FB24
FB86
FB63
FB6C
FBAF
FBB5
FB70
FB45
FB39
FAE4
FA60
FA5D
FAFD
FB6C
FB31
FAF4
FB53
FBA0
FAF5
FA27
FB56
FF2F
0396
05CF
057C
048B
0476
04CC
04AE
045B
047C
04CF
04AA
0448
047C
0545
05AE
0539
0492
0475
04A4
0491
0490
0537
05BC
0444
0060
FC36
FA3C
FA87
FB49
FB5F
FB3C
FB7F
FBCF
FB9F
FB35
FB3B
FB99
FB9A
FB1C
FACC
FAFE
FB34
FB1E
FB35
FBAA
FBB5
FADD
FA69
FC3B
0045
0421
05A9
0531
049A
04CC
0509
04AC
0440
046C
04CF
04BA
0460
046A
04CD
04F2
04C0
04AF
04D4
04B5
044D
0462
052F
054A
0300
FECC
FB51
FA6C
FB38
FBAB
FB3A
FAE7
FB42
FBA1
FB68
FAFA
FB00
FB5C
FB79
FB47
FB40
FB76
FB7B
FB42
FB4A
FB97
FB6C
FAB4
FAE9
FD78
01A3
04F4
05DF
0530
049B
04B0
04CC
0489
045B
049B
04EA
04E5
04C5
04DE
04FA
04D3
04A7
04C0
04D2
0483
044D
04E3
05BA
0501
01BC
FD65
FA97
FA40
FAF2
FB19
FAC6
FADE
FB6A
FBBA
FB95
FB68
FB5E
FB35
FAEA
FAE3
FB39
FB63
FB1B
FAF5
FB75
FBEC
FB51
FA42
FAFA
FE85
0303
05A7
05C4
04F6
04B4
04DF
04D3
04AB
04D6
0516
04D8
0453
0460
050C
0565
04F7
0487
04B7
04F1
0487
0425
04CB
05B6
04B6
00F8
FC86
FA26
FA4C
FB20
FB38
FB05
FB4B
FBA3
FB58
FACE
FADE
FB5F
FB70
FAF4
FABC
FB20
FB72
FB34
FAFA
FB6A
FBE3
FB63
FA98
FBAD
FF68
03B0
05DB
05A7
04E5
04D0
04FE
04D2
049D
04E2
0542
0512
0488
047D
050B
0558
04F7
0490
04AC
04D7
049B
0484
050F
053E
0368
FF91
FBE4
FA5F
FAC1
FB4E
FB2C
FAF4
FB2F
FB5F
FB0D
FAB2
FAE3
FB49
FB40
FAF2
FAFE
FB58
FB6B
FB31
FB48
FBBC
FBB0
FAD4
FA9D
FCD4
010B
04A4
05BC
051B
04A7
04EA
0522
04FB
04F8
0547
0557
04E1
0482
04CC
0545
051B
0478
0443
04A0
04B9
0456
045E
051E
050D
028B
FE58
FB15
FA4C
FB00
FB68
FB20
FAF3
FB27
FB21
FAAD
FA7F
FAFB
FB73
FB3B
FAC2
FACE
FB41
FB7A
FB78
FBB0
FBF0
FB7E
FAA5
FB1D
FE1D
0268
0554
05C0
0505
04CF
051A
0507
049D
04A0
051D
054F
04EB
0490
04C0
051C
0514
04D0
04C4
04C9
046E
040F
0483
055C
04B0
016C
FD24
FA81
FA4A
FAFA
FB0F
FAB1
FAC4
FB44
FB6C
FB13
FAE7
FB3E
FB8C
FB59
FB09
FB15
FB45
FB34
FB22
FB65
FB91
FB16
FAA3
FBE7
FF73
038B
05CA
05B3
04E3
04CE
0531
0521
04A1
046D
04B1
04EA
04D0
04B1
04CB
04EF
04ED
04DF
04DB
04B6
0472
048E
0539
0570
03AF
FFEC
FC20
FA4B
FA6B
FAFF
FB0D
FAE3
FB08
FB4E
FB44
FB04
FAFC
FB3A
FB5D
FB39
FB0F
FB0A
FB09
FB12
FB64
FBCB
FB93
FAB6
FA99
FCB9
00AE
043F
05A4
053D
04B7
04EF
0555
0537
04CC
04AA
04DF
0513
051F
0515
04E9
04A3
0497
04FA
055A
0519
0471
0456
04FD
050C
02F6
FF18
FBA9
FA5C
FABA
FB34
FB1B
FAE4
FAF1
FB06
FAED
FAE5
FB1E
FB4F
FB27
FAE9
FB08
FB61
FB67
FB1C
FB1C
FB82
FB86
FAD5
FAAE
FCB1
00AA
045F
05E1
056F
04BD
04C8
051F
0517
04D8
04DC
050D
0500
04BF
04AB
04CC
04C7
048D
0487
04D8
0505
04AB
0454
04D8
05F1
05FD
03A9
FF9C
FBFF
FA71
FABE
FB89
FBCA
FB72
FAF8
FAB9
FAC1
FAF7
FB37
FB58
FB47
FB21
FB1C
FB41
FB58
FB31
FAF1
FAE8
FB23
FB3C
FADF
FA8D
FB82
FE6F
025C
0535
05C1
04C1
03F2
0432
04ED
0545
0529
0516
052D
051B
04CE
04A7
04CB
04DF
04AD
049A
04FB
055D
0511
045E
0456
0524
0535
02E1
FEC1
FB6A
FA9C
FB79
FBF7
FB6B
FAD7
FB00
FB58
FB0F
FA6A
FA52
FAF0
FB82
FB8E
FB74
FB92
FB86
FAF2
FA68
FABF
FBA3
FBC3
FAC6
FA4F
FC45
0051
03F4
0535
049E
0423
04A0
0543
0524
049B
048E
0519
057E
0541
04B9
046D
0460
0457
0469
04D4
0555
054B
04AE
045C
04F0
0594
0490
014A
FD49
FACB
FA92
FB61
FBAA
FB33
FACF
FAF8
FB43
FB33
FAF1
FAF1
FB34
FB58
FB42
FB3E
FB63
FB5D
FB06
FAD8
FB41
FBC2
FB69
FA6C
FA82
FD17
0159
04C2
05B0
04EB
0455
04AA
0526
0510
04C7
04E8
053C
051A
048A
044C
04B6
052D
0514
04B9
04C5
0519
04FA
0461
044B
052C
05B5
03FE
FFFB
FBF9
FA40
FABE
FB8C
FB5A
FAAE
FA97
FB11
FB42
FAE5
FAA4
FB00
FB8A
FB94
FB33
FB09
FB3D
FB51
FB03
FAD2
FB2D
FB93
FB3F
FA9E
FB55
FE5F
0285
0559
05B8
04CB
0468
0501
0594
0559
04BD
0497
04F9
0545
051D
04C2
0482
0459
0446
048E
0536
05A3
0543
0487
0485
0554
0559
02F5
FEB1
FB0E
F9EB
FAAC
FB5A
FB0F
FA92
FAC5
FB55
FB67
FAEE
FAA6
FAE6
FB40
FB55
FB64
FBA3
FBA3
FB00
FA48
FA72
FB59
FBA1
FAA9
F9F8
FBC0
000A
0441
05F2
0558
0493
04DF
057E
055A
04B5
0497
0527
057E
050C
0468
0459
04BE
04EA
04CB
04E5
054C
0560
04DC
048A
052B
05F4
04F5
0166
FCF5
FA3E
FA24
FB39
FBA7
FB21
FAA2
FACC
FB3C
FB56
FB24
FB0D
FB29
FB2F
FB07
FAE7
FAE8
FAD8
FAB1
FACD
FB58
FBBD
FB4A
FA6D
FAC5
FD74
0198
04E9
05EB
053D
0489
04A6
051B
0530
04D9
0481
045F
046B
04AE
0525
057B
0550
04D6
04BA
0537
0599
0526
044F
0447
053C
0596
0398
FF91
FBC6
FA27
FA82
FB3C
FB4D
FB05
FB07
FB4A
FB5B
FB35
FB35
FB6D
FB7E
FB36
FAEA
FAF1
FB16
FAF4
FAA9
FAC2
FB51
FB90
FAF1
FA47
FB51
FEC4
0324
0601
0648
0516
043E
046B
04E9
04F3
04A8
0498
04D7
04FA
04CC
0493
049A
04C8
04E3
04ED
04FF
04F1
049B
0456
04BB
0589
054B
02BA
FE7A
FADF
F9AC
FA6E
FB56
FB5C
FAFA
FAFB
FB4D
FB63
FB2E
FB21
FB60
FB81
FB4B
FB15
FB33
FB5F
FB41
FB21
FB7C
FBFB
FBA9
FA7C
FA18
FC3F
008C
0481
060F
058C
04CE
04DE
0535
0510
049B
0479
04B4
04CC
0497
0482
04CB
050B
04D7
0474
0472
04C1
04BC
0448
042D
04FA
05BC
04A3
0111
FCB0
F9FE
F9E6
FB1C
FBCB
FB70
FADC
FACD
FB1D
FB4C
FB44
FB47
FB60
FB54
FB24
FB20
FB68
FB9E
FB75
FB41
FB79
FBCC
FB6B
FA7B
FA9F
FD51
01D3
0575
0646
0504
03F7
0442
0512
0542
04E5
04C1
04F3
04EB
0487
045C
04BD
0525
0503
049E
049A
04D7
04A4
0412
042C
0548
05D2
03CC
FF74
FB73
FA14
FAEA
FBC3
FB6E
FAB6
FAB3
FB32
FB4F
FAFB
FAF4
FB78
FBD2
FB76
FADD
FACF
FB36
FB5B
FB1C
FB24
FBB4
FBF6
FB2D
FA43
FB3B
FEC4
0314
0599
05A1
04B4
0482
051A
0573
051C
04B5
04CD
0513
04F8
0497
047C
04BC
04D6
0499
047D
04D7
0528
04CE
0427
0447
0538
054B
02D8
FE83
FAF0
F9FD
FAF2
FBB6
FB60
FAC2
FAC3
FB19
FB09
FAB3
FAD8
FB8B
FBFB
FBAB
FB25
FB19
FB58
FB49
FB04
FB31
FBBC
FBAF
FABD
FA63
FC72
00A1
0464
05A7
04ED
043E
048B
0502
04CD
0466
04AB
0564
0588
04D2
0427
0440
04AA
04A2
045D
049D
0550
0576
04B6
0425
04C5
05AD
04AB
00FD
FC98
FA31
FA64
FB7D
FBC6
FB4E
FB15
FB5D
FB83
FB33
FAF3
FB35
FB97
FB78
FB05
FAFE
FB8B
FBF2
FBA8
FB1E
FB09
FB3A
FAEC
FA4D
FAE3
FDD3
0222
0550
05E5
04D4
041F
0490
0544
0534
0487
041A
044E
04BD
04F1
04E9
04D0
04A7
0470
0467
04A7
04E0
04B9
0480
04E3
05C3
05BE
037E
FF72
FBBF
FA2C
FA7F
FB21
FB16
FACB
FAFA
FB7E
FBA3
FB41
FAEA
FB07
FB4A
FB42
FB0E
FB0F
FB39
FB2E
FB00
FB36
FBD3
FBEA
FADE
F9C7
FAC7
FE95
033D
05F2
05EA
04DE
04AB
0551
058C
04E7
043F
0463
04FC
0537
04FD
04D8
04F8
04F9
04BA
04B9
0538
058C
0502
041E
042B
0546
059F
0361
FF0E
FB3F
F9EE
FA91
FB41
FB12
FAB3
FAF2
FB86
FBA0
FB2B
FACD
FAEB
FB38
FB46
FB20
FB05
FAF3
FAD5
FAE5
FB5D
FBD4
FB7C
FA6C
FA1F
FC20
001D
03E1
0579
050D
0452
0474
0514
0546
04ED
04A5
04C3
04F9
04FA
04F2
0515
0530
04FA
04AC
04BC
0513
050C
047F
043B
04E7
05A3
049A
0136
FD31
FAEB
FAEE
FBAE
FBA2
FAF1
FAB5
FB3C
FBB6
FB81
FAF6
FABB
FAD4
FADE
FADA
FB1A
FB8B
FBA9
FB58
FB32
FB99
FBE0
FB2C
FA15
FA8E
FDB5
0222
051D
056C
045B
03EB
049E
0561
0546
0498
0438
047A
0502
0566
0585
055C
04EF
0478
044F
0470
046B
0409
03DA
048D
05BF
05D2
0377
FF4C
FB92
FA1C
FAB4
FBAB
FBBA
FB15
FAB6
FB0C
FBA2
FBD3
FB7F
FB02
FAB3
FAAC
FAE1
FB33
FB72
FB80
FB87
FBC6
FC0F
FBD0
FAE3
FA4A
FB8A
FF00
0317
0596
05BB
04C8
0466
04EC
0576
0555
04D0
0480
0480
0485
0482
04AF
0501
051A
04DB
049D
04A2
04A3
044E
0404
0470
053C
04E4
0245
FE44
FB34
FA7F
FB4D
FBC3
FB2A
FA60
FA5E
FAFB
FB64
FB4F
FB2C
FB50
FB7B
FB56
FB04
FAEC
FB22
FB5B
FB6D
FB7B
FB83
FB4B
FAEA
FB3D
FD36
009B
03D4
0552
0508
044B
044A
04F5
0574
0553
04E7
04B2
04CC
04FA
0513
050F
04EF
04C4
04BD
04EC
0505
04AF
0428
0432
0500
0579
0415
00AD
FCF8
FAEC
FAD9
FB74
FB8E
FB2A
FAEA
FAED
FADE
FAB7
FADE
FB56
FB84
FB0D
FA87
FAB6
FB6B
FBB2
FB3E
FAEA
FB74
FC3B
FBFE
FADF
FABE
FD26
0145
049D
059F
0502
0477
04B8
0530
0538
04F1
04D5
04ED
04EB
04BE
04A6
04BC
04C5
0499
0473
04A3
0510
0542
04F8
048A
048B
050A
053F
041D
014F
FDC0
FB0B
FA38
FAEA
FBCB
FBE3
FB5F
FB0B
FB38
FB71
FB40
FAD7
FAC5
FB2C
FB98
FBA0
FB6A
FB49
FB37
FAEE
FA82
FA70
FAF1
FB88
FB93
FB58
FC0A
FE88
022A
0520
0615
055E
046D
0447
04B4
04E6
049F
0463
04A2
050E
050A
0488
0423
044E
04C1
04E8
04BE
04C5
0525
0552
04DC
0444
0468
0507
0481
01A4
FD6C
FA58
F9DB
FAF5
FB98
FB0B
FA5E
FAA3
FB7C
FBCF
FB5F
FAF9
FB37
FBAC
FBA8
FB40
FB1D
FB6E
FBA3
FB56
FAF7
FB1E
FB93
FB81
FAB8
FA59
FBCD
FF35
0312
058C
05FA
0538
049F
04CE
055F
058E
051D
0486
045B
0499
04C5
04A2
047B
04A2
04D8
04A8
042C
041C
04CB
058D
0582
04D3
0476
0499
03F2
0144
FD4B
FA5D
F9EB
FB01
FB99
FB01
FA53
FA92
FB50
FB7F
FB08
FAC7
FB28
FB93
FB6C
FB16
FB52
FBFC
FC13
FB29
FA2B
FA44
FB4C
FBF7
FB90
FB0C
FC07
FEF3
0287
04FF
05AD
0541
04D1
04D8
0516
0525
04F4
04C6
04CB
04E8
04E7
04C4
04A7
049B
047B
0447
044E
04C5
0551
0549
0499
0410
0467
050A
0464
0199
FDC2
FAF9
FA47
FAD9
FB3D
FAFE
FABD
FAFE
FB6B
FB71
FB17
FAE6
FB14
FB41
FB1A
FADB
FAFE
FB7E
FBCC
FB88
FB10
FB0A
FB7F
FBBB
FB46
FAC9
FBA7
FE83
0253
052A
05F8
0561
04CA
04DB
051D
04F5
0487
0461
04A5
04E6
04E1
04DA
0515
0546
04F7
0454
041A
0493
050E
04CC
0424
0431
0532
05CD
0455
00BC
FCD4
FA8E
FA46
FAE2
FB46
FB3C
FB22
FB2C
FB46
FB60
FB80
FB93
FB64
FAF4
FAA4
FAD9
FB77
FBEA
FBBE
FB28
FAD5
FB22
FBA6
FB9E
FAE9
FA86
FBD3
FF26
0321
05C1
061B
0511
0440
045D
04D7
04E0
047A
043B
046C
04B9
04C9
04B5
04C1
04D4
04A3
0448
0449
04DC
056D
054A
049E
045F
04F3
0556
03FB
009B
FCC4
FA6E
FA26
FAD9
FB41
FB24
FB18
FB73
FBD9
FBD3
FB74
FB23
FB12
FB1B
FB29
FB64
FBCB
FBEE
FB65
FA81
FA25
FAC3
FBA7
FBBB
FAEC
FA97
FC35
FFB6
0364
0573
0594
04EA
04A3
04E5
0512
04C6
0449
0420
0462
04BB
04E4
04E2
04D5
04B6
047A
0457
049F
0539
0590
052D
0470
0442
04E5
053C
03BE
0034
FC4D
FA2B
FA5A
FB7C
FBE6
FB4F
FAAE
FAC7
FB50
FB96
FB7A
FB70
FBA8
FBB8
FB4F
FAC3
FAB2
FB1A
FB5C
FB21
FAE1
FB30
FBBF
FBAB
FAD7
FA8D
FC4C
FFF9
03AA
0572
052A
044A
042A
04C2
052F
0505
04AD
04A4
04C2
0499
0432
041C
04A4
0551
0572
0501
04A3
04C2
04FA
04B3
041E
0418
04E7
0568
0406
0092
FCC6
FAA7
FA98
FB48
FB69
FB05
FAF7
FB7A
FBDC
FB93
FB0B
FB04
FB77
FB9D
FB1B
FA90
FAC4
FB82
FBD5
FB58
FACE
FB1A
FBEF
FC22
FB4B
FAA0
FBD1
FF20
02EC
0543
05A2
0513
04C3
04DA
04CA
0459
03F9
0426
04B3
0509
04F2
04D6
050D
0549
04FF
0447
03E8
0454
04EF
04D2
041A
03EA
04CE
0589
042C
006F
FC5D
FA56
FAA5
FB97
FBAF
FB28
FB1A
FBB7
FC15
FB9B
FAE3
FAD5
FB60
FBA6
FB43
FAD8
FB16
FBBB
FBED
FB6F
FAFE
FB42
FBD4
FBC0
FAF3
FABB
FC7F
001C
03C1
0595
055D
0476
0436
04A4
04E1
0486
042B
0479
0528
0554
04B6
040E
041E
04A0
04BB
044D
0427
04C8
057C
0544
0459
0401
04B4
0512
0355
FF98
FC01
FA80
FAE4
FB80
FB53
FADC
FAF3
FB7B
FBAF
FB51
FAFB
FB3B
FBCB
FBFE
FBAF
FB61
FB78
FBB3
FB93
FB15
FAC3
FAFD
FB70
FB74
FB0A
FB39
FD1F
009C
040F
05BD
0571
048E
0478
0523
0579
04ED
042E
0423
04A9
04DA
045C
03E0
0423
04E1
0530
04C6
044C
0458
049F
048A
0444
0485
0541
0524
02E1
FEF3
FB73
FA19
FA9E
FB5E
FB48
FAC6
FAC2
FB58
FBD0
FBB5
FB64
FB6E
FBC1
FBCB
FB5C
FAEE
FAFF
FB5B
FB72
FB34
FB2C
FBA5
FC0A
FB9B
FAAC
FAC6
FD1A
0111
049D
0620
05C9
04FD
04C2
04F2
04EF
0496
044C
0456
047D
0478
045F
047E
04CC
04E6
049D
0457
048E
051E
0548
04A9
03E6
0400
04EB
0526
0328
FF33
FB64
F9BC
FA43
FB53
FB83
FAFA
FABE
FB37
FBC7
FBC8
FB65
FB37
FB65
FB86
FB5F
FB36
FB57
FB86
FB51
FAD3
FAB5
FB50
FC02
FBE5
FB1C
FB13
FD23
00FE
04B2
0663
05EC
04C4
0454
04B5
0509
04CB
0458
0442
047F
0492
0459
0443
0496
04FB
04F7
04B5
04CB
053D
054F
0498
03DA
0423
051E
04F9
025C
FE36
FAFA
FA1B
FAC7
FB3F
FAE9
FA98
FB0B
FBDE
FC2F
FBCB
FB55
FB54
FB98
FBA7
FB70
FB45
FB4A
FB4C
FB20
FAFE
FB35
FBA5
FBBB
FB28
FA8B
FB2F
FDD4
01AE
04D4
05E4
0542
0486
04BF
057A
059E
04EB
043C
044B
04C1
04C8
0447
03F7
044E
04D7
04DB
0467
042E
0479
04C2
048E
0446
04A3
0563
0513
0292
FE8E
FB2A
FA02
FABA
FBA5
FB97
FAEA
FAA2
FB0D
FB7D
FB50
FACB
FAB5
FB40
FBC9
FBB6
FB4C
FB47
FBC6
FC1E
FBD9
FB66
FB6B
FBBA
FB84
FAC3
FAD5
FD1B
0121
04B3
0602
0554
045E
0451
04EC
0559
054D
0513
04E7
04BB
0497
04B3
050F
0538
04CB
0414
03CA
042E
04AF
049A
040C
03E6
04B4
05BB
055F
02B3
FE9A
FB37
FA0D
FAB3
FB78
FB3F
FA7E
FA55
FAFA
FB8A
FB5E
FAED
FB10
FBB2
FBE7
FB50
FABD
FB12
FBF2
FC2A
FB68
FABC
FB1B
FBEA
FBD1
FAD6
FACC
FD46
0176
04D2
05B6
04ED
0467
04F3
05B9
05B9
0512
04A1
04C0
04F4
04C9
0475
0474
04C0
04D7
0485
043D
0475
04F1
0500
0487
0446
04D7
0591
04DD
01F8
FE08
FB31
FA86
FB2F
FB9C
FB39
FAA8
FA9B
FAE8
FB02
FAD9
FAE0
FB4B
FBAF
FB9E
FB51
FB55
FBB4
FBD6
FB5D
FAC5
FAD1
FB76
FBC1
FB12
FA3D
FAFB
FE14
0247
054A
05E5
04F0
0434
048D
0550
0578
04F5
0493
04CB
0523
04F3
0457
040E
0461
04BF
0490
0422
0444
0508
0589
0524
0479
049E
055F
0501
0230
FDDD
FA95
F9EA
FAFC
FBC3
FB5E
FAA4
FAA0
FB2D
FB6C
FB17
FAD1
FB1E
FBA8
FBCA
FB85
FB6C
FBBD
FBFA
FBA6
FB06
FACA
FB10
FB31
FAC2
FA7A
FBA7
FEAE
0258
04D6
0566
04D9
047F
04CF
053E
0531
04C5
0486
04A8
04D5
04C4
04A8
04D4
0522
050F
048A
042D
0475
04F1
04C3
03F0
03A1
0498
05CD
0529
01DE
FD8D
FABC
FA58
FB29
FB8D
FB2E
FACB
FAE6
FB3E
FB67
FB5F
FB5D
FB63
FB4A
FB18
FAFC
FAFD
FB02
FB0C
FB3E
FB87
FBA2
FB8B
FB94
FBCD
FBBE
FB18
FAA7
FBD1
FEFB
02B0
04F5
053A
04A6
0471
04B0
04D8
04D3
04F8
053F
0538
04CD
0486
04C5
0529
051A
04B1
048D
04D4
04FA
04AB
0452
0461
048A
0459
0421
048D
0537
0480
0173
FD53
FA93
FA46
FB38
FBB2
FB63
FB19
FB39
FB54
FB1C
FAE2
FB01
FB40
FB3A
FB06
FB06
FB35
FB37
FB07
FB15
FB84
FBD4
FBAB
FB6F
FB8F
FBA9
FB1B
FA79
FB75
FEE3
0343
0601
061E
04EF
0443
046F
04AE
0498
0488
04BA
04E2
04C4
04A3
04CC
0514
0519
04E4
04CA
04D0
04A7
0453
0443
0494
04C5
0492
0491
053E
05AF
0426
0042
FBFD
F9D6
FA41
FB83
FBEB
FB80
FB37
FB5F
FB7C
FB4A
FB13
FB0F
FB0E
FAF8
FB10
FB7C
FBDA
FBB6
FB47
FB27
FB6B
FB8A
FB49
FB19
FB38
FB21
FA82
FA5C
FC41
0038
042D
05F6
058A
04A8
0497
04F8
04F0
0492
048B
04EE
0523
04DE
0483
0477
049C
04A8
04A6
04C0
04D9
04B8
048E
04B6
04FE
04D3
044E
045C
054E
05C0
03E0
FFC8
FBD3
FA30
FAB4
FB7D
FB60
FAE3
FAEC
FB59
FB78
FB2D
FAFC
FB1B
FB3A
FB2B
FB2B
FB65
FB92
FB70
FB3A
FB4F
FB8B
FB83
FB4A
FB60
FBB3
FB77
FA84
FA47
FC68
0090
0459
05B9
0510
0449
047D
0510
051D
04BE
049A
04C8
04DB
04B8
04B5
04EC
0504
04C6
0481
048A
04B4
04A8
047E
048C
04B8
0490
0439
0477
0560
058C
0371
FF72
FBDB
FA83
FB00
FB8F
FB47
FAC3
FACF
FB40
FB76
FB61
FB64
FB8E
FB8A
FB41
FB05
FB0C
FB22
FB19
FB20
FB60
FB92
FB66
FB2A
FB6C
FBEE
FBBA
FAAF
FA62
FC88
00BC
0488
05E5
052F
0448
0452
04D6
0500
04C4
0496
0490
047D
046A
0493
04E4
0504
04DD
04BC
04C9
04D0
04AB
049C
04D2
04E6
046E
03EA
0459
0581
0581
02CD
FE5B
FAF2
FA43
FB55
FC14
FBC0
FB3A
FB4B
FB9B
FB85
FB2A
FB15
FB4A
FB59
FB29
FB19
FB4A
FB66
FB36
FB04
FB1E
FB4E
FB41
FB2B
FB76
FBDB
FB93
FACF
FB23
FDCD
01D6
04CA
0553
0477
040A
0487
04FB
04B9
043B
043B
04AB
0504
051F
052A
051E
04D2
0476
0471
04C2
04EE
04C2
04A6
04E9
0514
049C
03FA
0431
050F
04CC
0216
FDFF
FB11
FA89
FB4A
FB9E
FB43
FB21
FB9D
FC0C
FBD7
FB50
FB0C
FB04
FAE5
FAC3
FAF1
FB4F
FB6C
FB45
FB4A
FB94
FBA1
FB35
FAF6
FB81
FC39
FBE4
FAB5
FAB7
FD77
01D6
0511
05B9
04E9
0473
04BC
04EE
049D
0457
0496
04FF
0508
04CF
04BF
04D6
04CA
04A8
04B6
04DC
04B5
044D
0433
0499
04DE
047B
040F
0496
0597
0516
01F1
FD9D
FAC9
FA76
FB49
FB90
FB2C
FB03
FB5D
FB92
FB40
FAE4
FB05
FB65
FB81
FB63
FB6B
FB96
FB89
FB48
FB36
FB6F
FB8B
FB54
FB2D
FB66
FB83
FAF1
FA5D
FB73
FECD
02D0
0534
0568
04C4
049E
04E9
04F7
04BA
04B5
04FB
0509
04AB
045A
0474
04A8
048B
0455
0474
04C1
04BE
047F
049D
0528
0552
04A5
03FF
0473
0562
04AF
0159
FD10
FA82
FA70
FB51
FB8B
FB23
FAF7
FB35
FB4A
FB09
FAFA
FB67
FBD5
FBC2
FB6A
FB53
FB78
FB74
FB43
FB3F
FB6C
FB67
FB21
FB18
FB7F
FBAB
FB0C
FA85
FBD5
FF61
034E
0561
0557
04B5
04A9
04F0
04E2
049F
04B6
050D
0503
047B
0422
046B
04E9
050A
04E8
04E5
04EB
04A9
0454
0478
04F6
0500
045E
040A
04CC
058F
0437
005B
FC3F
FA66
FAE2
FBB8
FB8E
FAE8
FACD
FB32
FB5E
FB2D
FB26
FB68
FB6D
FB02
FABD
FB08
FB6A
FB49
FAF3
FB1D
FBAB
FBC7
FB49
FB0B
FB8E
FBF9
FB5D
FAA4
FBEE
FFC4
03EB
05C3
052D
043D
0468
0525
054F
04E4
04AE
04E4
04F3
04A5
0482
04DC
0538
0513
04B7
04B2
04EB
04EB
04BF
04DC
0523
04E3
0412
03C7
04B0
0580
0407
0000
FBD1
F9F4
FA5B
FB1C
FB17
FADD
FB21
FB79
FB36
FAA8
FAB7
FB6E
FBDD
FB7E
FAF1
FAEB
FB33
FB34
FB02
FB14
FB4B
FB1F
FAB7
FAE3
FBBD
FC22
FB4B
FA7F
FC05
002C
047B
064C
059F
048F
0488
0519
0548
050E
04F7
0511
04FA
04B7
04BC
050E
0519
04A9
045F
04B4
052D
051D
04BD
04C5
0524
0506
044E
040B
04DD
056A
03A3
FF86
FB9C
FA34
FAEF
FBB8
FB79
FAEC
FAEA
FB28
FAF7
FA7B
FA6B
FAE5
FB4B
FB48
FB36
FB5B
FB6D
FB33
FB10
FB57
FB9B
FB4F
FADA
FB21
FBFE
FC24
FB13
FA70
FC5F
00A8
0485
05B3
04D0
0410
046F
050F
0510
04CB
04F6
0568
056F
04FA
04A7
04BA
04CA
0494
0478
04C2
050C
04E9
04A6
04C8
050D
04C2
0416
041E
051A
0567
0327
FED3
FB26
FA29
FB19
FBCB
FB63
FAD2
FB03
FB97
FBC0
FB74
FB42
FB4D
FB3D
FAFE
FAF8
FB49
FB74
FB26
FACC
FAE6
FB3C
FB46
FB24
FB63
FBE5
FBCE
FAFE
FAED
FD32
0151
04D4
05EE
053E
049C
04C4
04F9
04A2
0432
044A
04B6
04CD
047E
0455
048E
04C9
04C4
04C3
0504
0539
0509
04BA
04C2
04F5
04C5
044C
0459
0506
04ED
0291
FE72
FAF7
F9ED
FAC2
FB9B
FB91
FB35
FB32
FB67
FB6E
FB5E
FB82
FBB5
FB9A
FB49
FB42
FB98
FBBB
FB5D
FAF4
FAFC
FB38
FB26
FAEF
FB1F
FB94
FB83
FAE7
FB33
FDCA
01EC
0519
05BC
04C9
043D
04B9
0541
0508
0476
0452
049F
04CC
04A4
047B
048B
04A4
0497
047D
046A
0447
0433
048A
0535
0572
04D5
0429
047F
0568
04EB
01D4
FD89
FABD
FA80
FB62
FB9F
FB2F
FB1D
FB99
FBCE
FB54
FAD8
FB06
FB8A
FBAD
FB6D
FB5C
FB98
FBA3
FB53
FB2D
FB7C
FBBA
FB71
FB1B
FB60
FBDA
FB8C
FABA
FB39
FE4B
02A1
057B
05A7
0492
0430
04B6
050F
04BF
0462
0476
04AD
04A4
0491
04CB
050A
04CE
0442
0419
047B
04C9
04A6
0488
04CE
04F4
0464
03AD
03E6
04CE
047D
01A2
FD76
FAAE
FA7C
FB8A
FBF3
FB70
FAFB
FB0D
FB29
FAFA
FAE3
FB40
FBB8
FBC1
FB75
FB5B
FB8F
FBA8
FB7C
FB66
FB98
FBBD
FB92
FB6C
FB9B
FBB2
FB2E
FAAD
FBBF
FEFE
02F0
055B
0586
04B3
0455
0496
04D3
04D5
04EA
0521
0527
04E9
04BB
04C3
04B0
044D
03F1
040E
0475
049C
0477
0484
04DA
04D8
0432
03B6
043F
0518
045D
013F
FD48
FAD6
FA9E
FB43
FB4F
FAD6
FAC7
FB52
FBAD
FB5A
FAD5
FACD
FB32
FB6B
FB40
FB20
FB71
FBF9
FC2B
FBEE
FBA7
FBA0
FBA6
FB73
FB33
FB49
FBA3
FBA4
FB0B
FAB1
FBF7
FF34
02F0
0528
0540
046F
042D
04AA
051B
0519
0513
0564
0593
0509
041B
03C5
0457
04F9
04D9
043F
040D
046B
04A0
0445
03F3
045F
052E
0558
04A5
041F
04A1
055D
0482
015C
FD62
FAD0
FA7D
FB56
FBD0
FB77
FAF2
FAD9
FB07
FB11
FAFB
FB20
FB85
FBC2
FB96
FB50
FB63
FBBC
FBD7
FB85
FB36
FB55
FB9C
FB7F
FB13
FB0D
FB9D
FBF2
FB55
FA8E
FB6C
FEA5
02B3
053B
057A
04BB
0484
04EA
0507
048F
0433
047F
050B
051E
04B9
0483
04C5
04FF
04B2
0428
0415
0496
050A
04EF
0492
0486
04C2
04B7
043F
0406
049A
054A
0482
0184
FD8A
FAC5
FA46
FB2B
FBD7
FBAC
FB43
FB3E
FB71
FB5D
FB07
FAF0
FB3C
FB79
FB4C
FB02
FB25
FBA6
FBE7
FB9A
FB32
FB3B
FB96
FBA9
FB56
FB2A
FB87
FBF4
FBC2
FB42
FBCE
FE44
01CC
0484
0553
04DB
0479
04C4
053F
0550
0507
04D0
04CA
04C4
04AC
04B4
04DE
04DA
047B
041B
0433
04A5
04D0
0472
041A
0465
0503
0510
045D
03EB
0491
0580
04C7
018C
FD52
FA9C
FA65
FB63
FBCE
FB4F
FAE2
FB26
FB8B
FB49
FA9A
FA70
FB20
FBE4
FBE4
FB55
FB1E
FB97
FC1C
FBF5
FB54
FAFD
FB42
FBAF
FBCE
FBBB
FBB7
FB91
FAFC
FA7B
FB53
FE2E
0204
04D4
058F
04F5
047C
04B2
050C
04FE
04BE
04C3
04FA
04EC
0488
044D
048D
04E4
04BC
0428
03DA
0430
04B0
04B4
0451
042E
047A
04A8
0451
0403
0493
05A5
0587
02FC
FEE6
FB9D
FA8B
FAEC
FB1C
FA9C
FA4D
FADA
FBAE
FBCE
FB42
FAF2
FB52
FBC2
FB94
FB16
FB1A
FBBE
FC38
FBFB
FB79
FB72
FBD4
FBE7
FB6D
FB0D
FB4F
FBAF
FB4E
FA6F
FA98
FCED
00B2
03E3
0538
052B
0504
0545
0571
051C
04A2
0494
04DC
04E3
0480
0442
049F
0530
0528
0469
03BC
03CD
0454
048D
0453
043F
049E
04E8
0492
041C
0488
05B6
05E8
038D
FF45
FB9B
FA72
FB3C
FBEF
FB73
FA86
FA56
FAED
FB66
FB45
FAFD
FB18
FB63
FB59
FB04
FAFA
FB7D
FC09
FC08
FB9C
FB64
FB99
FBCC
FBA6
FB70
FB8E
FBB4
FB3D
FA56
FA59
FC76
002D
0386
04FE
04DB
0480
04B4
0514
050B
04C3
04CF
0536
0565
050E
04A9
04C5
0533
0541
04B7
0434
0452
04CE
04E1
0456
03D1
03E9
0458
0472
0443
048D
057F
05E0
0422
0050
FC6F
FA97
FAEC
FBC4
FBB4
FAF0
FA8F
FAED
FB58
FB30
FAC1
FAAF
FB08
FB47
FB26
FAFA
FB19
FB56
FB5B
FB3E
FB63
FBCA
FBFC
FBC3
FB92
FBD1
FC0C
FB72
FA3B
F9FB
FC23
0034
03F2
0587
0527
0473
0483
0505
052C
04E7
04D1
0523
055F
0511
0488
0471
04E5
0542
050E
0498
047E
04C6
04E2
0493
0448
0470
04BC
048F
0409
040B
04E1
055F
03E0
0047
FC74
FA77
FA93
FB5B
FB8A
FB31
FB17
FB6A
FB96
FB3E
FABE
FAA9
FAFF
FB50
FB65
FB6F
FB8F
FB8B
FB38
FADD
FAE8
FB4E
FB90
FB6C
FB47
FB94
FC08
FBDF
FB0F
FAD6
FC90
0015
0396
0551
0535
04A0
04A4
0503
04EF
0454
03F4
0451
0506
0556
051E
04CF
04B2
048F
043C
0407
0454
04F5
0549
0509
049B
046F
0460
041B
03DE
0458
0572
05C5
03D1
FFD1
FBE4
FA21
FAA0
FBAF
FBD2
FB2D
FAD6
FB42
FBCA
FBB3
FB28
FAE8
FB37
FB93
FB7E
FB30
FB3B
FBB5
FC13
FBE5
FB5E
FB06
FB0A
FB39
FB76
FBD1
FC1D
FBD6
FAED
FA78
FBEB
FF70
0353
0584
0596
04E4
04CD
054B
057E
051C
04B7
04B6
04BA
045D
03FB
0436
04E5
0521
0483
03C6
03CF
0473
04C5
047D
0459
04DE
0564
04F7
03EA
03A4
04AC
0594
045E
00D7
FCFE
FAE4
FAAE
FAEF
FA97
F9FD
FA06
FACE
FB9B
FBD0
FB99
FB83
FBB3
FBD1
FB9A
FB46
FB3F
FB92
FBE4
FBDF
FB8C
FB2E
FAF4
FAF0
FB37
FBC3
FC29
FBD3
FAD2
FA58
FBCE
FF45
0310
054A
0599
0532
0534
058C
0586
0509
04B1
04CC
04E5
0481
03F4
03EF
047C
04E4
04AA
0439
0446
04D6
053D
0510
04AC
0499
04C0
049C
042B
041D
04D2
056A
045B
0120
FD16
FA62
F9EF
FAC6
FB59
FB26
FAD9
FB07
FB68
FB6A
FB1A
FB05
FB5B
FBAC
FB95
FB4F
FB49
FB73
FB5E
FB02
FAE4
FB43
FBA0
FB71
FB0B
FB37
FBF2
FC36
FB66
FA88
FB7B
FECE
02DD
0559
058F
04C8
0492
0523
0594
0547
04A5
046F
04C1
050A
04EC
04B5
04D6
0528
051A
0493
0430
0477
051D
0560
0505
048D
046B
0466
042C
0414
04A2
0550
048C
0180
FD6D
FAA1
FA1D
FAC8
FB0E
FAAE
FA81
FAEE
FB5C
FB41
FAFC
FB29
FB9A
FB9C
FB19
FACB
FB2C
FBB3
FB97
FAF5
FAB0
FB30
FBC8
FBB0
FB2A
FB27
FBD7
FC3A
FB82
FA7F
FB22
FE5E
02D4
05F2
066C
054E
048F
04F0
058D
0562
04A4
044F
04BF
0542
051B
0481
0438
047D
04CF
04CA
04AF
04D7
050A
04D4
0454
0427
0482
04D1
0496
0442
0494
052B
047A
0189
FD6F
FA7A
F9DF
FAB4
FB48
FB03
FA9E
FAD0
FB68
FBC4
FBBE
FBAD
FBB5
FB90
FB1A
FAAE
FAB7
FB17
FB53
FB42
FB42
FB8E
FBC8
FB76
FADC
FAD6
FBA4
FC54
FBE4
FADC
FB2D
FE0E
024D
0553
05C2
04B4
042D
04CD
057D
0537
0458
03F1
044A
04AD
0494
0461
04B1
055D
05AA
0546
04B3
0489
04BA
04CD
04A7
04A5
04E5
04F7
0482
03F2
0408
04AA
048B
026F
FEBB
FB63
FA14
FAAC
FB9B
FBB2
FB2B
FAED
FB47
FBB0
FBA8
FB4D
FB0D
FB09
FB0F
FB0E
FB26
FB4C
FB42
FB02
FAE8
FB2D
FB75
FB44
FAD2
FAED
FBCA
FC76
FBEC
FAAD
FAAB
FD37
0157
049D
0598
0505
048D
04D3
051F
04C5
042F
043F
0504
0591
0532
044F
03E6
0448
04D8
04F3
04BB
04BB
050E
0543
0514
04D5
04E2
050B
04E0
0488
049E
0520
04E1
02AD
FEE4
FB7B
FA1E
FA9B
FB67
FB6A
FAEB
FAC1
FB14
FB63
FB61
FB56
FB93
FBE9
FBF4
FBB0
FB78
FB77
FB71
FB2A
FAD0
FAB9
FAE1
FAFA
FAF4
FB1E
FB89
FBA7
FAF3
FA02
FA61
FD0B
011A
046C
0598
0512
045E
0465
04E5
053E
0542
051B
04D2
0450
03CA
03B5
0435
04D8
050F
04D0
048E
049D
04D3
04E7
04E7
051E
057E
058B
0504
0472
049B
055E
0569
0370
FFBD
FC33
FA89
FAB3
FB48
FB49
FAFE
FB13
FB77
FB95
FB4F
FB31
FB8E
FBF5
FBD2
FB4C
FB09
FB38
FB5E
FB23
FAD1
FACA
FAE9
FAD9
FAAB
FAAC
FAD7
FAE6
FAD8
FAF6
FB3B
FB38
FB00
FBAD
FE49
0228
0528
05F1
0544
04BD
04D6
04DB
046A
040A
043E
04BA
04F3
04F2
0517
0540
04F2
044F
0423
04C1
0574
058C
054F
0559
058A
054E
04C1
049C
0509
0540
04C6
0453
04B0
0503
0376
FFBE
FBF9
FA62
FAD7
FB81
FB5A
FB04
FB39
FB98
FB64
FAC4
FA8C
FAFD
FB7B
FB8A
FB5B
FB35
FAFB
FAAB
FAB9
FB54
FBCF
FB75
FAA5
FA63
FAE2
FB42
FAF8
FAAD
FB28
FBD8
FB8B
FA91
FB02
FE36
02BF
05C7
061D
050B
0463
0493
04F6
0528
054F
056D
0531
04AA
046A
04B8
0514
04F1
0490
0494
04F8
051D
04CA
048A
04D3
0550
0563
0515
04EC
0506
04F3
04A1
04B0
054A
0545
032C
FF41
FBA3
FA27
FA85
FB0A
FAC4
FA4A
FA70
FB05
FB4C
FB1C
FAFA
FB30
FB74
FB7B
FB6A
FB7A
FB8F
FB77
FB4B
FB40
FB27
FAB3
FA2D
FA4C
FB22
FBCA
FB8F
FAF5
FAF0
FB6A
FB6C
FAEE
FB86
FE8E
02F9
060B
064E
0506
0451
04B7
0536
0524
04F7
052D
056C
0526
0488
0437
0456
0474
045B
0467
04CD
052B
0528
0502
050C
0515
04CE
0475
048A
04DF
04C5
043A
042D
0507
056A
036C
FF2D
FB3E
F9F4
FAF8
FC1C
FC0C
FB50
FAEA
FAEF
FADE
FAAC
FAC0
FB2F
FB8B
FB8C
FB63
FB45
FB1C
FAE6
FAFD
FB87
FC02
FBD9
FB48
FB12
FB6F
FBC0
FB91
FB44
FB5D
FB82
FAFA
FA31
FADD
FE01
0254
0547
05A1
048A
03EC
0465
0520
054B
0502
04D6
04F4
051B
051B
050C
0507
0502
04F2
04D3
049B
044B
0414
0435
0498
04D3
04B1
0489
04C3
0523
050A
0482
046C
0530
05A8
0411
003A
FC2C
FA35
FA91
FB84
FB92
FAF2
FAB2
FB15
FB78
FB6B
FB33
FB31
FB49
FB35
FB05
FB05
FB3F
FB75
FB86
FB8B
FB79
FB24
FAB2
FA97
FAEE
FB31
FB06
FAD9
FB32
FBB9
FB97
FAFC
FB80
FE4C
024B
0505
0553
0474
042F
04BB
0515
04D2
0490
04C5
0509
04D6
0470
046D
04CD
0503
04E7
04DC
0509
0507
04B6
04AA
0546
05EC
05C7
0509
04A6
04DE
04F1
0474
0435
04E5
056A
03B2
FF7B
FB44
F9BB
FADB
FC56
FC70
FB8C
FAE5
FAD8
FADF
FAB9
FABB
FB13
FB68
FB62
FB22
FAEE
FACB
FAB8
FAE8
FB5C
FB96
FB34
FA9B
FA83
FAEF
FB22
FACE
FA9A
FB20
FBC8
FB8C
FACC
FB67
FE74
0297
054E
05AB
04F6
04BF
0526
055B
051C
04EA
0509
0513
04BF
047B
04C2
0555
058B
0545
04F9
04EC
04E6
04C3
04C8
0526
0573
0530
049D
047B
04F1
0542
04EE
0481
04A5
04B8
0330
FFAB
FBE2
FA04
FA5D
FB41
FB36
FA7D
FA3C
FAC1
FB4F
FB49
FAF6
FADD
FB02
FB0D
FAED
FAE3
FB0A
FB2F
FB2D
FB22
FB23
FB16
FAF9
FB03
FB41
FB60
FB2C
FB00
FB45
FBA7
FB73
FAE0
FB76
FE59
0289
0590
061B
053F
04C9
051F
0562
0526
0504
056E
05D0
056F
0494
043D
04B6
054A
0559
051A
04F4
04CF
0481
0462
04CB
0558
0549
04A4
043A
0474
04C1
0498
046B
04CE
04F8
033E
FF73
FBBA
FA4A
FAED
FB9A
FB24
FA52
FA3E
FABC
FAE4
FA97
FA90
FB0F
FB5F
FAF0
FA44
FA32
FAC5
FB61
FBAB
FBC0
FBB5
FB81
FB54
FB7E
FBD1
FBB4
FB12
FAC3
FB72
FC61
FC32
FB0A
FAFA
FDA2
01F1
0529
05DA
0515
04A6
04F8
0537
04F2
04B0
04FA
0583
05AD
056E
0532
0523
0510
04E8
04D8
04E8
04DF
04AA
0490
04C3
04F9
04D4
0476
044F
046A
0456
0405
041A
04DC
0539
0397
FFDD
FC07
FA3E
FAAA
FB99
FBAD
FB2C
FB0A
FB5C
FB61
FAD0
FA4C
FA76
FB0F
FB5E
FB26
FAD6
FACF
FAF5
FB05
FAFA
FAF1
FAF5
FB11
FB56
FB91
FB6A
FAF4
FAE1
FB99
FC5D
FC0C
FAEE
FB0A
FDED
026B
0588
05C2
048F
0436
050F
05B1
053B
045C
040C
044B
0491
04D8
0564
05DD
0590
04A5
042E
04B7
0575
057D
050B
04EA
051C
0504
049B
0492
050E
0537
0486
03D8
0436
04CE
0388
FFDD
FBFD
FA53
FABE
FB41
FAD6
FA5D
FAC3
FB8C
FBB3
FB37
FAF8
FB41
FB6F
FB17
FAB2
FAC3
FB0F
FB23
FB16
FB25
FB19
FAB9
FA7B
FAF2
FBBD
FBD6
FB1A
FAB5
FB72
FC4D
FBC7
FA6C
FAC6
FE37
02E3
05A3
058C
0474
0453
0528
05BF
058E
0516
04DB
04CC
04BC
04D6
052E
0565
052E
04C8
04A6
04BE
04B8
0497
04B6
0519
0549
050B
04C2
04CF
04E6
0480
03EB
0423
054B
05D2
03E5
FFAF
FB8C
F9B7
FA32
FB39
FB6A
FAF5
FABE
FB02
FB46
FB38
FB0C
FB07
FB0A
FAE4
FAB8
FACE
FB1B
FB49
FB2D
FAF4
FAD7
FAE2
FB1F
FB91
FBEE
FBB9
FAFC
FA8F
FB1A
FBFD
FBEA
FADD
FACD
FD8F
0249
05F1
0697
0557
0498
0521
05C0
056E
04A3
045C
04B0
04F7
04EC
04ED
0527
053F
0501
04C9
04E4
0511
0507
04F8
051F
052E
04CE
0459
0476
04F7
04F8
0447
03F7
04C9
057F
03EC
FFD1
FBA5
F9DD
FA4E
FAF0
FAA8
FA2F
FA70
FB20
FB68
FB2F
FB01
FB13
FB05
FAB5
FA90
FAD2
FB11
FAF3
FACE
FB13
FB7C
FB74
FB0C
FAE0
FB19
FB33
FAF5
FAF6
FBAF
FC69
FBFE
FABA
FAA9
FD60
01EF
05A6
06C9
05FC
050C
04F6
0566
05A4
0577
0520
04DF
04C7
04D3
04F1
0509
0513
0522
0540
0550
053E
052F
054C
0565
051B
0476
0409
0441
04B8
04AF
042B
0415
04E4
0578
0405
003D
FC13
F9DE
FA04
FAE9
FB0B
FA87
FA52
FAB3
FB0B
FAF0
FABC
FAEB
FB5D
FB9D
FB8A
FB5C
FB24
FABF
FA49
FA24
FA66
FAAB
FAB8
FADE
FB62
FBDE
FBC9
FB51
FB2A
FB77
FB92
FB46
FBAA
FDFF
01CB
04EE
05E8
0555
04D3
0500
0549
0537
0510
0526
0543
0516
04CE
04CC
0506
051A
04FF
050D
054E
0553
04FB
04C9
0519
0572
0533
0499
046C
04D0
0512
04C8
0479
04B0
04C3
0355
0023
FCA5
FA96
FA42
FAB9
FB19
FB31
FB16
FAD2
FA8C
FA86
FAC3
FAF7
FAF4
FAEB
FB0F
FB2B
FAEA
FA80
FA83
FB18
FBA1
FB99
FB42
FB2C
FB52
FB40
FAF5
FAFD
FB8B
FBF6
FB9C
FAFB
FB76
FDCB
011D
03CD
0506
053C
0547
057F
05A6
0579
0514
04DC
050C
0577
05A8
0564
04EB
04B2
04E4
053A
055A
053A
0512
04F1
04AD
043A
03E3
03F9
0475
04FD
053F
0525
04C8
0465
0451
04B2
051E
04AC
02BB
FFAC
FCBE
FAFE
FA78
FA82
FA91
FA9B
FAC2
FAEE
FAEE
FAC6
FAB0
FAC4
FADE
FADB
FAD2
FAEB
FB1A
FB2A
FB15
FB16
FB5A
FBAF
FBB7
FB69
FB27
FB4A
FBA0
FBA0
FB1E
FA96
FA98
FB0B
FB3D
FAE6
FADC
FC67
FFC7
038B
05C2
05CE
04D6
0467
04E0
056D
0553
04DC
04C3
0526
0568
051F
049B
046C
04A4
04EA
050A
051E
0532
0516
04B9
046E
048C
04E5
04F7
04A8
0477
04BF
0522
04FF
046C
0438
04D2
0570
049F
01C7
FDEC
FAE7
F9DA
FA60
FB38
FB76
FB28
FAE5
FAFF
FB3A
FB3B
FB02
FAD8
FADD
FAEC
FAEE
FB04
FB36
FB3D
FAE5
FA79
FA85
FB18
FB92
FB74
FB0A
FB06
FB75
FBAF
FB56
FAF1
FB1E
FB88
FB51
FA96
FAD8
FD62
0182
04E3
05D6
04E6
03EF
040F
04D3
0545
052C
0501
0513
052C
0512
04ED
04F9
051D
0510
04DA
04D8
0529
0562
051C
0494
0473
04E8
0562
054A
04CF
0495
04BF
04C2
043D
03B3
03FE
050C
0585
0405
0098
FCE4
FAB8
FA92
FB6D
FBE7
FB85
FAD8
FA9C
FADE
FB19
FB06
FAE7
FB06
FB36
FB16
FAB0
FA77
FAA7
FAE7
FAD5
FAA4
FACF
FB4F
FB98
FB6E
FB46
FB82
FBC8
FB8B
FB01
FAF2
FB7E
FBB8
FAF7
FA25
FB12
FE56
025F
04F7
0567
04CC
0483
04DC
0541
0532
04CB
0485
04A5
0506
054C
0544
0506
04D5
04D4
04F0
0507
050F
050C
04EC
049A
0442
042F
0467
04A2
04B8
04DD
0526
053E
04DC
0473
04C2
0593
0563
02DE
FEA6
FB19
FA02
FAE1
FBCB
FB9E
FAE0
FA93
FAD5
FAFC
FAB2
FA6A
FAB1
FB64
FBE1
FBD1
FB81
FB56
FB44
FB0F
FAD5
FAFB
FB8A
FBF9
FBCD
FB3F
FAF8
FB27
FB41
FADA
FA66
FA9A
FB46
FB6D
FACD
FAAE
FC92
004D
03EB
05A2
0578
04D4
04CA
053F
0586
0558
04FB
04BF
04B4
04C3
04C8
04AE
0481
046C
047C
0490
0494
04A1
04C4
04D2
04AA
0478
0484
04D0
0510
0528
054B
0580
0560
04BB
0445
04CC
05A4
04D4
0162
FCEC
FA24
F9F8
FAE8
FB2B
FAA8
FA6C
FAD8
FB35
FAFB
FA9A
FAAF
FB0A
FB27
FB10
FB36
FBA0
FBD7
FB9F
FB46
FB24
FB30
FB30
FB22
FB2E
FB55
FB64
FB3C
FAFE
FAD9
FADC
FAFD
FB13
FAE6
FAA1
FB34
FD98
0166
04B0
05DB
0550
04CB
0532
05CD
05AC
0516
0503
058D
05C7
052D
046F
0466
04DF
050F
04C8
048B
049F
04BB
04A1
048D
04C4
050A
04F1
0482
0446
048E
0501
0517
04D5
04C1
052A
05A1
0528
02F8
FF60
FBE2
FA1C
FA47
FB14
FB37
FAB8
FA88
FAFF
FB6C
FB24
FA76
FA33
FA8B
FAF1
FB09
FB1F
FB70
FBA0
FB4C
FAC6
FAB4
FB22
FB7A
FB6C
FB51
FB87
FBCD
FB96
FAEC
FA86
FAE0
FB83
FB94
FB07
FAF8
FC9D
FFF1
0378
056E
055F
0479
0441
04F8
0596
0550
0498
0468
04EE
0573
056D
0522
0518
0548
0543
04F4
04BB
04C8
04CC
0491
0464
0498
04F2
04F6
04AC
0498
04E8
051F
04C5
042C
042C
04FC
059B
0491
016F
FD73
FA98
F9EE
FAD1
FBAE
FB90
FADF
FA95
FAE6
FB29
FAED
FA9E
FAC7
FB3F
FB70
FB38
FB07
FB1F
FB39
FB13
FAF6
FB40
FBA4
FB7A
FAD1
FA8A
FB22
FBE3
FBD7
FB25
FAD0
FB45
FBB9
FB5B
FAA3
FB13
FD87
0126
0414
0524
04BF
043B
0487
0569
05F6
05A4
04E5
048A
04C8
051A
0512
04E3
04E3
04F2
04C3
0480
049F
0523
0574
0530
04C1
04C6
051C
050F
0478
0415
0466
04DE
04B3
042F
0459
0550
05A1
03C5
FFFF
FC54
FA9C
FAD7
FB96
FB9D
FAF2
FA5B
FA5C
FAC8
FB26
FB39
FB2A
FB2F
FB43
FB3B
FB19
FB06
FB05
FAEE
FACB
FAE0
FB3D
FB78
FB2B
FAA2
FA97
FB34
FBB2
FB5C
FAA3
FA9A
FB65
FBD9
FB2E
FA6C
FB7F
FEE5
02E5
054B
0586
04D9
04A3
050D
0554
0505
0479
0448
0492
04FE
0528
0508
04DE
04DB
04E4
04D1
04B6
04CD
0507
0511
04D2
04A4
04CE
0516
0510
04D2
04DE
054B
0579
04FB
0475
04D6
05A6
0502
01CD
FD62
FA6A
FA1C
FB3A
FBDD
FB7F
FB00
FB10
FB58
FB45
FAEA
FAC3
FAF0
FB24
FB35
FB47
FB67
FB62
FB17
FACA
FAD7
FB45
FBAC
FBB0
FB65
FB36
FB59
FB7F
FB38
FA90
FA25
FA6D
FB06
FB16
FA87
FAA9
FCEE
010B
04C7
061C
0538
040F
0418
04FD
0586
0540
04C8
04B5
04E7
04F7
04E2
04E5
04F6
04D0
047B
044B
0464
047C
044B
0408
0425
04A5
050B
04F8
04B9
04DC
055C
058D
04FF
0444
045F
056A
0601
0474
00A4
FC76
FA29
FA46
FB53
FB97
FAD3
FA18
FA46
FB11
FB98
FB80
FB34
FB2F
FB65
FB7B
FB5E
FB52
FB84
FBCE
FBF0
FBDC
FBAC
FB6E
FB25
FAF4
FB14
FB82
FBDA
FBBF
FB5F
FB4A
FB9C
FBA1
FAC0
F9B5
FA54
FDA4
025E
05D8
0688
0560
0474
04AE
0542
0530
0499
044F
048D
04CD
04B7
049D
04DD
0533
0511
0479
040B
042E
048F
04A5
0472
045C
0473
0459
03E9
03A7
041B
04FA
055A
04DC
0446
048B
0558
0508
026C
FE5D
FB28
FA55
FB43
FC1E
FBDE
FB0C
FAA6
FADC
FB1A
FB09
FAF7
FB31
FB7E
FB7F
FB48
FB3E
FB74
FB8D
FB51
FB10
FB27
FB76
FB8C
FB5A
FB53
FBB3
FC0F
FBDC
FB4F
FB2F
FBC5
FC4D
FBDD
FABE
FA7E
FC77
004B
040D
05F1
05C1
04BA
042F
0473
04F9
0531
051B
0506
0517
0522
04F8
04A9
0468
0452
0460
0484
04B3
04D6
04D7
04BD
04AB
04B4
04B9
0494
0461
0464
04A9
04D1
0484
0406
0408
04C0
053B
0410
00E0
FD04
FA78
FA16
FAF4
FB90
FB59
FAE6
FADE
FB25
FB2E
FADB
FAA4
FAE2
FB50
FB71
FB37
FB0B
FB37
FB86
FB9E
FB71
FB41
FB38
FB42
FB49
FB52
FB5E
FB47
FB07
FAED
FB4C
FBEA
FC04
FB3C
FA6B
FB1E
FDFF
01E8
04CE
059D
0512
04A2
04EC
0560
0558
04F5
04CE
0508
0534
0508
04CA
04D3
04F8
04CD
0459
042F
049C
0525
051B
0483
041B
045D
04E8
050F
04C2
0489
04B5
04FA
04FB
04E3
0511
0547
049D
0273
FF4D
FC7A
FAE8
FA7F
FA8F
FA9D
FA9E
FAA9
FAB8
FAC3
FADD
FB16
FB4D
FB4F
FB2C
FB2A
FB6C
FBB9
FBBD
FB7E
FB4C
FB52
FB57
FB1B
FAD3
FB00
FBB1
FC3F
FBF7
FB15
FA9A
FB1A
FBDD
FBAB
FA78
F9DD
FB8F
FF6D
036C
058E
05A3
050C
04F5
0552
057A
053F
050F
0527
053E
0507
04B3
049E
04C4
04CD
0499
046D
0481
04A9
04A8
049E
04CC
0515
0509
0498
0448
047F
04DF
04BE
0424
03E0
0470
0542
0573
04FE
04AF
04D7
048F
02BA
FF87
FC78
FAD4
FA83
FA8A
FA59
FA38
FA84
FB09
FB4B
FB3C
FB3C
FB7D
FBAB
FB61
FAC9
FA75
FAB6
FB41
FB96
FB95
FB7E
FB7E
FB6E
FB1A
FAA9
FA7D
FAC4
FB45
FBA2
FBAD
FB76
FB29
FAFE
FB22
FB79
FB8F
FB1A
FAA9
FB7C
FE49
0220
0502
05BF
050F
048E
04EC
056E
0537
047E
0429
048A
0507
0509
04C2
04BC
04FE
050C
04AD
0448
0455
04C3
0522
053F
053A
052D
0502
04B8
048C
049D
04AE
0483
044F
0477
04E1
04FB
048E
043A
0497
050C
0414
00FD
FD05
FA50
F9D4
FAA9
FB5A
FB6D
FB60
FB91
FBB5
FB68
FAD8
FA8A
FAB2
FB0A
FB4B
FB73
FB92
FB95
FB69
FB2A
FB03
FAF3
FAD8
FABD
FADA
FB3C
FB98
FBA5
FB7B
FB6B
FB85
FB88
FB61
FB62
FBC1
FC14
FBB2
FACA
FAAC
FC98
0041
03CB
057D
0544
0479
0444
049B
04CA
048F
0461
04A8
0521
053C
04DA
046E
0460
049D
04CB
04C7
04B3
04B0
04B8
04BC
04C4
04CE
04C2
049A
0484
049C
04AD
046D
03FD
03DE
043D
0497
0466
0402
0448
0537
055E
0344
FF50
FBB4
FA45
FABA
FB68
FB4B
FADC
FAE9
FB58
FB78
FB25
FAEC
FB22
FB62
FB3A
FAF0
FB12
FB93
FBCC
FB69
FAEB
FAEF
FB53
FB7F
FB4F
FB3D
FB99
FBFF
FBF5
FBA3
FB92
FBD5
FBEE
FBA5
FB6A
FB90
FB9A
FAE7
FA06
FAA2
FDAC
01EB
04FA
05AE
050F
04D0
055B
05C4
055A
049A
046D
04E5
0542
0505
0482
0455
0495
04DE
04E8
04C7
04A7
0492
0489
04A0
04D9
04F5
04BC
045A
0437
046A
0499
0475
043B
0454
04AF
04CC
048E
0492
053A
05AE
0453
00AE
FC5C
F9C1
F9B6
FAE9
FB8A
FB2B
FAAD
FABE
FB10
FB0E
FAD3
FAEE
FB74
FBCB
FB83
FAF4
FAC1
FB01
FB3E
FB28
FAF4
FB00
FB52
FBA6
FBC4
FBA4
FB4B
FADA
FAA4
FAEE
FB77
FB9F
FB2D
FABA
FAE8
FB75
FB80
FAED
FAFF
FD11
00CA
0436
05B0
0573
04EA
04F0
0535
0528
04E9
04EB
052F
053E
04F3
04B8
04EC
054E
055A
04FE
04A7
04A4
04CE
04D4
04AA
0485
048B
04BE
050E
0558
055A
04F0
0469
0457
04D6
053F
04E7
041D
03F4
04DA
05BC
04E7
01DF
FDFB
FB2D
FA48
FAA1
FB15
FB19
FAD9
FAA7
FAA2
FAB4
FAC4
FAC5
FAC6
FAE7
FB3B
FB9E
FBC5
FB90
FB2D
FAEB
FADD
FAE4
FAEF
FB19
FB63
FB86
FB46
FAD5
FABC
FB34
FBC4
FBC1
FB27
FAAF
FAF3
FB9C
FBBD
FB0E
FA8C
FBA3
FEAC
026B
0516
05DD
055B
04BB
04A5
04F7
054D
0576
0573
054D
050D
04D3
04C3
04D8
04E4
04CC
04AB
04AB
04CA
04DF
04D0
04A9
0486
0474
047E
04A7
04D7
04DF
04B2
0490
04C1
051C
0519
0488
0405
045D
055E
059B
03BA
0000
FC4B
FA62
FA69
FB19
FB49
FAF7
FACA
FB04
FB3E
FB17
FAC2
FAB3
FAFC
FB38
FB1E
FAE7
FAFF
FB66
FBAC
FB7F
FB20
FB16
FB82
FBEB
FBC3
FB11
FA6F
FA6F
FB07
FBA8
FBC8
FB60
FAED
FAF3
FB74
FBD8
FB88
FAC7
FAD3
FCDC
009E
0440
05E2
0562
0457
0448
052B
05D3
0592
04F1
04C2
0504
0517
04C5
048F
04D0
0526
04FF
0478
0438
047E
04C5
0488
0408
03F4
047C
0512
052E
04E8
04AC
04A3
04A5
049A
0490
0483
046B
047B
04EB
054B
046C
0194
FDB7
FAEC
FA66
FB3F
FBA8
FAFB
FA27
FA24
FAB4
FAFD
FAD5
FAD9
FB52
FBAD
FB66
FAE4
FAF4
FB9B
FC02
FBA4
FB06
FAFB
FB8B
FBF7
FBC5
FB43
FAFC
FB04
FB21
FB49
FB97
FBE1
FBD8
FB90
FB81
FBBE
FBA4
FAC6
FA15
FB4A
FEEF
0349
05D9
05D7
04C3
0478
0539
05E4
05AA
04F7
0497
04A8
04B8
049F
04AE
04FF
052E
04E1
0462
0444
049A
04E1
04BE
0474
0476
04BC
04E7
04D6
04CB
04DA
04B9
043D
03D2
03F9
0488
04C8
0487
046D
04EE
052D
03A3
0017
FC53
FA79
FAD0
FBB5
FBA6
FAD4
FA6B
FADD
FB76
FB83
FB3A
FB33
FB77
FB86
FB28
FABF
FAAE
FAD8
FAF1
FAFE
FB3E
FBA6
FBE5
FBD4
FBA9
FB90
FB65
FB15
FAF1
FB4C
FBCF
FBC1
FB12
FAA2
FB19
FBD1
FB9A
FA93
FA93
FD27
017E
04F9
05DA
04E0
040B
0448
04E4
04F5
049C
048F
04F8
054B
0528
04D1
04B5
04D4
04E6
04D8
04D0
04CF
04A8
0460
0440
0470
04AA
04A1
047B
0495
04E4
04E9
0473
0415
046B
0529
0559
04B8
0441
04E1
05E1
0545
0207
FD94
FA8E
FA2F
FB47
FBDD
FB54
FA9E
FAAB
FB49
FBA2
FB62
FAF1
FABB
FAB7
FAB9
FAD2
FB26
FB82
FB7F
FB03
FA72
FA37
FA64
FACA
FB44
FBAE
FBCC
FB7D
FB16
FB24
FBB1
FC14
FBC4
FB2C
FB29
FBB2
FBB8
FAAB
F9D4
FB3C
FF37
038D
05A1
051F
0404
0419
0519
0598
0519
0483
04AE
0544
0564
04E5
047D
04B4
0551
05C5
05D9
05A4
053A
04B8
046E
0499
04FE
0517
04CD
049E
04DA
0516
04C8
0438
0441
04F9
055A
04A4
03AC
03F3
0566
05E3
0392
FF40
FBB9
FABD
FB68
FBB6
FB09
FA62
FA98
FB2E
FB40
FADB
FAC0
FB2D
FB81
FB3C
FAB8
FA92
FAC6
FADC
FAB6
FABB
FB19
FB70
FB6B
FB57
FBA7
FC23
FC1A
FB6D
FAD5
FAE5
FB35
FB11
FAAF
FAEE
FBDA
FC33
FB11
F99C
FA36
FDB9
023E
0516
058A
0519
0536
05AD
0580
04A7
0421
0484
0540
0587
055C
054D
0578
0576
0525
04ED
0509
0519
04B6
0431
0434
04B2
04DF
045F
03E0
0430
04FF
0543
04B5
0434
0475
04F0
04C2
0434
047B
05C8
0668
048E
009D
FCE4
FB20
FAE9
FAD8
FA7A
FA71
FB00
FB68
FB03
FA46
FA1D
FAA1
FB0F
FAF4
FAB5
FAC5
FAEC
FAC4
FA88
FACA
FB74
FBBC
FB54
FB00
FB83
FC66
FC76
FB73
FA7F
FA96
FB42
FB65
FAF0
FAEE
FBC2
FC4D
FB6F
F9F1
F9FB
FC9C
0081
037D
04C2
0524
0580
05C0
058C
052E
0533
0586
058C
0514
04A6
04B1
04F0
04E8
04BA
04DD
053F
0536
0486
03E9
0425
04E2
0511
0465
03CE
042F
0523
057E
04EA
0443
0451
04B3
0495
040E
0415
0505
05C6
04E4
0234
FF01
FC9B
FB43
FA7D
FA14
FA3B
FAE6
FB81
FB7D
FAEB
FA58
FA37
FA88
FB07
FB6B
FB7C
FB3A
FAF5
FB18
FBA1
FC01
FBB2
FAF5
FA9B
FB0C
FBC2
FBF8
FB9E
FB57
FB7C
FBA2
FB56
FAED
FB2E
FC1C
FCA6
FBEA
FA85
FA37
FC17
FF6A
026F
041A
04BE
052F
05AB
05CC
055F
04C5
0490
04D6
052E
0534
04ED
04B1
04BC
04F3
050A
04D9
0490
0488
04E5
0550
0547
04A4
03DC
039C
0418
04DA
053C
0508
048B
0430
0421
0445
046D
0470
0437
03E2
03DC
0488
05A7
063F
0546
02A8
FF78
FD07
FBC8
FB2E
FA8F
F9FC
FA06
FAD7
FBBD
FBD0
FAF1
F9FE
F9EC
FACE
FBCF
FC17
FB92
FADB
FA89
FAB3
FB0F
FB58
FB74
FB74
FB75
FB90
FBBF
FBD0
FB9A
FB49
FB4C
FBD2
FC60
FC3C
FB4B
FA62
FA79
FB88
FC78
FC38
FAE5
F9BC
F9F4
FBC0
FE56
00B5
025F
037A
046A
0551
05E8
05D1
051F
0473
0469
04EF
0551
050F
0476
0438
0484
04DD
04D2
049B
04A8
04EA
04E0
0465
0407
044A
04E0
0507
048F
041E
0434
0476
0440
03BB
03C3
04A6
0581
0548
0434
03A1
046B
05DD
0677
0585
038D
0163
FF4F
FD34
FB41
FA00
F9D0
FA82
FB81
FC2D
FC25
FB79
FAC0
FAAF
FB60
FC14
FBFF
FB3C
FAAA
FAD2
FB3B
FB27
FAAF
FAAD
FB78
FC4C
FC3E
FB6A
FACC
FAF3
FB6F
FB9E
FB93
FBB5
FBE2
FB81
FAA0
FA42
FB2C
FCA2
FD07
FBC3
FA13
F9AE
FAF3
FCDA
FE74
FFED
01E0
0425
05C7
0613
054D
0457
03E5
0425
04DC
0590
05C5
0551
04A2
0460
04BA
0535
054A
0502
04C1
04AA
0486
0445
043A
049B
050E
0509
0498
044A
0465
047D
0436
03F3
045A
0532
055B
044B
030D
033E
050E
06D7
06D6
04FE
02A9
00D4
FF43
FD5F
FB5F
FA21
FA0F
FAAE
FB3F
FB74
FB67
FB25
FAB3
FA51
FA5E
FAE6
FB78
FB9B
FB43
FAC5
FA79
FA8D
FB07
FBB7
FC24
FBE5
FB2F
FABC
FB01
FB91
FBAF
FB4C
FB15
FB69
FBB8
FB53
FA96
FA9E
FBB7
FCA8
FC13
FA3F
F8FB
F9A1
FBB8
FDD6
FF67
0108
033E
056A
0671
060D
0514
047F
048C
04E6
053C
0577
0581
0539
04AE
0434
0420
0480
051B
059A
05A5
0515
043E
03D4
044B
0539
05AF
0542
0486
044F
04A7
04E9
04C6
04BA
052E
059D
0523
03E6
0339
0418
05C5
0681
057C
039D
0221
010E
FF65
FCC7
FA41
F93C
F9F7
FB55
FC0C
FBBE
FAF0
FA51
FA32
FA7F
FAF0
FB39
FB41
FB22
FB04
FAE8
FACA
FAD0
FB2C
FBBC
FBFC
FBA0
FB01
FAC8
FB15
FB53
FB13
FAAF
FAC8
FB4E
FB7C
FAF4
FA62
FA9D
FB6A
FB9F
FAB0
F98B
F99D
FB21
FD00
FE51
FF72
0150
03E7
05F9
0660
0557
042D
03F2
04A2
0576
05C7
0581
04FC
049C
0488
04A0
04B3
04C0
04F1
054E
0585
0542
04AA
0456
04A4
0543
059B
057E
053F
0512
04C7
0447
040C
0494
0582
05BA
04BF
0387
0380
04D2
0619
05F6
0485
02E6
01A5
0024
FDCB
FB35
F9C4
FA18
FB5D
FC37
FC0C
FB4B
FAAD
FA7C
FA8F
FAAE
FACA
FAEF
FB1F
FB41
FB29
FACC
FA6E
FA78
FAFC
FB86
FB8D
FB16
FAB0
FAB8
FAF3
FAF6
FAD2
FAEE
FB4A
FB55
FAC9
FA47
FAA8
FBBF
FC4C
FB82
FA26
F9C6
FAE7
FC80
FD72
FE0C
FF96
027A
0571
06C2
060F
0496
03D0
0421
04EF
0587
05B3
0590
0537
04C1
0468
0475
04F9
05A9
0601
05A6
04C3
0401
040D
04E6
05BF
05C4
0501
0452
0460
04E9
0544
054D
057C
05EF
0605
0537
041B
03E5
04D9
05C9
057C
0436
033E
02FC
023D
FFC3
FC28
F986
F94C
FACC
FC22
FC35
FB69
FAB2
FA81
FAA2
FACD
FAEA
FAF9
FAF3
FADD
FACC
FACF
FAE2
FB01
FB27
FB32
FB00
FAB1
FAA4
FB02
FB67
FB4E
FACE
FA92
FAF6
FB73
FB4A
FA9E
FA5F
FB09
FBD9
FBBB
FAC1
FA13
FA70
FB41
FBA9
FC0A
FDCA
015C
0530
0713
0675
04E1
042A
04A2
0555
0583
0557
0541
0538
04F3
048E
047F
04EE
057B
05B1
0582
0529
04D0
047D
0448
0454
0496
04CF
04D4
04B9
0497
046F
045E
04AD
0561
05E6
058B
0482
03E6
0480
05B0
061E
0561
0468
03FA
0366
015A
FDD9
FAAF
F98B
FA38
FB18
FB2B
FAEA
FB1E
FB8B
FB5B
FA7C
F9E2
FA4B
FB41
FBB0
FB33
FA73
FA44
FAC1
FB6A
FBD1
FBE7
FBC0
FB66
FAF9
FABF
FAED
FB6B
FBE6
FC10
FBD0
FB50
FAEB
FAF8
FB6A
FBBA
FB62
FA8F
FA18
FA8A
FB6B
FBD3
FBCD
FC9A
FF44
0311
05E6
066B
0550
0459
045F
04D2
04F5
04F4
055B
05F6
05EC
04FF
041A
043F
0539
05D7
0566
047B
0423
04A2
054C
056F
050C
049A
0466
0462
0470
048F
04C1
04EE
04F6
04CB
047F
044B
046C
04E6
055B
055A
04F0
04AC
04D4
04AD
0303
FFA1
FBFD
F9FB
FA1F
FB2D
FBA8
FB4D
FAE6
FAFF
FB41
FB2E
FAE9
FAF4
FB50
FB64
FAD9
FA34
FA40
FB04
FBB1
FB96
FAF6
FAAB
FB14
FBAE
FBBA
FB28
FA9F
FAB2
FB43
FBB9
FBAF
FB53
FB12
FB18
FB30
FB1C
FAF2
FAF7
FB2F
FB3F
FAE8
FAA5
FB8B
FE3B
01FD
0508
0606
053C
042D
0409
04B2
0540
0533
04DB
04B7
04CE
04D1
04B3
04B6
04EC
0506
04BF
0454
044B
04BB
0526
050E
0497
045F
04BF
0556
057C
0507
0479
0471
04EB
0546
04FB
0445
03EA
045A
0521
056C
050C
04AE
04E7
0530
0434
0151
FD91
FADF
FA41
FB02
FBA3
FB68
FAC9
FA8E
FAE3
FB50
FB6E
FB49
FB26
FB21
FB2B
FB3D
FB66
FBA1
FBC5
FBB2
FB81
FB6F
FB8E
FBA7
FB75
FAFA
FA90
FA96
FB0B
FB84
FB95
FB45
FB03
FB22
FB6F
FB74
FB1D
FAEA
FB4D
FBF1
FBF5
FB1A
FA7E
FBBF
FF35
0349
05C6
05E6
04D3
043B
049F
0535
052C
04A6
045E
04A9
0523
0547
050C
04CD
04C9
04EC
0503
04FF
04EE
04D2
04A0
045C
042B
042F
0463
04A1
04BE
04B2
049E
04AA
04D4
04EF
04D4
049D
0482
048F
048A
0451
042F
048E
052F
04F7
02D9
FF20
FB89
F9D7
FA3F
FB61
FBC9
FB46
FAB5
FABD
FB18
FB1D
FAB3
FA67
FAA6
FB31
FB6F
FB2E
FAD1
FACE
FB2A
FB83
FB8D
FB5E
FB3B
FB45
FB63
FB71
FB73
FB85
FBA3
FBA4
FB6B
FB20
FB0E
FB51
FBAD
FBCC
FBA7
FB82
FB81
FB65
FAF0
FA88
FB2C
FD84
0104
0425
05AD
05AB
052D
0513
055C
057A
0534
04E2
04F2
0552
058D
055D
04FF
04E5
0525
0564
054D
04F6
04C2
04DE
0507
04E6
0488
045B
049F
0511
0533
04DF
046B
0441
0469
049E
04B0
04AC
04A5
0480
042C
03F6
0457
0547
05D6
04CA
01D1
FE0A
FB38
FA49
FAB0
FB28
FAFE
FA87
FA6E
FACE
FB29
FB16
FABB
FA8D
FAB5
FAF2
FAF9
FAD7
FAD6
FB0E
FB45
FB34
FAE6
FAB3
FAE0
FB4E
FB96
FB7B
FB2D
FB0F
FB3B
FB6B
FB5D
FB31
FB3D
FB92
FBDB
FBC9
FB7F
FB60
FB84
FBA3
FB8A
FB77
FBB0
FBFB
FBC7
FB06
FAA7
FBD5
FEC4
0248
04C7
058B
052A
04BA
04CD
052D
0560
054C
053E
0572
05B5
05A2
052D
04C9
04E3
055A
0595
0537
048E
043F
0488
0503
0526
04DA
047E
0465
0482
0497
048F
048C
04A6
04C1
04B6
0492
048B
04BA
04EE
04E8
04AC
047A
0475
0478
0466
0475
04F2
0597
055F
0365
FFFC
FCAF
FAF3
FAE4
FB60
FB56
FAB9
FA3E
FA66
FAE8
FB1F
FAC7
FA44
FA35
FACE
FB99
FBE8
FB7A
FAC8
FA84
FAE4
FB72
FBA1
FB6B
FB36
FB43
FB6C
FB79
FB72
FB83
FBA3
FB96
FB4D
FB11
FB28
FB76
FBA2
FB89
FB5C
FB49
FB41
FB26
FB18
FB52
FBB5
FBBC
FB18
FA62
FAE1
FD61
0131
047B
05CA
0547
046C
0480
0572
062D
05EF
050C
0470
049B
053D
05AE
0598
052B
04CB
04B7
04DA
04EC
04BD
045E
0418
041E
045B
0494
04B0
04C0
04C7
04AD
0479
046B
04B2
051F
054E
051E
04CE
04A0
048D
0475
0473
04B8
0513
0508
0484
042A
0492
0540
04C8
0238
FE47
FAE6
F98D
FA18
FB2C
FB99
FB37
FAA4
FA76
FABB
FB1C
FB45
FB2B
FAFE
FAEE
FB06
FB30
FB54
FB65
FB65
FB5B
FB4F
FB47
FB4B
FB5C
FB74
FB82
FB7D
FB6F
FB66
FB62
FB54
FB38
FB27
FB3C
FB65
FB6A
FB3B
FB16
FB3C
FB95
FBC1
FB9D
FB71
FB75
FB77
FB3A
FB2E
FC52
FF15
028A
050C
05C3
0546
04B5
0499
04BE
04E6
051C
055F
056F
0520
04AC
047A
049F
04D0
04D6
04C5
04BE
04AE
047A
044D
0464
04B5
04EF
04E5
04BF
04AE
04A7
048A
0473
0497
04E0
04E3
0471
03EC
03E7
046A
04EC
04FD
04BC
048B
0485
048A
04A4
0508
0573
04F1
02B4
FF31
FC0C
FAA3
FAD3
FB54
FB3C
FACC
FAB8
FB19
FB66
FB4A
FB16
FB30
FB73
FB71
FB1E
FAE9
FB12
FB55
FB54
FB23
FB1C
FB52
FB7B
FB6A
FB4B
FB4D
FB58
FB44
FB3D
FB89
FBFE
FC15
FB9B
FB10
FB07
FB6B
FBAF
FB94
FB62
FB5D
FB64
FB52
FB5C
FBB0
FBE1
FB5B
FA8A
FAFC
FDBD
01D6
04F8
05C3
0506
0486
04F5
058A
0567
04BD
0459
0480
04C4
04C3
04AD
04CD
0505
04FB
04A7
0462
0471
04BB
04FF
052D
054C
0547
0503
04A7
048B
04C9
050D
04FD
04AE
047D
0497
04C8
04D9
04D0
04C3
049C
044B
0413
0442
04A8
04AE
0431
03EB
0481
053F
046D
013F
FD21
FA79
FA49
FB57
FBD6
FB57
FACA
FAE9
FB59
FB65
FB03
FAB9
FAC8
FAEC
FAEB
FAE8
FB0F
FB42
FB50
FB4C
FB69
FB93
FB7B
FB1B
FADD
FB10
FB72
FB90
FB61
FB3D
FB47
FB42
FB0F
FAF3
FB35
FB92
FB8D
FB33
FB18
FB7C
FBD9
FBA4
FB34
FB4D
FBE5
FBFC
FB1D
FA81
FC06
FFE4
040D
062D
05F2
04FC
04C8
0548
058F
0544
04E3
04DA
04FD
04F9
04DE
04E7
04FB
04D9
0491
0489
04DB
0522
04FF
04A7
048E
04C1
04DF
04B7
0499
04C7
04FC
04D0
0466
044B
04A6
04F6
04CE
047D
0494
0506
0532
04DE
0496
04CB
0512
04BF
0418
041B
04EA
050C
02E5
FED8
FB34
F9E1
FA8E
FB73
FB77
FAFF
FAD9
FB0B
FB16
FADE
FACD
FB10
FB4B
FB2B
FAEB
FAF6
FB3F
FB5A
FB1F
FAE7
FAFB
FB2E
FB2E
FB08
FB15
FB61
FB93
FB74
FB4A
FB6A
FBB0
FBAC
FB4C
FAFF
FB11
FB3F
FB27
FAEA
FAF9
FB5A
FB8F
FB5C
FB30
FB74
FBC8
FB82
FAFD
FBB5
FE9F
02A6
0579
05DE
04D2
0429
0483
051A
052C
04EB
04E9
0527
0530
04E6
04B5
04E7
0532
0529
04DD
04B4
04CE
04E6
04C8
049C
049A
04B2
04B1
0493
0488
049F
04B0
04A1
0495
04B2
04DA
04D8
04B3
04A6
04C0
04C8
049F
0479
0490
04B8
0498
044A
046A
0529
0592
0435
00C7
FCD5
FA77
FA54
FB37
FB95
FB1D
FA9E
FABA
FB2C
FB5B
FB34
FB1C
FB43
FB5E
FB34
FAFA
FB09
FB59
FB90
FB7F
FB50
FB3D
FB48
FB4F
FB49
FB44
FB46
FB4B
FB58
FB73
FB81
FB60
FB29
FB1C
FB49
FB68
FB4C
FB33
FB6C
FBCD
FBD0
FB5B
FB04
FB4B
FBC1
FB88
FAB2
FAA7
FCBE
008D
0414
05A9
056A
04BE
04AB
050B
052B
04D7
047A
047A
04C3
0501
050F
0504
04FB
04EE
04D5
04C0
04CB
04F9
0527
052E
04FE
04B3
047E
047C
049C
04AE
0491
0461
045B
048E
04BE
04B1
0485
048C
04D1
04F4
04B0
044A
044C
04B9
04F1
0495
0434
0496
0560
04FE
0257
FE53
FB35
FA5C
FB11
FBA1
FB49
FAAD
FA9C
FB07
FB58
FB52
FB3D
FB4F
FB63
FB4C
FB25
FB19
FB20
FB0D
FAE0
FAC6
FAD5
FAF5
FB13
FB34
FB52
FB4B
FB19
FAFF
FB37
FB95
FBB2
FB79
FB44
FB5A
FB85
FB68
FB1A
FB15
FB7E
FBD6
FBA2
FB26
FB19
FB8A
FBAA
FAF2
FA40
FB3F
FE89
02A9
0560
05C6
04F2
047F
04E2
0558
053C
04CF
04AE
04F1
052B
051D
04FD
0508
051C
04FD
04BE
04AF
04DE
0508
04FF
04E5
04EB
04FB
04EE
04CF
04CA
04D4
04BE
048C
0484
04BE
04EF
04CE
048D
0496
04E1
04F3
04A3
046F
04B9
0512
04C8
0412
03FD
04E2
056C
03D5
0009
FC17
FA28
FA6C
FB52
FB82
FB0F
FAC8
FAF6
FB2E
FB19
FAE4
FAE1
FB04
FB0A
FAEA
FAE2
FB11
FB45
FB47
FB24
FB0F
FB18
FB21
FB19
FB12
FB18
FB14
FAF8
FAE2
FAF7
FB23
FB2C
FB04
FAE4
FAF3
FB06
FAEE
FADD
FB2A
FBB3
FBE2
FB7E
FB1F
FB64
FBF2
FBCE
FAEE
FADC
FD26
014C
04E7
061A
0559
0483
049D
0517
0518
04B9
04A5
04FD
0537
0507
04CA
04E5
052C
052C
04DE
04A4
04AD
04C7
04C9
04D6
0512
054D
053E
04F6
04C9
04DB
04F5
04EC
04E2
0503
0524
04FD
04A9
0494
04D9
050D
04D1
0470
0477
04E3
0507
0494
0432
04A7
0573
04E2
01EE
FDB9
FAAA
FA07
FAE3
FB77
FB24
FAAB
FAC9
FB31
FB31
FAC0
FA7D
FAB5
FB0B
FB19
FB03
FB1F
FB5D
FB66
FB33
FB1B
FB47
FB6C
FB44
FAF7
FAE0
FAFC
FB05
FAF2
FB0C
FB61
FB89
FB3F
FADF
FAEB
FB46
FB62
FB1B
FAF8
FB56
FBC4
FBA1
FB24
FB1C
FBAA
FBDB
FB0F
FA51
FB83
FF22
0360
05E1
0602
051C
04C0
0527
0589
0567
0513
0508
053A
054D
0529
050B
051A
052E
050F
04CB
049F
04A5
04B5
04AE
04A5
04BB
04E3
04EF
04DF
04D9
04E8
04E6
04C1
04A5
04B9
04D6
04B8
0470
0465
04B8
0502
04D7
0473
046B
04C2
04DA
0476
043A
04A8
04EA
036B
FFD2
FBE3
F9DB
FA27
FB2C
FB53
FAA3
FA2B
FA6E
FAEF
FB17
FAEC
FACB
FAD6
FAEB
FAF0
FAF5
FB06
FB19
FB27
FB3A
FB4E
FB4C
FB33
FB20
FB1B
FB0A
FAEA
FAF3
FB49
FBB3
FBD7
FBA9
FB74
FB72
FB88
FB7A
FB49
FB33
FB5D
FBA4
FBC3
FBA2
FB64
FB43
FB5D
FB94
FBA8
FB86
FB7E
FBD8
FC42
FC0E
FB41
FB15
FCE2
007B
040B
05C8
059F
04F5
04EE
0569
05A4
0567
051F
051E
0542
0547
0527
0508
04FC
04F9
04EE
04DD
04D9
04F3
051E
052F
0504
04B8
0494
04BC
04EA
04C4
0464
0442
048F
04EA
04EC
04B5
04AB
04E0
04FF
04D6
048E
046A
046E
047D
0493
04B5
04C1
049D
047D
04A3
04DC
04B0
0440
0449
04EC
04EB
02D4
FEF0
FB63
FA08
FA9F
FB69
FB4E
FAC4
FAA2
FAE2
FAED
FAA7
FA82
FAB1
FAE5
FADD
FAC7
FAED
FB3B
FB5F
FB3A
FAFF
FAEB
FB04
FB2B
FB4B
FB59
FB55
FB5A
FB8A
FBCA
FBC4
FB5F
FAF5
FAF0
FB45
FB92
FB9D
FB80
FB6D
FB6E
FB6E
FB62
FB4C
FB2F
FB1D
FB34
FB6B
FB80
FB54
FB43
FBA9
FC1F
FBCF
FADB
FAD8
FD36
015E
04F3
0631
0587
04B2
04B3
0520
054A
0534
053C
0555
0533
04E7
04CD
04F7
0519
0505
04E5
04EC
050B
051B
0513
04FE
04DE
04BA
04B3
04DF
0503
04D0
0465
0447
04A4
0508
0501
04C1
04C0
0504
0523
04EA
04A1
0494
04B1
04BA
04A9
049E
0497
047B
046F
049D
04C7
0488
0425
0466
0541
0534
02C8
FE95
FAFF
F9D2
FA89
FB4F
FB32
FABE
FAB3
FAED
FAE9
FAB5
FABD
FB09
FB36
FB21
FB14
FB3E
FB6D
FB64
FB36
FB21
FB3A
FB5A
FB5C
FB41
FB19
FAF6
FAF9
FB37
FB7F
FB7E
FB32
FAF8
FB07
FB24
FB11
FAF9
FB24
FB7B
FBA9
FBA0
FB99
FBAF
FBB2
FB84
FB61
FB7B
FB96
FB6C
FB45
FB8F
FBF7
FB9C
FAA1
FAB6
FD52
01A8
052B
0634
057C
04D6
0506
0564
0549
04F7
04EF
0515
0507
04D3
04D2
04FF
04FE
04BF
0496
04B5
04E2
04D6
049F
047A
047E
048D
0499
04B2
04D2
04D5
04B7
04AA
04C0
04CD
04C0
04C8
04F8
050E
04D5
047F
0460
046E
0461
0434
0432
046E
0496
0479
046C
04BD
0507
04B0
040A
041B
04E2
04B7
0226
FE0B
FAED
FA45
FB1F
FB9E
FB37
FACC
FB08
FB7B
FB7F
FB34
FB1B
FB36
FB2B
FAF9
FAFB
FB3F
FB6A
FB45
FB0C
FB0C
FB37
FB4E
FB43
FB41
FB5B
FB6F
FB66
FB5D
FB6C
FB7F
FB84
FB88
FB8F
FB7A
FB48
FB32
FB5A
FB8F
FBA1
FBA8
FBC8
FBD8
FBA4
FB61
FB7C
FBEF
FC20
FBBE
FB53
FB7E
FBCD
FB52
FA64
FAE4
FE05
026D
056C
05DA
04FC
0496
04EC
051F
04C5
046D
048B
04CF
04D0
04C0
04FA
0550
0555
0514
04F8
0518
051F
04E6
04AD
04AF
04C8
04B6
0485
0473
0482
047B
0455
0451
0486
04AC
0499
0487
04AE
04DA
04C0
0471
0437
0423
041A
0427
046B
04C6
04E1
04B6
04A5
04DC
04E6
0469
03F8
046C
054A
04B6
01A7
FD7E
FABC
FA52
FB01
FB3A
FAD9
FAAD
FAFE
FB3F
FB0F
FAC3
FAC5
FAF1
FAF5
FAEB
FB1C
FB6F
FB8A
FB64
FB44
FB4C
FB5B
FB58
FB55
FB5E
FB5B
FB47
FB46
FB6C
FB86
FB5F
FB1F
FB20
FB58
FB5B
FB0C
FADC
FB16
FB6F
FB81
FB6B
FB7D
FB9F
FB83
FB3E
FB37
FB76
FB81
FB2B
FB0B
FB94
FC20
FBBD
FAF2
FBAB
FEDD
02F5
0575
05B4
0527
0533
05A8
05A0
0508
049A
04AA
04C7
0499
0477
04BA
0513
050D
04CC
04D0
0523
055B
0542
0510
04FE
04FC
04E7
04CA
04B9
04A9
048D
0481
04A5
04D5
04CB
049F
04AE
0504
0534
0506
04D0
04E8
051A
0511
04EB
04F1
0501
04BC
043F
0417
0467
0492
0432
03EF
0490
0553
044A
00CC
FCB2
FA6E
FA6E
FB23
FB40
FAF7
FAFE
FB4A
FB50
FAFF
FAD1
FAED
FAEE
FAA9
FA8C
FAE7
FB51
FB4A
FAFE
FAF0
FB26
FB3D
FB16
FAFD
FB1B
FB3B
FB2E
FB1D
FB3B
FB67
FB60
FB3C
FB45
FB70
FB5B
FAF9
FAC2
FAF6
FB39
FB30
FB14
FB3C
FB7A
FB73
FB49
FB71
FBE2
FC14
FBDF
FBD5
FC44
FC74
FBA7
FAB5
FB9B
FEFF
0307
054C
0568
04DA
04DA
053C
0554
051D
04FC
0500
04E8
04B9
04C4
0509
0521
04EE
04D8
051A
054C
0510
04B6
04BE
0507
0512
04D6
04C6
050A
053C
050A
04B9
04B3
04E0
04D3
048D
0481
04C9
04EB
04A4
045C
0470
0494
0465
0425
0448
04A5
04AF
0463
0459
04BC
04E3
0463
03FA
0487
0549
0438
00A0
FC6B
FA26
FA40
FB13
FB33
FACC
FAAE
FAFA
FB2F
FB15
FAF4
FB02
FB19
FB14
FB11
FB1C
FB09
FAD1
FAC4
FB07
FB43
FB2E
FB09
FB2F
FB72
FB64
FB0D
FAE9
FB2C
FB76
FB69
FB33
FB36
FB63
FB5C
FB26
FB2E
FB82
FBAD
FB81
FB6D
FBB4
FBE1
FB8C
FB25
FB4D
FBC3
FBB8
FB26
FB02
FBB8
FC3D
FB90
FAAD
FBDA
FFA7
03CF
05BE
0565
04B6
04E5
055C
053B
04BB
04A2
0504
054B
052F
050A
0520
052E
04FF
04D9
0500
0533
051B
04E2
04DD
04F2
04C9
0477
046E
04CC
0525
051C
04DC
04C7
04E4
04E5
04B3
0490
049D
04AA
0494
0482
0486
046F
043D
0446
04A4
04E4
04AB
045E
0490
0504
04EF
0447
0418
04EE
057F
03DD
FFFD
FC29
FA7C
FAB4
FB1C
FAE0
FA8E
FAB6
FB0A
FB0D
FADD
FAD8
FAF2
FADC
FAAC
FAC7
FB2F
FB63
FB2C
FAFE
FB2F
FB64
FB2F
FAD3
FADE
FB3C
FB56
FB04
FACB
FB0E
FB79
FB80
FB27
FAEB
FAFF
FB13
FAF2
FADD
FB0C
FB49
FB5B
FB63
FB8C
FBA4
FB7A
FB4B
FB6D
FBB4
FBB2
FB77
FB80
FBD6
FBC6
FB02
FAAF
FC6C
0033
03F1
05AA
057A
04F0
0501
055B
056A
053B
0523
052E
0531
0533
0551
056A
053D
04EA
04DA
0519
0531
04EE
04BD
04FF
0560
0553
04EF
04C9
0506
0524
04CB
0453
044E
04B6
0507
04FD
04DA
04DD
04E2
04C0
04A0
04AD
04BF
04AA
0495
04B3
04DD
04CD
04A1
04A4
04C0
048E
0419
0412
04BB
04FB
0347
FFA1
FC06
FA63
FAA4
FB36
FB0F
FA8E
FA79
FADE
FB34
FB2A
FAEE
FAC7
FAC3
FAD3
FAEF
FB06
FAF7
FACD
FAB9
FAC8
FAC4
FAA1
FAAB
FB11
FB79
FB74
FB1A
FAF4
FB3A
FB8B
FB7A
FB1F
FAE8
FAF6
FB0B
FB00
FAFE
FB21
FB3E
FB31
FB29
FB57
FBA2
FBD3
FBE9
FBEC
FBBC
FB52
FB10
FB5C
FBE2
FBC7
FAF9
FADF
FD00
00FB
0487
05D4
055A
04D6
0511
0560
0519
04A8
04CE
0570
05C3
0574
050F
0519
0553
0538
04D0
0499
04C9
050F
051D
0504
04F7
04FA
04FB
0504
052C
055B
0554
050B
04BA
049A
049A
048D
0478
0486
04B6
04D3
04C1
04A9
04BC
04DE
04C3
0462
042D
048A
050A
0473
01EA
FE21
FB00
F9E5
FA66
FAFE
FACB
FA55
FA7E
FB2B
FB79
FB0D
FA8C
FAA5
FB1B
FB46
FB14
FB14
FB81
FBD6
FB93
FAFE
FAC7
FB15
FB5C
FB39
FAF1
FAE9
FB09
FAFE
FAD3
FAE2
FB39
FB7D
FB72
FB4C
FB4E
FB5B
FB36
FAFF
FB0F
FB62
FB89
FB5F
FB4C
FB8E
FBB1
FB3C
FAE0
FC24
FF9A
03C5
065A
0688
0595
0528
0585
05CC
057B
0511
0524
057F
0584
0517
04BB
04C9
04FB
04E6
04A0
048E
04C8
04F5
04D4
0495
0492
04CC
04FB
04F6
04DB
04CB
04C2
04BB
04CF
050A
0534
0513
04C1
0493
04A5
04B8
04A5
04A6
04EF
052F
04E3
043B
041B
04D6
0544
03B7
0000
FC02
F9E6
F9F9
FAB6
FAC0
FA41
FA2A
FAB0
FB20
FAFA
FA9E
FAA5
FB03
FB30
FB02
FADF
FB19
FB6E
FB73
FB31
FB0E
FB35
FB68
FB6A
FB55
FB5C
FB74
FB72
FB5B
FB5D
FB76
FB6B
FB2D
FB06
FB2B
FB66
FB61
FB31
FB38
FB80
FB8F
FB23
FAC0
FB08
FBAB
FBAB
FAEF
FAF4
FD4B
017E
052A
0664
0599
04B5
04D2
055F
056D
0510
0500
055D
0587
0525
04A4
0491
04D3
04EF
04CF
04D2
051C
054F
051F
04C6
04AD
04D2
04E5
04D8
04F1
0538
054F
04F8
0484
046E
04A8
04B7
047B
0460
04A6
04E3
049F
0429
0439
04DA
0534
04C4
043F
049B
0563
04C8
01B7
FD6D
FA64
F9CC
FA97
FB0D
FABA
FA70
FACC
FB68
FB98
FB55
FB1E
FB22
FB18
FAD5
FAA1
FAC4
FB10
FB20
FAF1
FAE2
FB1A
FB53
FB40
FB03
FAEB
FAFD
FAFC
FAE0
FAF4
FB59
FBB9
FBAF
FB5B
FB35
FB5E
FB7B
FB57
FB41
FB8B
FBE7
FBCC
FB4E
FB25
FB92
FBD3
FB3D
FAA4
FBDC
FF7B
03B8
0615
05F5
04EF
04B3
053E
0575
04F5
047B
04A8
0521
053A
04F6
04D5
04ED
04D4
046D
043F
04B4
056C
05AE
055F
050B
050E
051F
04ED
04B2
04D3
052A
0536
04E3
04AD
04E3
052C
050C
04A8
0488
04C4
04E6
04B5
0497
04DF
051B
04B6
0407
0414
04F8
052D
030D
FEEF
FB23
F9A4
FA36
FB13
FB15
FAA8
FAAF
FB37
FB96
FB7A
FB3D
FB3F
FB59
FB36
FAF0
FAEC
FB39
FB6C
FB3B
FAE7
FAE8
FB3E
FB78
FB51
FB01
FADB
FADE
FAD0
FAB5
FAC7
FB0E
FB38
FB06
FAB6
FAB0
FAFE
FB4B
FB69
FB7D
FB96
FB7D
FB26
FAFD
FB56
FBBA
FB5C
FA81
FAD5
FDB0
022D
05AC
0680
058A
04D7
052A
0591
052A
046B
044D
04D2
0526
04E8
04AD
04F7
0562
0544
04C0
048E
04EE
0553
0541
04F2
04DE
0505
0503
04C9
04BA
0503
0546
0526
04D3
04BA
04D9
04DA
04AB
049D
04CB
04E4
04B1
0488
04D4
054E
0540
04A2
0461
0515
05BA
0479
00D2
FC8F
FA1D
FA2B
FB40
FBA2
FB17
FA9B
FAD2
FB48
FB53
FB0A
FB09
FB77
FBC6
FB80
FAE4
FA86
FA8F
FAAA
FA9E
FA9F
FAE4
FB39
FB42
FB04
FAE1
FB07
FB3B
FB46
FB47
FB6C
FB8E
FB6A
FB19
FAF9
FB21
FB3B
FB0F
FAE3
FB07
FB40
FB26
FAF2
FB45
FC06
FC27
FB2C
FA6E
FBF7
FFFE
0433
0617
0590
049A
04AD
0549
0540
048F
0432
049D
0530
054A
0523
0540
058D
0586
051A
04D2
0503
0550
0542
04F3
04D1
04E5
04D2
0483
045C
049F
04FA
04FE
04C5
04CD
0531
0572
052F
04AF
0478
048A
047F
044B
0462
04E9
0546
04E6
0444
046F
0562
056F
02F9
FE94
FAD4
F9B3
FAAC
FBAA
FB81
FAD8
FAB7
FB14
FB2F
FADF
FAC1
FB20
FB6B
FB0F
FA63
FA3B
FAC3
FB4D
FB55
FB25
FB34
FB5F
FB33
FAC2
FA9D
FAFA
FB58
FB3F
FAF0
FAF7
FB4B
FB5C
FAFA
FAAC
FAE3
FB54
FB77
FB57
FB67
FBAC
FBAA
FB49
FB2A
FBB6
FC36
FBB1
FA97
FADA
FDC5
022F
0572
0628
054E
04BA
04FF
0555
0523
04D3
04FA
0560
055A
04D8
0484
04CD
054C
055A
04F5
04AD
04CE
050A
050B
04F1
0509
0543
0545
04FC
04C1
04D7
0509
0501
04CC
04BA
04D4
04D0
048F
045A
046C
0492
0482
0466
049E
0501
04F2
0452
03F3
0477
0504
03D3
005A
FC56
FA1B
FA32
FB18
FB46
FAC4
FA89
FAEF
FB60
FB64
FB42
FB5F
FB8B
FB51
FAC7
FA79
FAAB
FB05
FB22
FB0A
FB01
FB0D
FB07
FAF4
FB04
FB3A
FB4D
FB17
FAD5
FAD4
FAFE
FB0D
FB05
FB37
FBB0
FC0B
FBF1
FB98
FB7B
FBA9
FBAF
FB56
FB11
FB5E
FBEB
FBE0
FB2C
FB21
FD2B
010B
04B4
063B
05A8
049D
046D
04F0
0542
0517
04E8
0506
0522
04EE
04B2
04D9
0546
056F
052C
04EA
0505
053B
051D
04BB
048A
04B1
04D9
04CF
04DB
0534
0584
0557
04D4
048F
04B3
04C1
0463
0401
0427
04A9
04D0
0472
042E
0468
049F
0445
03CB
041C
0501
04DB
0267
FE73
FB3B
FA22
FA8B
FAF7
FACD
FA8A
FAAB
FB01
FB2C
FB37
FB60
FB9C
FB9D
FB55
FB11
FB0D
FB22
FAFF
FAAA
FA78
FAA0
FAFC
FB47
FB68
FB68
FB42
FAF6
FAAE
FAB3
FB12
FB7F
FBA2
FB83
FB73
FB9E
FBCC
FBBA
FB7B
FB57
FB5C
FB53
FB32
FB38
FB82
FBAD
FB5F
FB22
FC3A
FF40
0312
05AC
0621
0559
04CB
04E4
0501
04B5
0462
0487
04EE
0510
04E5
04EF
055D
05B0
0575
04EE
04B2
04DC
04FD
04D6
04A1
049E
04A9
048B
0470
04AC
0520
0542
04DF
046C
0466
04A4
04A5
0459
0430
0461
049B
048B
0466
0482
04B3
0487
041E
0430
04E4
0513
0352
FFBE
FC30
FA71
FA8E
FB2C
FB39
FADE
FAC5
FB08
FB31
FB0D
FAEB
FB19
FB64
FB64
FB0C
FAB4
FAA6
FAD9
FB19
FB4F
FB76
FB7E
FB5A
FB2C
FB2E
FB64
FB88
FB68
FB2F
FB30
FB77
FBBA
FBBE
FB9F
FB9A
FBB1
FBB1
FB91
FB81
FB96
FB96
FB5A
FB1F
FB36
FB6A
FB2D
FA9C
FAE4
FD2B
0101
0471
05D8
0571
04C7
04D8
0542
0543
04E2
04BA
04F5
051B
04D8
047E
047E
04BF
04D2
04A5
049B
04E5
0531
052E
04FC
04E6
04DE
049E
043D
0428
0484
04DE
04C2
045B
042F
0465
049D
0499
0497
04CB
04EA
04A2
0443
046A
050B
0556
04DA
044D
04A0
056D
04F6
021C
FDE5
FA99
F98D
FA22
FAEE
FB39
FB3B
FB41
FB38
FB0E
FAFE
FB3E
FB95
FB9D
FB4D
FB07
FB14
FB4F
FB6E
FB5F
FB49
FB3F
FB3B
FB46
FB75
FBB5
FBC7
FB8E
FB4C
FB54
FB92
FBA7
FB6F
FB36
FB43
FB63
FB37
FADC
FADC
FB56
FB9D
FB1A
FA76
FB47
FE51
025B
0535
05DD
053E
04D8
0517
055A
052D
04E3
04EA
051B
0503
04A9
0483
04B6
04DE
04B2
0480
04B7
0531
055A
04FE
0488
046A
048E
049C
0487
047E
047E
044E
0405
0411
0492
0501
04E3
047A
046E
04C2
04D2
0463
0432
04D9
0579
044E
00DD
FCDF
FA98
FA86
FB40
FB5F
FAEE
FAB9
FAFD
FB3D
FB2F
FB21
FB4E
FB69
FB1F
FAB9
FAC5
FB3D
FB82
FB3C
FAD5
FADD
FB40
FB6D
FB29
FAD7
FAE6
FB3E
FB7E
FB80
FB68
FB46
FB0E
FADD
FAF1
FB41
FB68
FB2C
FAE9
FB17
FB71
FB2D
FA43
FA14
FC30
0067
048A
0669
05E4
04AD
0448
04AC
04F7
04CC
049E
04C9
0509
04FF
04CF
04DB
0514
050C
04AA
0468
04AE
052F
0550
04FB
04B1
04C5
04E9
04B3
0448
042C
0484
04E6
04EC
04B4
0494
04A5
04CC
0503
053A
052A
04A1
0416
0455
054A
0578
035A
FF55
FBB3
FA59
FAE3
FB78
FB15
FA70
FA92
FB59
FBD1
FB97
FB3B
FB42
FB71
FB59
FB18
FB18
FB4B
FB3A
FAC7
FA74
FAAF
FB30
FB60
FB25
FAEF
FB09
FB3C
FB46
FB48
FB7C
FBC1
FBBF
FB70
FB21
FAFB
FADE
FACE
FB16
FBBC
FC14
FB79
FA81
FADF
FD9D
01B4
04D8
05BB
051B
0493
04C8
0524
0509
04A7
0487
04B7
04CE
04A7
048E
04C2
0509
0506
04C5
04A5
04CF
0505
0503
04DD
04D4
04EE
04F6
04D5
04B1
04AB
04B3
04AC
04A3
04AF
04B9
04A6
0493
04BC
0505
0500
048E
0442
04A7
052E
045D
0173
FD96
FAEE
FA75
FB2A
FB7C
FB0A
FAA2
FAD7
FB48
FB5D
FB26
FB20
FB52
FB4A
FAE4
FA95
FABD
FB15
FB26
FB02
FB21
FB96
FBDF
FB98
FB0B
FAC3
FAD1
FADF
FAD1
FAEB
FB41
FB7E
FB65
FB41
FB66
FB97
FB62
FAF0
FAEE
FB6E
FB8B
FAAB
F9E2
FB25
FEF7
0367
05F1
05FF
0515
04C0
050A
0528
04E1
04B6
04ED
0528
0510
04E9
050A
053C
050C
0495
0478
04F3
0574
055B
04CB
046E
048A
04BF
04AE
0480
0488
04B7
04C4
04B1
04C4
04FC
04F7
0491
0442
0474
04D5
04C1
0457
0481
0581
05FE
0433
0021
FBFD
FA08
FA58
FB2C
FB27
FA99
FA7D
FAF2
FB3B
FAFD
FAB0
FAC7
FAFB
FAD0
FA72
FA86
FB23
FB9A
FB65
FAE5
FACC
FB20
FB4C
FB0E
FAD5
FB0C
FB75
FB8C
FB4E
FB27
FB3C
FB42
FB1B
FB20
FB7E
FBBE
FB6D
FAF1
FB17
FBC0
FBD3
FAE4
FA65
FC49
0078
047A
0608
0569
04A9
04F8
05A0
058E
04EC
04AB
04FB
0523
04C2
0472
04CE
0575
0594
051C
04CA
0503
0550
0522
04B1
0499
04F0
0533
0516
04E6
04FB
0528
051F
04FD
050E
052B
04E2
0445
0407
0481
050B
04D3
042A
0432
051C
0555
032F
FF10
FB59
F9EF
FA70
FB1B
FAFC
FA98
FAA9
FB01
FB02
FAB4
FAB4
FB2B
FB80
FB2E
FA8A
FA51
FAA8
FB01
FAF4
FAC0
FACF
FB0C
FB0F
FAC8
FA94
FAB6
FAFF
FB27
FB34
FB51
FB6B
FB4D
FB0A
FAF8
FB28
FB47
FB24
FB17
FB67
FBA8
FB38
FA7B
FB02
FDE1
0215
053E
0603
054C
04DC
0536
0581
0519
0484
0491
0525
0577
0540
050A
053F
057C
0535
0495
0451
04B2
0545
0586
0574
054D
0518
04B7
044F
043C
048E
04EC
050F
0511
0518
0505
04C0
0491
04C3
050C
04D2
0429
040D
0508
05F7
04D9
0126
FCC4
FA41
FA42
FB43
FB9A
FB26
FAC9
FAE8
FB09
FAC8
FA79
FA9B
FB15
FB57
FB27
FAD7
FAC0
FAD6
FAE3
FADE
FAE3
FAF5
FB01
FB12
FB39
FB5C
FB42
FAF6
FACB
FAEF
FB16
FAEE
FAAB
FAD0
FB66
FBCF
FBA4
FB5C
FBA8
FC46
FC25
FAF7
FA2F
FBB0
FF8B
039A
059D
0563
0491
0488
051F
0574
054C
0526
0549
055B
04FE
046E
042F
0462
04BE
050D
0552
057A
054F
04DA
048D
04BD
0526
0544
050A
04EA
051D
0546
050A
04AF
04B3
04F6
04DB
0447
03F6
0466
04FE
04D6
042D
0434
0533
058A
0366
FF28
FB5A
FA08
FABC
FB81
FB53
FAD1
FAD0
FB22
FB20
FAC5
FA9E
FADF
FB21
FB22
FB2D
FB74
FB8D
FB0D
FA4D
FA21
FAB2
FB44
FB3B
FAE6
FAEC
FB47
FB5C
FB02
FACF
FB26
FB90
FB6B
FAF0
FAE1
FB5F
FBB4
FB79
FB4C
FBCF
FC6D
FBF7
FA9F
FA65
FCF8
0174
0517
0620
055E
04BE
0501
056C
0557
051A
0545
059A
0578
04E2
0484
04B6
050A
0508
04E7
051A
0582
058E
051E
04C7
04F5
0540
050C
0479
0441
049E
04F5
04BB
0443
043C
04A5
04DF
04AC
048C
04CD
04F2
047D
03F8
045A
054F
0504
022E
FDF5
FAF7
FA78
FB39
FB52
FA81
F9FA
FA6E
FB24
FB31
FABF
FA9D
FAF4
FB25
FADE
FA95
FABE
FB06
FADD
FA6D
FA63
FAEF
FB72
FB6A
FB25
FB34
FB83
FB88
FB29
FAFB
FB56
FBCC
FBC4
FB5F
FB30
FB52
FB55
FB1F
FB30
FBBE
FC01
FB3B
FA3F
FB11
FE95
031E
05EC
0604
04E0
0467
04E3
054E
0519
04CE
0508
0580
058E
052E
04FA
053B
058F
0588
0548
0531
054B
054C
051D
04FA
0504
0504
04D2
04A5
04C4
0508
050C
04BE
047E
0484
0492
0468
0443
0483
04EE
04DC
0445
0410
04D6
0596
046F
00D1
FC8B
FA20
FA41
FB5F
FBB0
FB06
FA6E
FA8B
FAED
FAEE
FA9C
FA79
FAB2
FAF7
FB01
FADD
FAB5
FA90
FA7A
FA97
FAE7
FB1B
FAF1
FAA3
FAA5
FB07
FB57
FB46
FB19
FB36
FB7D
FB6C
FAF4
FAA5
FAE1
FB4E
FB69
FB5C
FBB1
FC46
FC35
FB34
FA91
FC17
FFE2
03E4
05D9
057C
0466
0418
04A5
0543
057E
0586
058E
0581
054A
050F
04ED
04C9
0495
0493
04FA
0583
05A6
0551
0504
0520
0562
054F
04F7
04E4
053F
058A
0550
04D5
04A8
04CA
04B6
043C
03E0
0413
0480
048C
0454
048B
052B
04EF
02A8
FEEC
FBD2
FAD1
FB5E
FBDA
FB80
FAEB
FADE
FB32
FB41
FAE6
FA93
FA8E
FAA1
FA93
FA91
FAD2
FB27
FB2E
FAF2
FAE0
FB26
FB6A
FB52
FB08
FAF0
FB07
FAF9
FAC3
FAD7
FB67
FBF2
FBDD
FB4C
FAF2
FB0D
FB1E
FAD0
FAA8
FB3F
FC15
FBFD
FAE9
FA9C
FCE4
0149
052F
0677
058A
046C
045B
04E3
051E
050A
053B
05C3
060B
05B5
051E
04D0
04D6
04E0
04D8
04E8
0510
0512
04DD
04B7
04C9
04D5
049A
0455
0479
04F5
0524
04B7
0438
0453
04D7
04FD
04A1
0496
055E
05F4
04A8
0132
FD5A
FB31
FAF1
FB27
FAB5
FA05
FA16
FAE5
FB6C
FB09
FA4A
FA19
FA93
FB08
FAFE
FABB
FABE
FB0F
FB57
FB5D
FB3C
FB1F
FB1A
FB3D
FB92
FBE3
FBCE
FB3D
FAA6
FA93
FAEF
FB24
FAF6
FAE8
FB6F
FC12
FBDE
FAD9
FA7E
FC55
001C
03D8
05B4
05A3
04F2
04AA
04CA
04E6
04F8
053C
0598
059B
0526
04AF
04B1
0514
0556
053C
050B
0513
053C
0534
04E5
048C
0468
047F
04B8
04F8
051C
04FE
04AA
047D
04BD
0524
0517
0479
0409
0482
0565
0518
0288
FE8B
FB41
FA16
FA96
FB4A
FB5C
FB1A
FB15
FB41
FB30
FAD1
FA8E
FABB
FB2B
FB7A
FB85
FB6F
FB51
FB21
FAE0
FAAD
FA9D
FA9E
FAA9
FADA
FB3D
FB91
FB7D
FB09
FAB0
FACA
FB23
FB53
FB66
FBC7
FC6C
FC91
FBAD
FA9F
FB37
FE4F
028B
0578
05E9
04DE
0420
0455
04CC
04D9
04AF
04D2
0530
0545
04F7
04BD
04E8
0529
0512
04BE
04A8
04F1
0530
0516
04DE
04E4
0518
0522
04FC
04F3
0522
0536
04FA
04C0
04E6
0520
04CE
0406
03C2
0489
053C
03FB
0058
FC32
F9ED
FA16
FB24
FB7E
FB19
FAE5
FB3D
FB84
FB3E
FAD4
FAF0
FB75
FBA8
FB3D
FAB6
FA9E
FACE
FAC9
FA81
FA66
FAB0
FB13
FB3C
FB42
FB64
FB86
FB5D
FAF9
FAC4
FADF
FAEA
FAB5
FAAE
FB3C
FBDC
FB95
FA80
FA48
FC8C
00D2
04BC
0657
05E2
050B
04E6
0522
0515
04C8
04B8
04F3
0510
04DB
04A7
04C4
0505
0511
04F4
0503
054A
056F
0546
051F
0548
057F
053E
0490
0427
0476
050E
0537
04F1
04DA
0524
0527
0471
03BD
0428
0563
057B
02F3
FEAB
FB2C
FA0B
FA94
FB1B
FAFB
FAC0
FAD9
FAE8
FA93
FA3F
FA7B
FB0E
FB3D
FAE6
FAB5
FB1F
FBAB
FB96
FAF2
FA88
FABF
FB1F
FB1C
FAE4
FAF8
FB4D
FB51
FADE
FA85
FABE
FB35
FB50
FB26
FB66
FC25
FC70
FB85
FA4D
FAD6
FE14
0281
0579
05D8
04D5
045B
04F0
059B
0584
04FF
04E0
0542
057E
052E
04AF
0483
04A5
04B4
04A1
04B4
0501
052F
04F8
0497
047D
04B3
04E9
04FB
0517
054F
055D
051D
04E1
04F6
0514
04AC
03E7
03B2
0477
051B
03EF
00A6
FCF8
FAEB
FAD3
FB58
FB3F
FAA9
FA76
FAF0
FB80
FB85
FB12
FAAC
FAA9
FAEF
FB3B
FB5F
FB4A
FB0A
FAD7
FAF3
FB61
FBCF
FBE5
FBA0
FB44
FB0F
FB01
FB07
FB1B
FB2B
FB05
FA99
FA4B
FAAF
FBB5
FC67
FBE2
FAA6
FA81
FCD2
00E9
0482
05EC
0579
04BA
04A3
04E0
04DA
04B2
04E7
056F
05A7
0539
0492
0453
048E
04D6
04EA
04ED
0500
04FC
04C4
0490
04A4
04DE
04E3
04B0
04A3
04ED
053E
0539
04FD
04F6
0528
0526
04D1
04B9
0548
05C2
04A3
0160
FD58
FABA
FA66
FB46
FBB7
FB47
FAC3
FAD7
FB2A
FB01
FA61
FA07
FA6A
FB1F
FB75
FB4D
FB20
FB3F
FB76
FB71
FB3B
FB18
FB10
FAEC
FAAA
FA98
FAE4
FB55
FB91
FB8C
FB71
FB4D
FB17
FB05
FB69
FC0D
FC21
FB39
FA53
FB2F
FE69
0280
0538
05BF
051F
04BB
04E3
0510
0503
050F
0562
059D
0562
04F0
04D1
0515
0542
0504
0496
0467
048A
04BE
04DB
04F6
051E
0535
0526
050A
04FE
04EA
04B5
048A
04A2
04CF
0490
03CC
0345
03D1
0519
0581
03A1
FFE0
FC44
FA8A
FAAA
FB46
FB53
FAFA
FAE4
FB2D
FB5A
FB1F
FAC9
FABB
FADE
FADC
FAB4
FAC5
FB30
FB92
FB86
FB31
FB06
FB1B
FB10
FAB3
FA65
FAA3
FB4D
FBC4
FBAC
FB46
FAF7
FAD6
FADB
FB2C
FBD9
FC5B
FC05
FB29
FB55
FDCE
01DB
051F
05F1
04F6
0420
046D
0528
054B
04E5
04C1
051C
0561
0523
04C1
04C3
04FC
04D7
0453
0419
048E
053A
0569
0520
04FC
053E
0575
053D
04DC
04CC
04FD
04EE
0489
044B
047C
04AE
0470
042A
0499
0568
04FB
0228
FDE6
FAA0
F9CF
FAA7
FB53
FB08
FA6F
FA55
FAA6
FADE
FAF0
FB33
FBAB
FBDF
FB91
FB21
FB07
FB29
FB1A
FAD7
FAD3
FB3E
FB9F
FB6D
FAD8
FA8F
FAE1
FB66
FB9E
FB85
FB5B
FB2A
FADE
FABD
FB26
FBD4
FBD5
FAD0
FA08
FB6E
FF60
03D2
0628
05CB
0480
043B
051C
05D8
0594
04CC
0468
0496
04DB
04EB
04EE
0509
0513
04EF
04CE
04E6
0508
04E1
048D
0483
04DE
0523
04E6
0474
0474
04F0
0548
0516
04BA
04B2
04C8
0476
03FD
0448
056D
05DE
03CB
FF74
FB52
F9A9
FA51
FB49
FB2D
FA6F
FA2C
FA90
FAE4
FAC8
FAAF
FB06
FB7E
FB8B
FB38
FB0A
FB2E
FB47
FB11
FAD5
FAEF
FB37
FB3F
FB00
FAEB
FB35
FB7C
FB60
FB1D
FB2D
FB84
FB96
FB3E
FB0E
FB6D
FBC9
FB4D
FA60
FAC4
FDB4
0223
0583
0645
053E
046A
04B8
0579
05B7
056A
0530
054B
0566
0548
052E
0558
058C
0560
04DA
0472
047D
04CC
0508
051A
0525
0528
04FD
04A9
046F
0474
0490
0494
0496
04BC
04D2
047D
03EA
03DD
04B4
0574
046D
010C
FCD9
FA32
FA11
FB4C
FC05
FB89
FA9A
FA2D
FA63
FABD
FAE7
FAF8
FB12
FB27
FB2B
FB33
FB41
FB27
FAC9
FA71
FA8F
FB22
FBAA
FBBD
FB83
FB66
FB6F
FB4D
FAED
FAB4
FAF0
FB59
FB83
FB84
FBCB
FC42
FC25
FB2B
FA81
FBDC
FF78
0381
05D8
061D
059D
0579
0589
0531
0491
045A
04AF
04F7
04CA
048F
04C6
0531
0531
04C3
048A
04CE
050B
04C3
044F
0467
04FF
0544
04D4
045D
049F
054B
0572
04DF
0464
0490
04DD
0489
03E8
0409
04FD
052B
02FC
FEEE
FB54
FA02
FA9B
FB67
FB55
FAC7
FA99
FAEB
FB34
FB25
FAFE
FB0F
FB3D
FB46
FB3A
FB5D
FBAA
FBC0
FB6E
FB06
FAF8
FB3B
FB53
FB06
FAAB
FAA8
FADE
FAE9
FACB
FAED
FB65
FBB7
FB8C
FB43
FB68
FBBF
FB89
FADC
FB27
FDAF
01C2
0512
060D
0559
04B7
04EA
054E
0534
04DC
04E0
053A
0564
052C
04EC
04EB
04FB
04E0
04C0
04DB
0513
051A
04FC
050D
0550
055F
0504
04A5
04C2
053C
056D
050A
048D
0481
04BF
04B5
045A
044C
04CD
0508
03C6
00E2
FDA8
FB90
FADF
FAB5
FA67
FA37
FAA2
FB60
FB98
FB09
FA71
FA92
FB33
FB85
FB3D
FADE
FADC
FAEE
FA9F
FA2B
FA3C
FAE0
FB58
FB22
FAB1
FABB
FB32
FB6D
FB30
FAF0
FB06
FB1E
FADE
FA9D
FAF4
FBAC
FBDA
FB4C
FB46
FD31
00C6
0421
05A8
057C
04E7
04CE
0504
0503
04C5
04B9
050F
0563
0542
04C8
0491
0500
05BB
05F8
0569
04A7
047F
04F4
054A
0519
04DA
051E
05AB
05BC
0517
0450
03FD
0409
0421
0460
04F3
0535
03EF
00D5
FD42
FAF6
FA5E
FA87
FA95
FA95
FAE3
FB4D
FB4B
FAE0
FAA6
FAFE
FB87
FBA2
FB49
FAFF
FB19
FB62
FB72
FB2B
FAC6
FA96
FAB0
FAE2
FAF0
FAE2
FAF5
FB3A
FB73
FB77
FB73
FBA1
FBCC
FB7E
FAF3
FB6A
FDF4
01F4
0553
0683
05F2
0522
04DB
04B9
0452
0405
0457
0508
0546
04CA
0431
0422
047F
04B4
0497
0484
04BD
0512
052E
0503
04C6
04A6
04AA
04CE
050F
055A
056C
0508
0455
03F4
0462
0533
0511
02E0
FF0A
FB76
F9E3
FA51
FB46
FB8F
FB57
FB61
FBC0
FBDA
FB7A
FB31
FB79
FBF2
FBD6
FB1C
FA97
FADD
FB87
FBC2
FB69
FB14
FB39
FB9A
FBAE
FB60
FB0A
FAED
FAE7
FAC8
FAB4
FAF1
FB5B
FB63
FAEA
FADD
FC88
0018
0400
0633
060F
04D3
0423
045E
04B0
0483
043C
0472
04F2
0507
048A
041F
044B
04CB
0505
04E2
04D7
0523
0570
055B
0508
04E5
0506
0514
04EC
04DD
0525
0570
052E
047B
0439
04FC
05E6
051E
01C0
FD25
F9D9
F936
FA4B
FB3C
FB45
FB11
FB52
FBB8
FB99
FB1A
FB07
FB8F
FBE4
FB62
FA8C
FA69
FB13
FB99
FB4A
FA89
FA30
FA68
FAA8
FAA0
FAA8
FB12
FB89
FB81
FB18
FAFA
FB62
FBA0
FB00
F9FA
FA23
FCA8
00E6
04B2
064D
05E4
0518
051E
05A8
05B3
04FD
0447
0441
04A9
04D4
04AD
04BD
052E
0576
0527
04A9
04B0
053D
05A6
0594
0572
05A5
05D7
056D
048B
040D
0461
04E1
04C3
0451
048F
059A
05FB
040C
FFF0
FBBE
F997
F9BD
FAB3
FB16
FADE
FAD4
FB3E
FB92
FB68
FB1A
FB38
FBA1
FBA7
FB14
FA89
FAAE
FB48
FB85
FB1D
FA9A
FA85
FAAE
FAA9
FA95
FAE8
FB8D
FBC9
FB40
FA97
FAB9
FB88
FBDD
FB15
FA3E
FB42
FEC8
0344
064F
06D6
05D4
0500
0507
0545
0501
047F
047D
0501
0544
04D5
0449
046B
0516
0567
0508
04B1
050F
05B0
0593
04A9
03FF
044C
04F4
0502
0489
046C
04ED
054C
04FC
0498
04FA
05AF
050B
0215
FDE9
FABF
F9C6
FA54
FB03
FB23
FAFB
FAFB
FB2B
FB47
FB32
FB1A
FB29
FB42
FB2F
FAF7
FAD6
FAE4
FAEE
FAC5
FA8F
FA9C
FAEC
FB20
FB13
FB2F
FBD3
FC7C
FC29
FACB
F9B4
FA17
FB6E
FC03
FB40
FABB
FC7D
007E
0479
0654
0624
0581
0566
056F
04FB
0455
0442
04DB
0559
051E
048C
0484
0536
05D8
05AA
04F4
04AC
0532
05D7
05B5
04D9
042D
044F
04E0
051C
04E0
04A1
0495
0479
0441
0475
054D
05CB
0465
00CD
FCAB
FA1D
F9C3
FA7B
FAEE
FAE4
FAE8
FB33
FB6E
FB54
FB1C
FB11
FB27
FB18
FAD1
FA8C
FA7B
FA90
FA9E
FAA9
FAD9
FB26
FB42
FAF6
FA8C
FA97
FB43
FBF7
FBEB
FB28
FAA1
FB07
FBC0
FBAD
FAEF
FB3D
FDF4
022F
0573
0648
058A
04F8
0512
050E
0490
0460
0519
05FB
05D7
04CB
0430
04D1
05D4
05EB
050A
045E
04AD
0569
059B
0527
04BC
04C4
04F3
04EA
04C8
04D5
04F1
04BA
043F
0426
04E1
05CC
0563
02B1
FE79
FAD8
F97D
FA47
FB8F
FBDF
FB39
FAAB
FAD6
FB4A
FB48
FACB
FA6E
FA8E
FAE2
FB02
FAF6
FB03
FB22
FB0E
FAC9
FABE
FB21
FB90
FB8C
FB31
FB0E
FB4C
FB6C
FB11
FAAB
FAE6
FB90
FBB9
FB19
FADC
FC80
FFF3
0372
0558
05AA
058C
0597
055F
049D
03FB
0445
0530
059F
0514
045A
046D
0539
05C1
0576
04D9
04AD
04FE
053B
0514
04CE
04C6
04F3
050A
04ED
04C4
04B7
04AD
0479
043E
0470
0536
05C4
04AD
013E
FCAD
F97A
F938
FAF3
FC37
FBB3
FA60
F9F6
FAC1
FB98
FB8D
FAFA
FAB0
FAD0
FAE5
FAD3
FAFA
FB6F
FBB1
FB69
FB04
FB09
FB4C
FB38
FAC5
FA90
FAF4
FB85
FBBA
FBA8
FBBD
FBD9
FB61
FA4D
F9BC
FAF6
FE05
0199
0442
0588
05D9
05D3
05BA
0586
0534
04FB
0516
0575
05B1
057D
050E
04EF
054E
05AB
056E
04BE
0456
048B
04D8
04A7
0432
041E
0484
04D5
04C1
04B0
0509
0560
0504
043B
0429
0524
05AB
03D0
FF9A
FB69
F9A3
FA5C
FB96
FB9D
FA9D
F9ED
FA44
FB13
FB6D
FB16
FA88
FA3A
FA3E
FA6C
FAA6
FAD4
FAD7
FAAD
FA92
FAD9
FB86
FC35
FC6D
FC13
FB74
FAF2
FABD
FAD1
FB16
FB5F
FB66
FAFF
FA7D
FAB9
FC88
FFE3
0394
05F9
064F
0551
046C
0467
04E1
051A
04F5
04EC
0542
059D
0596
0556
0557
05A0
05C0
0583
0541
0542
0536
04B7
0411
0403
04AB
053B
04FE
0459
043D
04BE
04F2
0454
03B7
0424
0523
04D9
021B
FDF8
FACB
F9F5
FAC0
FB7F
FB50
FAB3
FA90
FB1E
FBBF
FBC4
FB22
FA6C
FA32
FA77
FACE
FAE4
FAC4
FA9C
FA7E
FA7A
FAB5
FB33
FBA8
FBB2
FB5E
FB2D
FB70
FBD7
FBE3
FBA2
FB90
FBBB
FB9B
FB0D
FB1E
FD21
00EA
0486
0609
0575
0476
046D
0525
0594
054D
04CB
0493
0499
04A1
04B8
0504
055A
055A
0506
04D2
0508
054F
0521
0490
0442
049F
053D
055B
04D2
0437
041F
046E
0497
046D
0452
0487
0473
0306
FFEB
FC4A
F9FE
F9E6
FB10
FBC8
FB63
FAB3
FAC5
FB7F
FBE3
FB71
FAC6
FABA
FB43
FBAC
FBA3
FB81
FB8B
FB7E
FB26
FAE4
FB20
FB84
FB64
FAC9
FA8F
FB28
FBDA
FBBC
FB16
FAFE
FBA0
FBDA
FB03
FA55
FBC2
FF84
03A7
0608
0646
0586
04DA
047D
0454
046E
04D0
0525
051D
04D6
04A4
0497
0489
046E
0459
0442
0423
041F
045C
04B5
04DD
04D3
04F0
0554
0591
053A
0499
0458
048B
049F
045F
045B
04C3
047F
0248
FE89
FB64
FA7A
FB30
FBA5
FB02
FA2A
FA35
FAF7
FB75
FB4D
FB03
FB15
FB63
FB97
FBA4
FBAE
FBB5
FB99
FB65
FB50
FB6E
FB8E
FB6D
FB0F
FABB
FAB0
FAF9
FB78
FBF6
FC2D
FBE9
FB37
FA7A
FA4A
FB2D
FD3F
000F
02CD
04D1
05E5
062F
05F1
056B
04EE
04C0
04EB
0525
051A
04CC
048E
04A5
04EC
0504
04CF
0493
04A3
04E4
04EA
047D
03FC
03FD
0490
0511
04F6
0482
0464
04B8
04E9
04B6
04AB
0531
0572
03F5
0084
FCD7
FAE5
FAD5
FB2F
FAED
FA81
FAA6
FB0D
FAE3
FA34
F9E9
FA7D
FB5A
FBB3
FB76
FB2C
FB24
FB39
FB3E
FB3F
FB3C
FB1C
FAFB
FB1B
FB5D
FB51
FB06
FB34
FC18
FCB0
FBE2
FA56
FA36
FCD7
010B
0455
057F
0557
0521
0521
050B
04EF
0511
0544
052C
04F4
0515
057E
058C
0501
047D
049D
050F
0505
0475
0432
04B4
055D
0568
04FA
04B9
04C0
04AD
0484
04C5
0565
0546
0351
FFE5
FCAD
FAF9
FAA2
FAB9
FABD
FAD7
FB22
FB54
FB2F
FAE6
FAD6
FB14
FB5D
FB62
FB09
FA84
FA35
FA6E
FB15
FB9C
FB8A
FB0F
FACE
FB07
FB42
FB0B
FAC1
FB18
FBE3
FBF4
FAB8
F981
FA76
FE18
0266
04E7
0525
04B1
04F0
05AB
05E8
0576
0502
04EE
04DF
048E
0455
048A
04D9
04C2
047D
04B8
057F
0601
0598
04B1
044E
04C7
057F
05B7
0541
046A
03AE
03A5
04A3
05FD
061C
03F1
003E
FCEF
FB3E
FAD1
FAB4
FA90
FAA6
FAFC
FB2A
FB03
FAD3
FAD7
FAE3
FADD
FB0A
FB7C
FBBC
FB68
FAEC
FAF7
FB70
FB88
FAEA
FA40
FA39
FA96
FAB9
FAD0
FB80
FC72
FC4C
FAB6
F986
FAE5
FE9B
022D
03BC
03D9
0431
052D
05BA
052A
0443
0425
04D2
056C
057B
0546
051B
04E7
049B
047C
04C5
0532
0544
04DD
046E
0478
050D
05C9
061D
05A7
0490
03AA
03DF
052B
063E
058D
02DB
FF70
FCD6
FB89
FB04
FAC6
FAD1
FB30
FB91
FB8E
FB33
FAE3
FACB
FAC4
FABB
FAE3
FB48
FB8C
FB54
FAE0
FACD
FB40
FBAB
FB91
FB1B
FAC0
FAA5
FAB8
FB19
FBDA
FC64
FBC4
FA17
F91D
FA9F
FE50
01F3
03DF
0489
0540
061B
061C
04FE
03E8
03F8
04DD
056B
0531
04CA
04BB
04CB
04A8
0492
04D5
0527
0515
04B9
0486
0490
0493
0486
049C
04BA
0478
03F4
0410
0545
067A
05E6
032D
FFDC
FD82
FC16
FAD2
F9D8
F9F4
FB13
FBF3
FBAF
FAD1
FA72
FAC7
FB1E
FB1F
FB31
FB8F
FBB9
FB4B
FAC1
FAD3
FB6E
FBE1
FBD0
FB77
FB1E
FAE0
FB04
FBCE
FCBF
FC96
FACC
F8D4
F902
FBF9
FFD0
023F
030A
03A6
04ED
0618
060B
04EC
03F2
03F5
04B6
0569
0586
050B
044B
03CF
0408
04D7
0585
057A
04E3
0461
043C
043D
044D
04AE
055A
059A
04D7
03AF
038E
04E4
0641
05BA
0306
FFB1
FD43
FBDE
FADA
FA27
FA4C
FB32
FBD4
FB80
FAC6
FAB1
FB59
FBDC
FBA9
FB30
FB23
FB78
FB9A
FB4D
FAF8
FAF6
FB27
FB38
FB13
FACF
FA94
FAB9
FB78
FC48
FC18
FAB0
F983
FA57
FD1A
FFD3
0105
0187
0329
05E6
0795
06A9
0440
02CB
0354
04E1
05FD
060A
052D
03EF
0330
03B1
0528
0626
058F
0411
0368
0439
056E
05E2
05B6
057F
0515
042F
0393
0469
0649
0719
0563
0220
FF76
FE10
FCCC
FAEE
F981
F9CA
FB4B
FC4B
FBF7
FB16
FAB1
FADE
FB1C
FB31
FB43
FB5D
FB55
FB28
FB07
FB06
FB0E
FB28
FB6E
FB97
FB2C
FA67
FA4C
FB56
FC69
FBFA
FA24
F8E0
F9CE
FC5E
FEC0
0040
01D8
044A
0696
0712
0595
03C9
0353
043F
056A
05E1
058A
04CB
0422
040C
04BC
05B5
0605
054D
0444
03F2
0480
0538
0578
054E
04F8
047A
03F9
041E
0555
06C7
06C9
04C3
01FB
0004
FED7
FD39
FADB
F923
F96F
FB32
FC74
FC1A
FAE8
FA30
FA52
FAD1
FB4D
FBB5
FBDB
FB85
FAE9
FA99
FADA
FB63
FBC6
FBCF
FB6A
FA96
F9D0
FA00
FB66
FCB6
FC41
FA3A
F8E7
F9FF
FCAD
FEE4
0024
01B7
0449
0683
06B4
052C
03E6
0418
050C
0592
0588
0567
0529
0494
0413
0456
0525
0579
04DC
0414
040D
04B0
052F
053D
052D
0516
049D
03ED
03F9
052D
0675
0653
04AA
02AB
010B
FF36
FC95
F9F2
F8D8
F9BD
FB63
FC35
FBCE
FAE8
FA4C
FA47
FAC7
FB79
FBD5
FB8C
FAF5
FAB0
FAF2
FB58
FB88
FB91
FB88
FB30
FA7E
FA2D
FB13
FCB1
FD36
FB91
F919
F856
FA31
FD15
FF16
003D
01F6
04A9
06DD
0710
05A0
0448
0414
04A2
0526
056C
0586
053F
0471
03B4
03EA
0503
05D6
0584
0484
03FA
044D
04EC
053B
052F
04F4
0496
0441
0464
0523
05D1
0586
0437
02A0
0110
FEF6
FC1A
F99C
F8F9
FA34
FBB5
FC02
FB27
FA4B
FA3C
FAD8
FB89
FBD8
FB8E
FAD6
FA5A
FAB4
FB92
FBF1
FB72
FAEC
FB25
FBA5
FB79
FAC8
FAB2
FB89
FC18
FB4B
F9EF
F9D0
FB4D
FD00
FE07
FF64
0241
05AD
0761
0689
04BA
03E6
044E
04F1
0541
0583
05BD
0561
0464
03C4
0457
0581
05DC
04FD
03DB
0389
0420
04FC
058C
0594
050A
0436
03C6
044D
0579
0635
05C9
047D
02E6
00FA
FE5D
FB6D
F968
F942
FA91
FBE8
FC21
FB3F
FA32
F9E7
FA90
FB89
FBEF
FB7A
FAD2
FADF
FBA4
FC2A
FBB9
FAD8
FAAA
FB63
FC04
FBB3
FAE9
FABA
FB40
FB86
FAFF
FA5F
FA8F
FB6C
FC46
FD4C
FF83
0301
0610
06D5
058A
043D
0450
051E
0569
0524
051B
055A
050B
03FD
0354
0415
0597
0629
0531
03D5
0378
042A
0509
0575
0564
04EE
0440
03E7
0462
0561
05D9
0535
03F3
02CC
0188
FF57
FC51
F9E8
F974
FAAC
FC0A
FC5F
FBAC
FABF
FA69
FAE9
FBC0
FC0C
FB6D
FA88
FA56
FAF0
FB6C
FB25
FAA9
FAE6
FBAA
FBD0
FB03
FA5E
FAD0
FBBE
FBFB
FB87
FB60
FBC3
FBDA
FB77
FC1A
FF2C
0397
066A
0625
0460
0393
0433
04D8
04B1
0474
04D9
0551
04F8
041C
03F2
04DE
05D2
05BA
04D3
043C
047D
0523
0592
059A
054D
04BC
0421
03EC
044D
04E4
0516
04BE
0426
0359
01D9
FF44
FC2D
F9E4
F95B
FA5B
FBBF
FC63
FBF1
FAFE
FA76
FACE
FB99
FC02
FBA9
FAFF
FAB6
FAF7
FB5B
FB8E
FB98
FB82
FB23
FA95
FA68
FAF9
FBBC
FBAF
FAC9
FA37
FAD5
FBCF
FBC2
FB0B
FBE3
FF8B
0436
06B6
0609
0445
03D2
04B5
0546
04D3
045C
04BA
054E
0522
047C
0460
04EE
053A
04BD
0415
0404
045F
0478
0446
0463
04F7
0560
0527
04C0
04D9
0564
05CD
05C2
0538
03E5
016A
FE2B
FB64
FA1E
FA38
FAC4
FB1D
FB4A
FB6B
FB5B
FB13
FAEE
FB2A
FB7F
FB86
FB5A
FB58
FB89
FBA5
FB9C
FB9C
FBA2
FB69
FAF8
FAD7
FB4F
FBC9
FB78
FAA0
FA5C
FAFE
FB70
FADE
FA5E
FBF8
0000
0444
0656
0602
0507
04C2
04EF
04C5
0461
046E
04F3
0533
04CE
0444
043A
049F
04E2
04C3
048B
048B
04B9
04E2
04F5
04F0
04C3
0473
044A
0483
04EB
051A
0509
0505
04F4
03F6
0151
FDA9
FACA
F9F9
FABA
FB83
FB78
FB06
FAF1
FB42
FB79
FB62
FB48
FB66
FB8F
FB8A
FB70
FB6B
FB5F
FB21
FAD9
FAE1
FB3D
FB8E
FB92
FB74
FB77
FB7F
FB3F
FADA
FAFB
FC43
FEAF
01A7
0452
05E3
05F6
0504
0432
0450
0507
0561
0501
048B
04AA
051D
051B
0479
03F1
041C
04AE
04F9
04CA
0478
0454
046B
04B1
04FD
04F6
0475
03F4
0430
04F2
04B8
022C
FE00
FAA0
F9BB
FA9E
FB5B
FB21
FAC0
FB0F
FBAE
FBB7
FB1E
FAB4
FAFB
FB7E
FB8E
FB2B
FADF
FAF3
FB33
FB64
FB8C
FBAA
FB8F
FB37
FB0C
FB74
FC26
FC44
FB68
FA71
FAF2
FDA8
0197
04CD
0605
0591
04CC
04BB
054C
05BA
057F
04D7
0461
046F
04C2
04E6
04B6
0471
0461
0487
04B0
04B2
049A
048D
049B
04B1
04AD
047D
0440
044D
04D9
056D
04E5
0267
FE91
FB48
FA14
FAB1
FB84
FB6B
FAC2
FA81
FADA
FB25
FAFC
FACA
FB02
FB6E
FB88
FB55
FB43
FB73
FB89
FB5A
FB3D
FB82
FBD5
FBB0
FB33
FB0C
FB6C
FB9D
FB05
FA4A
FAE0
FD74
0123
043C
05AA
058E
04DB
0474
049D
04FB
050A
04AE
045B
0481
04FA
0527
04C1
043A
042C
049D
050F
051A
04C4
0457
041A
0434
0490
04D9
04CA
0498
04C8
0552
052A
0326
FF83
FC12
FA7C
FAB3
FB51
FB55
FAF9
FAE8
FB38
FB73
FB62
FB4A
FB69
FB98
FB9A
FB7B
FB68
FB61
FB4F
FB4B
FB7A
FBAC
FB77
FAD3
FA59
FAA1
FB77
FBF3
FB7F
FAAA
FACD
FCCC
0037
0390
056B
057D
04AF
0436
0483
0513
052F
04C5
0457
0448
046F
0478
046F
049A
04EB
04F6
048A
0411
0419
049E
0514
0519
04D0
048F
0476
0491
04FF
0592
055F
0358
FFA4
FC05
FA56
FABE
FBB8
FBD8
FB32
FACA
FB17
FB95
FBA7
FB60
FB35
FB53
FB8A
FBAF
FBB4
FB83
FB15
FAB8
FACF
FB49
FB92
FB4C
FADC
FAF3
FB8C
FBD2
FB35
FA55
FA93
FCBD
0040
039A
056E
0573
0490
040A
045E
04F2
04F2
0462
0410
0475
0509
0509
048F
0466
04D0
0521
04D0
0459
0480
051F
054E
04C0
0433
0462
04FE
0541
051E
0513
04E9
0376
0034
FC70
FA3B
FA36
FB21
FB8D
FB5B
FB51
FBB6
FBF8
FBA6
FB1D
FB04
FB6F
FBD1
FBB6
FB2F
FAA3
FA75
FACE
FB72
FBCF
FB7B
FAC0
FA74
FB0E
FBF6
FC06
FADB
F98B
F9CC
FC61
0058
03D0
0569
0537
0470
043D
04BC
0529
04EB
044E
0418
0487
0504
04EF
046E
0431
047C
04E0
04ED
04C9
04DB
0513
050A
04B9
0499
04E8
0531
04F0
0475
0476
04BE
03F0
011D
FD45
FAA1
FA57
FB6C
FC18
FBC9
FB48
FB4B
FB86
FB62
FAF8
FADB
FB2A
FB69
FB42
FB04
FB1E
FB77
FB9B
FB60
FB17
FB06
FB18
FB28
FB51
FBA7
FBD9
FB83
FAE5
FAFF
FCA4
FF92
028A
0466
04EA
04AC
0457
0429
041A
042B
0477
04EE
0540
051E
04A0
0443
0469
04E7
0534
050D
04B4
048D
04A0
04B6
04BB
04C9
04CA
0478
03EA
03D0
049B
056E
0486
0126
FCD3
FA24
FA33
FBA7
FC66
FBD5
FB09
FB07
FB8B
FBB3
FB5C
FB2C
FB74
FBB3
FB63
FAD8
FAD1
FB5F
FBC5
FB7D
FAF3
FAE8
FB64
FBBB
FB90
FB44
FB46
FB5F
FB26
FB04
FC1F
FEFA
028E
0513
05B2
051A
0479
0453
0471
0493
04C4
0500
0506
04AE
0448
0445
04A2
04E2
04B2
0458
0453
04B2
0502
04DF
0478
0443
045E
0479
0462
046A
04DE
0535
0437
014A
FD7D
FADA
FA70
FB53
FBC3
FB2A
FA7A
FAAD
FB6C
FBAC
FB2D
FAC6
FB22
FBD1
FBEE
FB6C
FB0F
FB4A
FBA7
FB97
FB4C
FB58
FBB6
FBCD
FB6F
FB2C
FB6F
FBB5
FB49
FAA6
FB61
FE5C
0269
0546
05D3
04F6
044D
047C
04F8
0523
0506
04FB
0509
04EF
04A1
046B
0479
049B
048F
0467
046C
04AC
04DE
04C0
047D
046F
04A3
04C6
04A7
0492
04D8
050B
0415
0159
FDB1
FAE3
FA0C
FAAB
FB67
FB84
FB4F
FB40
FB3D
FAFE
FAB4
FAE2
FB80
FBDD
FB82
FAED
FAEF
FB92
FC02
FBB5
FB1F
FAFC
FB45
FB5F
FB20
FB16
FB8F
FBEC
FB71
FAA9
FB3A
FE17
022D
053D
0607
053D
0468
0456
04B6
04F3
04EE
04DD
04DB
04D6
04CD
04D5
04E8
04D8
049D
0477
04A3
04F3
04F4
0488
0424
044C
04D7
0505
047F
03E9
0425
04EE
04BE
025B
FE6E
FB22
FA0B
FABF
FB99
FB9B
FB20
FAEA
FB0F
FB2A
FB1F
FB2E
FB5D
FB4F
FAE5
FA92
FACA
FB47
FB5D
FAF7
FAC5
FB3A
FBCF
FBB8
FB18
FAE3
FB82
FC1E
FBBE
FAD9
FB2B
FDC7
01B5
04C7
05BA
052D
0490
049B
04ED
04F2
04A9
047B
049A
04CC
04D4
04C6
04D6
0502
0515
0502
04F9
051B
0535
0502
049D
0474
04B4
04F3
04C1
0465
048C
0528
04F4
02B2
FEC9
FB40
F9D7
FA60
FB45
FB68
FB0E
FAFB
FB44
FB67
FB37
FB18
FB41
FB5B
FB10
FAA7
FAB2
FB2E
FB77
FB2F
FACD
FAF1
FB78
FBAE
FB54
FAFB
FB25
FB73
FB29
FA7C
FAC8
FD2F
011C
048E
05EE
056F
048B
0464
04E2
053D
0516
04C9
04CD
0517
0541
0517
04D0
04B5
04CA
04E6
04F1
04F0
04DC
04A7
0472
0486
04E9
052A
04E3
0460
0464
0502
050F
0331
FF89
FBEB
FA30
FA70
FB3E
FB67
FB0E
FAF5
FB3B
FB51
FAF4
FA9F
FAD3
FB4C
FB60
FAF0
FA91
FAC1
FB3F
FB82
FB6E
FB55
FB4F
FB1C
FAB3
FA91
FB0C
FBA4
FB7D
FAB5
FAB7
FCDE
00C2
0457
05DD
056C
0486
045D
04D6
0531
0521
04F4
04F3
04F9
04D2
04A4
04B9
0505
052A
04FC
04BA
04B2
04D1
04D2
04BD
04E2
054B
057A
0510
047A
048E
054C
0561
0367
FF98
FBE8
FA30
FA74
FB32
FB3B
FAC3
FAA6
FB13
FB6C
FB42
FAF4
FB10
FB82
FBBA
FB7F
FB2E
FB1F
FB26
FAF5
FAB2
FAC6
FB2C
FB5E
FB1A
FAD3
FB0F
FB7D
FB46
FA6D
FA56
FC6C
0062
042E
05FC
05D4
0520
04F1
051E
050B
04B6
0499
04D9
0504
04C5
0467
0469
04C2
04F5
04CD
04AB
04EA
054B
0547
04E1
04B4
0514
057C
0538
047F
044E
04FB
055B
03C8
001B
FC28
FA0C
FA32
FB36
FB9B
FB2C
FAA9
FA9D
FADE
FB15
FB34
FB4E
FB4E
FB1B
FAE7
FB01
FB55
FB77
FB31
FAD6
FACB
FAF8
FAFB
FAD2
FAF7
FB94
FC0B
FB9D
FA93
FA5B
FC2F
FFB9
0340
0537
0572
04F5
04C6
0515
056E
056C
0523
04EB
04EB
04FD
04EF
04C7
04AB
04B0
04C2
04D0
04E3
0502
0516
050C
0500
0515
0524
04E4
0479
047A
0518
0565
03F5
0082
FC99
FA47
FA1F
FAE9
FB3E
FAFA
FADF
FB40
FB9D
FB6F
FAE0
FA7F
FA8E
FAE3
FB42
FB87
FB85
FB25
FAAB
FA91
FAF0
FB4F
FB4D
FB23
FB2C
FB43
FB0F
FAFB
FC33
FF46
030C
0589
05EB
0533
04C9
04FA
0523
04EC
04AF
04C2
04F8
04FB
04CE
04B0
04B2
04B4
04B9
04DE
0507
04F5
04BB
04BD
0503
0511
04B6
0486
04FA
0543
03CD
003E
FC5B
FA64
FAAE
FB85
FB60
FA84
FA21
FA94
FB27
FB44
FB21
FB2E
FB65
FB7C
FB68
FB54
FB4A
FB2F
FB10
FB11
FB16
FAF1
FADA
FB41
FBE7
FBDB
FAE4
FA79
FC62
0068
0421
0570
04B9
040B
047F
054A
0562
0501
04F5
053E
0531
04B3
046D
04B7
050A
04DC
0478
0484
04F9
0531
04F6
04B7
04AB
0473
0407
0423
050B
056B
0378
FF55
FB78
FA22
FAFF
FBE8
FB9C
FADE
FAD5
FB61
FB94
FB35
FAD8
FADC
FAFC
FAF5
FAF2
FB16
FB27
FAFE
FAF2
FB56
FBCC
FBB9
FB3F
FB24
FB88
FB8E
FAE2
FAD7
FD08
010D
0483
0597
04E6
045A
04BA
0531
04F4
0471
046A
04C9
04F9
04E8
04FE
0541
0540
04E4
04AB
04D4
04F0
0491
041C
043C
04BF
04D2
0462
045A
050B
0517
02EA
FEF9
FB92
FA63
FAD6
FB49
FB23
FB05
FB4C
FB6F
FB0B
FAA7
FAE2
FB66
FB6C
FAF4
FABB
FB16
FB80
FB7D
FB4C
FB58
FB7A
FB4D
FB0F
FB51
FBDD
FBB7
FAC8
FAAB
FCFD
0125
04AA
05D1
0537
049F
04CC
0529
0525
0500
0516
0534
0507
04BE
04B2
04C3
049B
0459
0471
04D6
04EE
0480
042F
048A
0517
04F9
045D
045A
051B
050D
02A6
FE94
FB47
FA4D
FAED
FB79
FB4B
FAF5
FAEA
FAE3
FAA6
FA8F
FAF1
FB74
FB94
FB65
FB55
FB66
FB40
FAE9
FAE1
FB4E
FB96
FB42
FAD2
FB0C
FBB1
FBB2
FB00
FB33
FDB7
01C5
04F1
05C3
0507
046E
0495
04E6
04E6
04D1
04ED
04F8
04B2
0468
0481
04D8
04F7
04D3
04C1
04D2
04C4
0494
04A9
0518
0546
04C2
0433
0492
056D
04DA
01B7
FD6E
FAA3
FA5B
FB35
FB79
FB06
FADB
FB4C
FBA2
FB5E
FAF5
FB03
FB59
FB67
FB2B
FB0B
FB1B
FB12
FAEE
FB0D
FB7B
FBAB
FB4C
FAE7
FB25
FBA8
FB83
FADF
FB5A
FE19
020C
04E5
0593
0511
04CC
04F9
04F2
0492
046F
04CA
0525
050D
04C2
04B3
04CA
04BB
04A4
04D1
0512
04EC
047C
0472
04FF
0557
04D4
042A
0480
0564
04BE
0163
FCF6
FA55
FA71
FB98
FBDA
FB2C
FABC
FAFE
FB3D
FAFB
FAAF
FAE6
FB58
FB74
FB4A
FB55
FB9C
FBAA
FB59
FB0C
FB03
FB06
FAEF
FB09
FB7C
FBAA
FB01
FA4F
FB65
FEDC
02F1
0540
0551
04AE
04B2
0524
052E
04D3
04C3
0520
0542
04D5
0461
0471
04C0
04CE
04AC
04BB
04DD
04AA
044E
0474
0522
0571
04D7
0431
049A
056A
0485
010D
FCDF
FA8F
FA8D
FB22
FAF8
FA90
FAE5
FBAE
FBD4
FB2C
FAB1
FAFF
FB78
FB5B
FAF2
FAF9
FB60
FB75
FB15
FAEB
FB51
FBBF
FB9E
FB29
FAF6
FAF3
FAAD
FA97
FC0A
FF7D
0364
0599
05A0
04D9
049E
04ED
0516
04E8
04C2
04C7
04BB
049C
04C1
0529
054A
04E4
047F
04A1
04FC
04EF
0492
048C
04EF
0503
0483
0452
0521
05CD
0438
0010
FBBD
F9E0
FA81
FB81
FB6C
FAD5
FAD8
FB5E
FB83
FB1F
FAE8
FB30
FB5D
FAFB
FA8E
FAC7
FB68
FBA5
FB4E
FAF2
FAEA
FAF4
FADE
FAF2
FB53
FB75
FAF8
FACE
FC8E
004E
040B
05B0
0552
04AA
04C5
0517
04DE
046D
048E
0531
057F
0523
04B8
04C2
04EB
04BC
0471
0495
050E
0541
050D
04EB
0511
050F
04A5
045F
04B1
04C6
031A
FF86
FBED
FA4E
FAA5
FB5B
FB5C
FB05
FB01
FB2F
FB10
FAC3
FADD
FB63
FBAD
FB5D
FAE2
FABD
FAD5
FAD7
FAE4
FB3A
FB93
FB77
FB1A
FB2A
FBAB
FBB5
FAE4
FA96
FCA2
00D8
04AF
05F4
051C
044D
04A2
0553
055B
04EE
04DA
052C
053F
04E5
04AF
04F8
0550
0539
04E4
04C7
04D8
04BF
048A
0490
04B9
049A
044D
048C
056C
0582
033E
FF10
FB6C
FA35
FAD8
FB70
FB26
FAB5
FAD4
FB28
FB0B
FAA0
FA88
FADE
FB1E
FB0A
FAF8
FB1C
FB27
FAEA
FAD2
FB39
FBAF
FB8D
FB02
FADB
FB38
FB4C
FACA
FAED
FD34
013D
04BC
05EE
055A
04B9
04CE
050A
04ED
04C4
04F2
0540
0547
0526
0536
0556
0515
0489
045B
04C1
0516
04D9
047A
049E
0506
04FB
04A0
04DD
05B2
057C
02BA
FE45
FACE
F9F9
FACC
FB50
FAF6
FAA2
FAE7
FB46
FB2A
FAC9
FAAA
FACD
FADA
FADA
FB20
FB90
FBA3
FB3B
FAE5
FAF8
FB13
FAD9
FAB5
FB23
FB9D
FB36
FA4B
FABF
FDD3
023F
054F
05C7
04EB
048C
04EE
0536
0512
0500
053C
0556
0502
04A5
04A7
04C8
049C
0467
04B9
055E
0570
04C2
0451
04D6
059C
0588
04D6
04BD
0549
04BF
01BD
FD69
FA78
FA27
FB1C
FB73
FAF3
FAA0
FAE6
FB2F
FB10
FAEB
FB2D
FB99
FBB2
FB77
FB38
FB05
FABD
FA9A
FB00
FBA3
FBAA
FAE4
FA49
FAA2
FB51
FB3F
FAC7
FBAA
FEC9
02B2
051C
0573
0515
052E
056F
0521
048E
047E
04E2
04F2
0483
0455
04DC
0578
055F
04CA
0490
04D4
04F1
04AC
04A0
0516
0550
04B4
0405
046B
0563
04D1
018E
FD26
FA57
FA18
FAF5
FB41
FAEC
FAD5
FB33
FB7C
FB6E
FB53
FB4E
FB1C
FAB5
FA89
FAD6
FB29
FB06
FAC2
FB05
FBAA
FBD0
FB47
FAF4
FB6B
FBD3
FB2E
FA4B
FB51
FF02
0364
05C8
05A4
04B9
0493
04F7
04FC
04AB
04B9
052C
0554
04F0
049A
04CF
053C
054E
0509
04DB
04CB
048D
043A
045B
04F1
053B
04DD
0494
0516
0587
041F
0079
FC7B
FA6F
FA9F
FB6E
FB81
FB06
FAC2
FACB
FABE
FAA4
FADA
FB48
FB65
FB11
FAC9
FAEB
FB32
FB49
FB64
FBCD
FC16
FB91
FA88
FA33
FB01
FBC1
FB44
FA6E
FB83
FF46
03AD
05FE
05BE
04C1
04AD
0548
057C
0517
04C7
04DE
04F8
04CB
04A4
04D4
051E
0515
04BF
047E
047A
0482
0488
04B9
0506
050F
04D1
04D9
055E
0564
0394
FFF8
FC59
FA7E
FA73
FADB
FABF
FA71
FA9A
FB24
FB7A
FB6D
FB4F
FB4B
FB36
FB01
FAEE
FB29
FB6F
FB6A
FB30
FB14
FB23
FB20
FB17
FB5A
FBD7
FBE1
FB31
FAC9
FC2F
FFA3
0386
05D9
061B
0568
04FC
050F
0526
04FB
04B9
049B
04A7
04D0
04FB
04FD
04C6
048D
049C
04E8
050B
04D8
049F
04B3
04DC
04B0
0465
04AB
0572
0555
02F7
FEDF
FB53
FA1C
FACE
FB8C
FB44
FA8B
FA6D
FAFD
FB72
FB5A
FB0E
FB04
FB2F
FB3B
FB1A
FB0C
FB2C
FB44
FB27
FAFE
FB15
FB65
FB80
FB17
FA8F
FAF0
FD0F
009A
0411
05E0
05C4
04EB
04AD
0538
05AF
0564
04A9
0445
0476
04C9
04E1
04DF
04FC
050B
04CD
0477
0485
04F5
052D
04D3
0476
04DC
05B8
0586
031A
FF1A
FB99
FA23
FA71
FB12
FB19
FAC8
FAC9
FB28
FB5E
FB28
FAE7
FB07
FB5E
FB6A
FB17
FAE8
FB36
FB9B
FB74
FAD6
FA99
FB2F
FBD4
FB6C
FA2E
F9ED
FC3F
0093
0483
0623
05AE
04D7
04C5
052C
0544
04F5
04CC
04FD
0518
04BB
043B
0431
04A6
0501
04DF
049F
04D6
055F
056C
04AF
03FC
0461
0593
05C5
0371
FF35
FB7B
FA29
FAD4
FB8B
FB1E
FA32
FA0E
FAE2
FBAB
FBA1
FB20
FAFA
FB4D
FB81
FB44
FB02
FB2B
FB72
FB41
FAB6
FAA2
FB57
FC00
FB9A
FA84
FA84
FCED
00FD
046A
05A0
0519
047D
04C1
056D
059A
0527
04B5
04B1
04D9
04C2
0481
0486
04E7
052F
0500
049D
048F
04DA
04EA
0477
0415
0487
0573
0549
02D6
FECE
FB63
FA35
FADC
FBA6
FB82
FAD9
FA96
FAE6
FB32
FB1D
FAF1
FB0E
FB45
FB2E
FAD9
FAC9
FB2B
FB89
FB70
FB28
FB51
FBDB
FBE7
FAF7
F9FC
FAB0
FDC4
01E5
04E5
05B2
0512
0484
04AF
051C
0521
04C2
048B
04C9
052E
0547
0509
04CE
04CC
04D7
04B3
0483
0494
04DC
04E5
047D
042E
04A0
0572
0524
0297
FE85
FB1A
F9E4
FA71
FB20
FB04
FA9E
FAC2
FB5B
FBA5
FB53
FAE7
FAED
FB3A
FB46
FAFE
FAE0
FB34
FB9D
FB99
FB43
FB30
FB8C
FBC0
FB40
FA8B
FB0B
FDA2
0186
04BA
05DF
0558
04AA
04CC
0563
0592
052C
04C3
04C0
04DC
04A7
0448
0444
04B0
0503
04E3
04AB
04D9
0530
04FB
042F
03C7
0484
0597
0520
0237
FE20
FB25
FA60
FAF6
FB5F
FB0A
FA8A
FA84
FADB
FB0F
FAF9
FAF2
FB3A
FB9B
FBB1
FB72
FB34
FB2B
FB2A
FAFA
FAD3
FB20
FBCA
FC06
FB49
FA57
FAE5
FDD9
020A
052B
05FB
0546
04B2
04E5
053A
050F
04B6
04D4
054C
055D
04BF
041B
0429
04B9
0503
04BF
047F
04C4
0528
04E6
040B
03A8
047B
05AB
0552
026E
FE20
FAC2
F9C1
FA7A
FB3C
FB20
FAAE
FAC4
FB59
FBA2
FB36
FAA5
FAB0
FB4A
FBB0
FB76
FB0B
FB0A
FB5C
FB76
FB3C
FB34
FBA2
FBF4
FB7F
FABE
FB40
FDFA
01F8
050F
05F1
0540
0491
04B0
0526
053D
04F4
04CE
04FE
052F
0513
04D9
04D3
04EB
04C0
044E
0417
0478
0506
04FD
0456
0409
04C4
05AF
04E6
0193
FD30
FA47
F9F7
FB01
FB76
FADE
FA58
FAC2
FB8D
FB94
FAC3
FA28
FA7F
FB3C
FB62
FAE9
FAB4
FB3E
FBE4
FBD4
FB4B
FB3B
FBD5
FC15
FB39
FA32
FB06
FE87
0312
0608
0655
0535
048D
04F2
0586
056B
04D5
048C
04D4
0535
0538
0501
04FA
0533
0553
0525
04E1
04C8
04B7
045F
03EA
03FA
04C7
056A
0477
0174
FD9E
FADC
FA0E
FA77
FAD8
FAC1
FAA8
FAE5
FB2E
FB1A
FACF
FACA
FB16
FB2F
FACC
FA68
FAA9
FB68
FBBF
FB36
FA81
FAA3
FB8E
FC0F
FB63
FA7C
FB42
FE77
02B0
0592
060F
051D
046C
04A8
053C
0569
052E
0507
0521
052B
04EC
04A3
04AD
04FA
0527
050E
04FF
0535
0566
051D
0481
0455
04F5
057F
0471
0146
FD48
FA89
F9FD
FAC6
FB54
FB02
FA6B
FA62
FAE8
FB53
FB3B
FAEB
FADD
FB13
FB31
FB10
FAEF
FB01
FB0F
FAD8
FA97
FACC
FB6E
FBB7
FB25
FA8B
FB8F
FED3
02E9
058A
05D4
04F4
0496
0514
0585
0543
04C3
04C2
052C
054C
04E5
048E
04CE
0548
0541
04B1
0460
04C9
0558
052D
046A
042B
0505
05DD
04D2
0152
FCFC
FA30
F9D9
FADA
FB86
FB54
FAED
FAF4
FB37
FB32
FAE6
FACE
FB16
FB4C
FB14
FABE
FADF
FB6B
FBA6
FB30
FAA6
FADD
FBA2
FBD4
FAEE
FA1C
FB3A
FEB7
02DE
0570
05C1
0506
04B9
051B
056D
052B
04A8
0477
04A8
04DA
04D7
04D0
04F1
0517
0504
04D1
04D0
050F
052C
04D5
045B
046B
051E
0577
0425
00EF
FD2D
FAB6
FA3A
FAD1
FB24
FACF
FA77
FAB9
FB54
FB97
FB54
FB07
FB1A
FB51
FB39
FAE3
FACD
FB1B
FB51
FB0E
FAB3
FAE5
FB88
FBB3
FB05
FA93
FBFF
FF8B
037A
05B1
05B4
04D8
048D
04FE
055B
0522
04A9
047F
04AB
04C9
04AC
0499
04D3
0536
055E
052A
04DC
04C1
04CA
04AF
0478
0493
052B
0570
0411
00AC
FCA5
FA21
F9FE
FB0C
FB7E
FAE9
FA60
FAC4
FB97
FBCC
FB47
FAE5
FB27
FB82
FB41
FAA8
FA8F
FB20
FB91
FB51
FAE9
FB26
FBC7
FBBD
FAC9
FA4D
FBF0
FFB0
03A2
05CA
05DE
0520
04CC
0508
053E
0514
04C4
04AA
04C9
04D7
04B4
0495
04B7
0501
051A
04E7
04AD
04AB
04BB
0495
0461
04A6
0567
0592
03D4
002C
FC4D
FA28
FA1E
FAF2
FB4F
FB10
FAE2
FB1F
FB68
FB53
FB09
FAF8
FB28
FB3B
FB04
FAD4
FB0A
FB86
FBC9
FB9D
FB53
FB4D
FB65
FB16
FA69
FA6A
FC4D
0002
03DA
05EE
05D4
04D6
046F
04CF
051D
04D9
0477
0494
0503
051E
04C7
0498
04F9
0570
053D
046B
03D8
0419
04BF
04FD
04C8
04D2
055B
0570
03BC
0025
FC43
FA0F
FA1D
FB3C
FBD8
FB7D
FAEA
FADF
FB3C
FB68
FB37
FB0C
FB28
FB3F
FAFE
FAB0
FAE4
FB86
FBCF
FB58
FAC8
FAFC
FBBC
FBE8
FB1B
FAA8
FC4D
0014
03F4
05D1
0586
04A2
047A
04F2
052E
04DF
0486
049E
04F8
050F
04C9
0492
04C3
0524
0543
0507
04D1
04E5
0502
04BF
0443
043D
04DD
050F
035E
FFB4
FBE5
FA05
FA5D
FB5D
FB86
FAF1
FAB4
FB30
FBA6
FB6F
FAF2
FAF9
FB79
FB9F
FB0C
FA71
FA9C
FB54
FBA0
FB1C
FA87
FAC0
FB84
FBC5
FB31
FB00
FCBF
006B
042E
060F
05D3
04EC
04B4
051A
0531
04A9
0437
047D
051C
0542
04D0
0481
04D1
0547
052B
049B
0468
04DA
0539
04D9
043A
0464
0549
055A
0329
FF2E
FB8A
F9F4
FA43
FB05
FB37
FB05
FB0B
FB57
FB73
FB24
FAC5
FACB
FB25
FB53
FB18
FAD1
FAFC
FB80
FBC6
FB7F
FB1A
FB22
FB74
FB6A
FAF3
FB1D
FD1A
00B3
0426
05CC
05A5
0505
04F5
0542
0531
04B1
0466
04B9
0540
054F
04DC
0481
049B
04D5
04BA
046F
0486
0515
0575
051D
0487
04A4
055E
0522
028A
FE4B
FADB
F9F4
FAE8
FBB8
FB76
FAEA
FB05
FB76
FB5E
FAC3
FA8B
FB10
FB96
FB71
FB0B
FB23
FB8B
FB6E
FABE
FA7A
FB26
FBD0
FB63
FA96
FB85
FF0B
035E
05E4
05EF
0501
04A3
04E2
0507
04EC
04F8
0536
0532
04CE
0487
04AA
04CF
048D
0441
0489
0529
053E
0495
0436
04F5
05EA
0513
01AF
FD69
FABC
FA75
FB3D
FB77
FAEE
FA7D
FAA4
FB04
FB23
FB17
FB31
FB5E
FB47
FAFB
FAF2
FB51
FB92
FB40
FAC1
FADA
FB74
FB94
FADD
FA9E
FC9D
00C5
04B7
062A
0550
044B
048C
0572
05AC
051E
04B2
04D1
04F0
049F
044D
0486
04FD
0504
04B2
04C1
0548
056B
04B4
040C
0472
0529
0428
00AB
FC84
FA41
FA6A
FB4D
FB55
FAB5
FA79
FAD8
FB25
FB0D
FAFF
FB45
FB7F
FB55
FB1B
FB47
FB8D
FB42
FA89
FA68
FB47
FC11
FB93
FA77
FAEF
FE20
0285
056B
05CA
04F9
04B5
0531
0575
0516
04B0
04D0
051E
0509
04B1
04A9
04FA
0514
04C1
048F
04E9
0547
04E1
040D
040D
0527
05A5
0389
FF24
FB21
F9B8
FA78
FB43
FAFF
FA78
FAB0
FB54
FB6B
FAE7
FAA9
FB12
FB74
FB33
FAB9
FAC1
FB23
FB22
FABA
FAC3
FB85
FBFC
FB45
FA62
FB7E
FF3A
0389
05D4
05B4
04E7
04E2
0555
0549
04C3
0499
050B
056B
0537
04D5
04D9
0517
050A
04CD
04F4
0572
0579
04B5
0411
048E
058A
0508
01FD
FDC5
FAD1
FA27
FAC1
FB2A
FB11
FAFB
FB18
FB0E
FAC0
FA9D
FAE9
FB42
FB30
FAE4
FAE9
FB3C
FB41
FAC6
FA7A
FAFB
FBC4
FBB2
FAC0
FA90
FCB7
00C1
046A
05E7
057B
04B7
049C
04ED
051D
0526
0547
0564
0533
04CA
04A0
04D9
050A
04DF
04A6
04D3
0534
0523
0496
0462
0505
0582
0425
0094
FC97
FA66
FA74
FB4B
FB76
FAF4
FAA7
FAE6
FB31
FB1A
FADF
FAE5
FB1D
FB39
FB39
FB5C
FB88
FB60
FAF0
FACF
FB39
FB80
FAEA
FA21
FAEB
FE23
025C
0525
058C
04D1
049C
0520
056C
050B
048F
048D
04CB
04C8
0496
04A5
04E9
04E1
0482
046E
04FB
057B
0529
0475
0497
05A8
05E3
0389
FF2D
FB6B
FA2C
FAD4
FB71
FB1D
FA90
FA9C
FB06
FB26
FB08
FB3A
FBC1
FBF3
FB80
FAF6
FAF5
FB3A
FB19
FA9F
FA96
FB34
FB8E
FAEA
FA3D
FB77
FF24
0361
05B6
059E
04B3
048C
051D
0566
0516
04C4
04D2
04E1
0492
0439
045C
04D3
0503
04D5
04D3
053A
0573
0502
0480
04DA
05AB
0520
0219
FDD1
FAD0
FA3E
FAF2
FB34
FAB9
FA72
FAE1
FB77
FB92
FB5C
FB4D
FB57
FB24
FADC
FAFF
FB7A
FB92
FAF7
FA6D
FAC1
FB7D
FB64
FA69
FA4A
FCA6
00CF
0452
058B
0520
04C1
0515
0572
0543
04D6
04B4
04CA
04B8
0493
04BD
0522
052F
04BA
0462
04B6
054E
0552
04CF
04C2
0592
05FF
044D
0074
FC7D
FA7A
FA84
FB1A
FB1A
FAC4
FAC4
FB0E
FB19
FADF
FAF0
FB75
FBCA
FB61
FAAB
FA8A
FB11
FB6E
FB2A
FAD3
FB0A
FB59
FADF
FA06
FAA7
FDE9
026D
0577
05D1
04DB
048A
0525
058B
0528
04B3
04DB
052F
04E9
0446
043E
04FE
0592
0543
04A3
0498
04F9
04EE
0475
0496
0597
05DD
038C
FF11
FB21
F9E3
FAC3
FB93
FB3E
FA92
FA98
FB1E
FB4E
FB0E
FAFC
FB56
FB95
FB52
FAED
FAF4
FB45
FB57
FB2B
FB45
FBA8
FB90
FAAA
FA21
FBAE
FF80
0398
05B5
0586
04A4
047E
04FB
053A
04F9
04C4
04F0
051F
04ED
0497
0496
04DE
04F6
04BD
049D
04CE
04EC
04A1
0467
04E7
05A5
04F5
01DD
FD9B
FAA8
FA38
FB29
FBA0
FB24
FAA4
FACF
FB3D
FB46
FB0A
FB0F
FB53
FB5F
FB1F
FB0C
FB59
FB87
FB2D
FABF
FAED
FB73
FB52
FA7B
FA7F
FCE7
011D
04BA
05F5
054E
0487
0499
0516
0547
0521
04F3
04C4
0480
0463
04B3
052D
0538
04C4
047C
04D6
0553
0533
049C
048B
054F
05A6
03EC
0019
FC19
F9FD
FA1C
FB22
FBA8
FB62
FAE0
FAA7
FAC5
FB12
FB6B
FB9F
FB77
FB01
FAA8
FAC4
FB1F
FB3D
FB09
FAFE
FB62
FBB1
FB43
FA90
FB3A
FE4C
02A8
05CA
0642
050F
043D
04A5
056A
0588
0515
04C9
04D5
04CF
0496
0490
04ED
0541
052A
04EE
04F9
0512
04B4
0421
0442
052A
0545
02EE
FEA8
FB00
F9E2
FAB3
FB6F
FB22
FA8A
FA8D
FAF9
FB23
FB07
FB22
FB7E
FB97
FB43
FB04
FB34
FB66
FB20
FACB
FB22
FBEA
FBFE
FB06
FA78
FC30
0017
03F5
05BE
0586
04E5
04E9
0540
0549
0511
04FF
050B
04DA
0474
0456
04A9
04EE
04BA
0461
047F
04F6
0500
0466
0406
04A4
057C
04B3
017B
FD4A
FA87
FA20
FAE8
FB40
FAD5
FA79
FAB2
FB22
FB43
FB30
FB4B
FB8D
FB91
FB4E
FB2F
FB65
FB91
FB5C
FB18
FB4B
FBB8
FB8C
FAC2
FAC1
FCFE
010C
04AB
0601
0564
04A1
04D4
0579
0594
0513
04A7
04AD
04D0
04B5
0486
048F
04BB
04C3
04AD
04BB
04E2
04C8
0474
0484
053C
059D
0412
0059
FC42
FA14
FA4B
FB55
FB87
FAD0
FA4C
FA94
FB25
FB4F
FB23
FB21
FB5D
FB76
FB44
FB15
FB1E
FB2A
FB14
FB21
FB80
FBAD
FB13
FA4E
FB1A
FE6A
02D6
05B5
05DE
04B9
0457
0518
05BE
0574
04D1
04BB
050E
0503
0487
0450
04B3
051A
04FA
04AE
04D3
052E
0505
046A
0459
0515
052F
02F9
FED6
FB3C
FA1B
FAE8
FBA5
FB59
FAC1
FAC2
FB27
FB3D
FAFF
FAFF
FB56
FB7C
FB32
FAFB
FB40
FB92
FB4B
FAB5
FAC1
FB93
FC14
FB7D
FAD2
FC06
FF8D
0382
0591
0558
046E
044A
04DF
0545
0524
04E9
04EC
0502
04F2
04D9
04DC
04D1
0491
0462
04A8
0524
051A
046A
0404
04B6
05B3
0506
01C9
FD7F
FAB9
FA7B
FB70
FBC1
FB18
FA81
FAB1
FB38
FB57
FB14
FAFA
FB31
FB58
FB3B
FB25
FB50
FB77
FB4D
FB1A
FB4A
FB94
FB32
FA41
FA52
FCD7
012D
04DB
0604
0537
0469
04A0
052F
0528
04AB
0474
04AA
04D4
04BE
04C0
0502
0518
04B8
0455
0489
0513
051C
0496
0485
056C
0602
0459
004F
FC1C
FA1A
FA70
FB5B
FB7D
FB16
FB0B
FB73
FBAE
FB78
FB36
FB37
FB49
FB30
FB1D
FB4B
FB76
FB30
FAAB
FA9D
FB32
FB94
FB02
FA39
FB07
FE39
0263
052B
05A0
04E1
0485
04DB
0516
04C4
046B
049F
0513
0514
0498
044B
0489
04E3
04E0
04BF
04FB
0560
0545
04B4
0497
0547
0570
0353
FF25
FB50
F9EB
FA9C
FB76
FB6A
FB0A
FB17
FB52
FB2A
FAD9
FB00
FB7D
FB83
FAFB
FAC2
FB49
FBBF
FB54
FA9F
FAC0
FB7D
FB65
FA29
F9BB
FC22
00B0
0477
058C
04D7
0451
0497
04F0
04FB
0513
0552
053F
04BE
0475
04D5
054A
0511
047B
0478
050A
0526
047B
042A
04F5
058E
03E7
FFF4
FC08
FA44
FA80
FB24
FB47
FB36
FB3F
FB1A
FAAE
FA86
FAF1
FB62
FB47
FAF4
FB06
FB54
FB45
FAF6
FB18
FBAB
FBB8
FAEC
FAAC
FCB0
009E
041C
0574
0541
050D
0536
051F
04B2
049A
050D
056B
0534
04C7
04AD
04C8
04B2
0499
04E9
054E
0502
0446
0458
0567
0587
02E6
FE6E
FB0A
FA5F
FB37
FB86
FAF0
FA98
FB05
FB71
FB36
FACE
FADF
FB30
FB3B
FB23
FB4C
FB7F
FB4B
FAF5
FB25
FBA4
FB75
FA8F
FAA7
FD59
01CB
052E
05DA
04EB
046B
04DD
054D
0526
04D1
04C1
04D4
04D4
04E0
0510
0525
04F1
04C3
04E8
0508
04AB
0440
04A7
057F
04EA
01CC
FD97
FAE3
FA9B
FB62
FB9C
FB28
FACF
FAE0
FB01
FB0C
FB41
FB8F
FB7D
FAFD
FAA7
FAD2
FB09
FAF6
FB00
FB77
FBB0
FB01
FA50
FB8A
FF30
0344
054E
0508
043F
0450
04D5
04F3
04D4
0504
054E
051C
0498
0478
04D6
0518
04FA
04E5
050E
04F9
046E
043D
051B
05E5
0469
004F
FC16
FA65
FB19
FC02
FBD3
FB34
FB18
FB4D
FB29
FAC8
FAC7
FB2B
FB5A
FB2E
FB21
FB58
FB53
FAF3
FAE5
FB67
FB8B
FAB4
FA2F
FC0A
0048
045C
05DD
0512
0420
043F
04C5
04CE
0498
04C3
0523
0530
0504
0507
0520
04EC
0499
04A9
04FD
04EE
0478
0484
0561
0598
0359
FF10
FB6A
FA5F
FB2B
FBD0
FB9B
FB49
FB54
FB56
FB06
FACA
FAF2
FB24
FAFC
FAC8
FB03
FB6C
FB5C
FAFD
FB1C
FBA6
FB7E
FA7C
FA76
FD2A
01A5
04FF
05A3
04BF
044F
04B4
04F5
04AB
0486
04E7
0533
04EE
0497
04C0
0511
04FC
04BF
04E4
0524
04D8
0451
0496
0587
0546
0254
FDE1
FAD0
FA78
FB64
FBA0
FB18
FADF
FB31
FB51
FAFD
FACC
FB16
FB65
FB4F
FB19
FB29
FB4A
FB20
FAF9
FB5B
FBD0
FB60
FA72
FB0F
FE5B
02B3
054E
0560
0491
0482
050D
0539
04EC
04DB
052E
0546
04E2
0495
04C0
04F6
04D5
04B7
04EB
04F9
047D
0428
04CB
059A
048C
00E8
FCA1
FA5E
FA96
FB73
FB71
FAEF
FAE2
FB2C
FB18
FAB8
FAB1
FB0F
FB41
FB17
FB00
FB2B
FB3C
FB0E
FB1A
FB9E
FBDB
FB26
FA86
FC02
FFF0
0404
05D1
0569
04B1
04BE
0503
04DA
049D
04D7
0541
053E
04EA
04E2
052D
052B
04C3
04A0
04F8
050F
048F
0457
0505
0557
035B
FF2B
FB50
F9FE
FAB6
FB63
FB23
FAD9
FB40
FBB1
FB6D
FAE3
FAE1
FB33
FB1F
FAB3
FAA6
FB17
FB5E
FB32
FB1B
FB5F
FB5E
FAC3
FACC
FD2F
018B
0534
061A
0511
0459
04C1
0547
051C
04B1
04B7
0503
050B
04DA
04E2
051D
0517
04C9
04AA
04D1
04C3
0483
04C9
0591
0546
0275
FE00
FA92
F9CB
FAC3
FB88
FB69
FB14
FB11
FB16
FAE5
FAD9
FB26
FB56
FB17
FADC
FB17
FB69
FB4A
FB0B
FB50
FBC7
FB74
FA87
FAE2
FDEF
0273
0590
05F9
0515
04BC
0502
04FA
0496
049A
0520
0568
0517
04C0
04DB
0505
04C0
0466
0494
04FF
04D9
0454
0487
055E
04EA
01C2
FD4B
FA6A
FA34
FB18
FB42
FABF
FAAE
FB44
FB99
FB3B
FAD0
FAEC
FB35
FB2E
FB15
FB4A
FB81
FB57
FB26
FB6C
FBBD
FB4F
FA9B
FB70
FEC1
02FF
0589
0591
04B5
04A7
0545
057F
0520
04CE
04D1
04DB
04C6
04C4
04CE
049F
0451
0465
04EC
0530
04BB
044B
04C8
0573
043F
008E
FC70
FA6E
FAB9
FB7E
FB73
FAFF
FAEE
FB21
FB10
FAD6
FAF7
FB60
FB78
FB33
FB2B
FB83
FB98
FB24
FAE0
FB43
FB88
FAEE
FA7B
FC21
001C
0420
05CB
053C
0471
0498
050B
04F7
04B6
04F3
0565
0556
04DE
04A0
04B4
04A8
0474
048D
04F6
050A
049B
047E
053C
0599
03AA
FF82
FBAA
FA50
FAEE
FB7A
FB25
FAC3
FAFF
FB58
FB2B
FAB9
FAA4
FAEF
FB1F
FB21
FB46
FB81
FB68
FB17
FB35
FBB1
FB91
FAA6
FA95
FD06
0137
047C
053D
0488
0448
04DF
0542
04F7
04BB
0518
057C
054A
04E2
04E3
050F
04D7
046E
046D
04B4
0497
042D
0464
054F
0545
02AD
FE68
FB3F
FABA
FB99
FBDF
FB50
FB01
FB4D
FB7E
FB2D
FADA
FAF6
FB31
FB20
FAFF
FB36
FB8C
FB81
FB42
FB6C
FBCB
FB78
FAA4
FB1A
FE15
023C
04E9
0528
0469
044C
04C7
04E1
0473
043B
0486
04C9
04AF
04A7
04F7
0529
04E5
049E
04C0
04D8
0463
03FE
0492
0582
04C1
015B
FD1B
FABE
FAE6
FBBF
FBAD
FB13
FB08
FB7C
FBA2
FB67
FB66
FBB3
FBBC
FB56
FB0E
FB33
FB50
FB0A
FAE0
FB59
FBE0
FB80
FAD3
FBDA
FF5D
0365
0563
0513
0450
0468
04E2
04D9
0473
0467
04BB
04D3
0488
045B
047E
048C
0467
0489
050B
0531
04A1
0440
04D3
054C
03B1
FFC5
FBD2
FA35
FAD4
FBB2
FB98
FB23
FB36
FB99
FBA6
FB77
FB7E
FB99
FB65
FB1B
FB3C
FBA1
FBA5
FB42
FB33
FBB0
FBDB
FB26
FACC
FCBA
00D9
04A0
05E3
0528
047A
04B1
0506
04C9
045D
0456
0489
0487
0463
047D
04BE
04C0
0496
04AC
04DE
048B
03D5
03D4
04CF
0520
02F4
FECF
FB4A
FA39
FAE5
FB75
FB38
FAE7
FB13
FB5D
FB59
FB4E
FB8E
FBC2
FB8B
FB35
FB3C
FB7A
FB87
FB82
FBC6
FC11
FBB7
FB01
FB73
FE1C
01F1
04AC
0548
04D5
04BA
050F
052E
0505
04F8
04FD
04BE
045E
0464
04C5
04DC
046E
0420
046E
04BD
044A
03A4
0411
0544
04FE
01CF
FD4B
FA73
FA57
FB68
FBCC
FB59
FAEB
FAD3
FAC0
FAAC
FAF7
FB83
FBA5
FB3A
FAFE
FB5F
FBCA
FBB4
FB8F
FBE4
FC26
FB82
FAAB
FBA2
FF30
0372
05BB
0586
04A3
0493
04F8
04E5
048B
04AE
0535
055E
0506
04CE
04F8
050D
04C7
0492
04BE
04D1
0452
03E4
046F
053B
0423
0054
FBE3
F9AE
FA2E
FB62
FB95
FB09
FADA
FB30
FB54
FAFE
FAB5
FAD6
FB10
FB09
FAF0
FB01
FB16
FB18
FB4F
FBC2
FBD0
FB2B
FAE9
FCA6
006C
0431
05E5
058A
04CC
04CB
0521
0513
04C6
04C8
0515
0547
0552
0568
0569
0517
04B4
04C0
051B
050D
046B
0410
0491
04D2
0307
FF2F
FB8E
FA31
FAB0
FB32
FAEB
FAA0
FAF8
FB70
FB54
FAE1
FAD1
FB23
FB2D
FABF
FA71
FA9D
FAE3
FAF6
FB32
FBC2
FBEF
FB44
FAE7
FCBA
00D1
04CD
064E
0590
04C1
0514
059C
052E
0447
0429
04EA
056D
0520
04B8
04E9
0557
0544
04CD
04AA
04EF
04EB
046E
0453
051F
05A8
0413
0034
FC26
FA28
FA6C
FB4D
FB6E
FAF6
FAC3
FB15
FB63
FB4E
FB0F
FAF7
FAF6
FADE
FACA
FAF5
FB3F
FB44
FAF6
FACD
FB21
FB88
FB5C
FAE8
FB8E
FE4D
023B
051F
05B0
04CC
0441
04B1
053C
050E
048A
0492
0528
057C
052F
04CE
04DB
050B
04E1
0496
04B6
0519
0503
046A
0440
04F5
0536
0333
FF23
FB87
FA71
FB42
FBC4
FB0E
FA42
FA8A
FB65
FB94
FAF7
FA93
FAEF
FB64
FB4E
FB10
FB49
FBAA
FB74
FAD8
FADA
FBAD
FC16
FB3A
FA56
FBA8
FF89
039E
0565
04EE
0446
04B5
0581
0580
04D4
047A
04B5
04DB
0494
0465
04B9
0513
04CE
0444
045C
051A
056D
04C5
0414
0483
057A
04E5
01BB
FD86
FADA
FA99
FB67
FBA6
FB33
FAE7
FB17
FB48
FB2A
FB14
FB5B
FBA6
FB7E
FB16
FB13
FB81
FBAF
FB3A
FABA
FAEA
FB77
FB61
FA9E
FAB2
FD14
0137
04CB
060C
055C
046F
044F
04A6
04C9
04AF
04B3
04D7
04CC
0491
0483
04BD
04DE
04A7
0476
04C0
0538
051F
047B
044A
0518
05B7
042F
002D
FBD4
F9B6
FA34
FB71
FBB5
FB23
FAE6
FB55
FBA6
FB4D
FAC8
FAD6
FB59
FB9A
FB62
FB30
FB55
FB79
FB41
FB01
FB2A
FB6F
FB1D
FA87
FB3F
FE57
02AF
05BD
0624
0502
0459
04C6
054D
0513
0481
0471
04E7
0530
0503
04CB
04D7
04DE
0496
0456
048F
04FB
04EE
047A
047B
0523
0515
02C3
FE9E
FB1A
FA1F
FB13
FBDC
FB6E
FAA1
FA93
FB1F
FB66
FB31
FB0E
FB3A
FB43
FAF2
FACF
FB45
FBC8
FB87
FAC6
FAA7
FB70
FBEF
FB3B
FA7A
FBE4
FFDF
040B
05C4
04FC
03E5
041A
0511
0578
051E
04DE
051B
0546
04F7
049F
04C8
0526
0519
04BB
04B7
051D
0526
047A
03F8
048F
0581
04C1
0169
FD20
FA8B
FA83
FB8B
FBDA
FB45
FACC
FAEF
FB26
FAEC
FA90
FAA1
FB0B
FB44
FB21
FAFC
FB08
FB03
FACB
FAD2
FB6D
FC07
FBB2
FAAE
FABE
FD4F
018F
04F3
05CC
04E2
0433
0499
0545
0549
04D6
04B6
050F
0556
053D
050B
04FD
04DF
0490
0476
04EB
0570
0531
0456
0412
04EE
0585
03D8
FFD2
FBC6
FA07
FA90
FB7A
FB6A
FAC8
FA94
FAE9
FB1F
FAF8
FADA
FAFE
FB12
FADE
FAC8
FB31
FBBC
FBB3
FB1A
FAC7
FB2B
FB95
FB3C
FAB3
FB9E
FEBE
02C3
057A
05F6
052D
0497
04B0
0501
0520
0525
0535
0526
04DC
04A3
04D1
0533
0540
04D8
047B
0492
04D0
04A9
0449
046D
0517
04ED
0290
FE7C
FAFB
F9DB
FAA8
FB7E
FB4B
FAAC
FA9A
FB04
FB29
FAE7
FADA
FB48
FBA2
FB69
FAFA
FAEE
FB29
FB1D
FAE0
FB27
FBFB
FC48
FB6A
FAAE
FC3D
0050
046D
0609
0547
045E
04B2
0580
057C
04CB
0483
04EF
0534
04C9
0449
0468
04D8
04DF
0499
04BC
0547
054B
0464
039A
0406
04F4
0448
010C
FCE3
FA5B
FA41
FB2A
FB7D
FB1A
FAD6
FB0B
FB4B
FB42
FB2E
FB55
FB81
FB60
FB21
FB30
FB7C
FB77
FAF9
FAAF
FB2D
FBF5
FBFC
FB3E
FB47
FD91
0194
04FE
0608
052F
0456
0485
051F
052A
04B0
046D
04A3
04DA
04BA
0491
04B6
04F1
04DE
04A8
04C7
0513
04DD
041A
03C6
047C
0515
03A0
FFD7
FBE2
FA22
FAAF
FB9E
FB8D
FAF8
FAF0
FB67
FB7E
FB04
FABC
FB19
FB88
FB65
FAFC
FB04
FB73
FB8E
FB2E
FB1C
FBC4
FC48
FBA9
FA9F
FB47
FEA0
0305
05BB
05CE
04B8
044F
04C6
0516
04C1
0462
0493
0507
051C
04D0
04AA
04D8
04F0
04B1
046E
0480
04A1
045E
03FE
044C
0535
0532
02C9
FE8C
FAEF
F9D9
FAC4
FBAF
FB82
FAE8
FAE8
FB6B
FB9F
FB4B
FB08
FB32
FB61
FB31
FAF3
FB23
FB89
FB86
FB25
FB20
FBA4
FBD0
FB0E
FA7F
FC15
000C
0427
05F9
0574
0485
048E
0517
051A
04A2
047E
04D3
04EB
047A
042B
0494
0530
0522
048D
0463
04EF
055A
04FB
046E
04A7
052E
044B
012D
FD47
FAE1
FAA6
FB3B
FB39
FAB9
FAB0
FB4F
FBC5
FB7B
FAE4
FAC7
FB36
FB97
FB8D
FB55
FB39
FB21
FAEE
FADA
FB22
FB76
FB46
FAC9
FB3D
FDA2
0156
0467
057C
050E
049D
04E6
0559
0535
049E
044D
048F
04F8
050B
04C8
0479
0448
0444
048E
0518
0563
04F9
043F
0439
0528
05AD
0402
0023
FC30
FA5E
FAC1
FB97
FB79
FAB3
FA5F
FACE
FB5A
FB79
FB56
FB4B
FB52
FB45
FB4B
FB95
FBD6
FB8B
FAD8
FA90
FB1F
FBC2
FB7C
FAAD
FB1B
FDEE
0215
0529
05D5
04F8
044E
048C
0517
0544
052C
0526
0514
04A5
0412
03FF
0493
0525
0511
048D
0453
04A0
04FD
0512
051D
053C
04B1
0289
FF0E
FBF1
FAA9
FAF8
FB78
FB59
FB06
FB13
FB48
FB1E
FABB
FACB
FB61
FBBF
FB6D
FAF0
FAFE
FB69
FB75
FB13
FAF9
FB63
FB80
FAC8
FA5B
FC0C
FFF4
03CF
0563
04DC
0439
04A3
055B
0543
048D
0448
04C2
053C
0528
04EC
0508
053B
0502
0490
0488
04E6
04F3
0473
0437
04ED
05B6
04C9
0194
FDAA
FB38
FADE
FB73
FBA5
FB3D
FACE
FAC7
FB11
FB5D
FB68
FB17
FA8F
FA45
FA9C
FB53
FBA8
FB3C
FAA5
FABE
FB81
FBF5
FB6D
FA8F
FAD8
FD1B
00A7
03E2
059D
05BD
04F7
042A
03EF
0471
0550
05DA
0593
04C0
0438
0499
0589
0604
0575
046F
03FF
0478
0526
054B
050A
04F2
04D2
0394
00A1
FD06
FAB2
FA79
FB53
FBB8
FB4C
FADC
FAFC
FB4B
FB27
FAA4
FA60
FAA7
FB1E
FB49
FB1D
FADE
FACA
FAFE
FB6D
FBBD
FB69
FA84
FA27
FBA2
FF04
02B5
04E4
0534
04BE
049B
04DC
050A
0506
0508
0512
04EE
04B6
04D4
054F
0590
052D
049D
04A6
0527
0530
046D
03E4
0499
05CD
0564
0258
FE25
FB5C
FAF2
FB98
FBA3
FAE9
FA6F
FAB6
FB21
FB07
FAB1
FAD3
FB6A
FBB5
FB4D
FAC7
FAE3
FB76
FB9F
FB08
FA76
FABE
FB95
FBFB
FBD0
FC65
FEF7
02E1
05DD
064E
04E3
03BC
0417
0548
05EF
0599
04F2
04A9
04BB
04C6
04AA
0497
04AE
04D1
04DC
04D1
04D2
04FE
0552
0581
04F1
0327
0062
FD92
FB94
FA8E
FA3A
FA7B
FB41
FC05
FBF2
FAE8
F9F6
FA37
FB60
FC11
FB9D
FADD
FAD0
FB2C
FAFE
FA68
FA97
FBD1
FC86
FB5C
F996
FA2F
FE3A
032D
059C
0503
03DE
0449
05A7
0610
051B
042F
0467
052D
0556
04D0
047D
04D0
0547
054F
0509
04EC
0505
04FE
04B9
047F
0483
0462
0353
00E7
FD95
FAA0
F94C
F9E1
FB49
FC00
FB7F
FAA7
FA85
FB11
FB67
FB1C
FABF
FAEB
FB56
FB4C
FAD1
FAAC
FB36
FBC4
FB95
FAED
FAA7
FAF8
FB53
FB9A
FCB4
FF66
02F6
0581
05EF
0507
0461
04A2
0528
0538
04F3
04F4
0565
05C0
057B
04B7
042A
0455
04F5
0547
04F1
046E
047C
051C
0581
051A
045A
03F6
0379
017C
FDB2
FA0F
F910
FADD
FCDF
FCA3
FA8F
F91E
F9B2
FB26
FBA1
FAFB
FA90
FB27
FBFC
FBFD
FB38
FA9D
FAB4
FB20
FB57
FB44
FB17
FADD
FAB6
FB30
FCF3
FFF3
0332
056F
060F
0573
049D
0468
04EE
0590
059D
0512
0492
049A
04EB
04EC
048F
0461
04B5
0522
0519
04AC
0461
0471
049F
04C5
0500
0501
03BE
0087
FC5F
F994
F97D
FB0C
FC0B
FB81
FA70
FA41
FB0F
FBC8
FBA1
FAEF
FA92
FAF0
FBA2
FBFE
FBBB
FB2C
FAFA
FB6E
FC08
FBF3
FB0D
FA36
FA65
FBB7
FD9E
FFD8
028E
0560
06FA
065C
046B
035C
0442
05D0
060B
04C3
03AC
0412
0547
05B1
04DE
03E3
03D8
049B
0540
0535
04AC
042C
042B
04CC
058A
0546
031C
FF74
FBF4
FA1E
FA17
FAD7
FB63
FB7F
FB60
FB37
FB2D
FB64
FBAF
FB96
FB01
FA97
FB02
FBE6
FC20
FB42
FA44
FA5C
FB66
FC17
FBAC
FAD4
FAAA
FB8A
FD43
FFE1
034D
0660
0754
05B9
0377
02FE
0498
0634
05F9
046E
038C
0439
056A
05B0
04E6
0416
041D
04CB
0550
0521
0474
0410
049B
05CD
0655
04E6
01A1
FE2F
FC21
FB7A
FB19
FA6E
FA17
FAB3
FBAE
FBD9
FAF9
FA27
FA62
FB54
FBE5
FBB4
FB5D
FB61
FB6F
FB12
FA9F
FADE
FBC8
FC36
FB44
F9B0
F969
FB82
FF03
01FC
0385
0453
0555
0650
0642
04FD
03C4
03EA
0533
0624
05CC
04C7
0433
0444
0464
045D
04B1
057D
05D8
04F5
039D
0390
0541
06E8
066E
03D2
00E5
FEED
FD64
FB5E
F956
F8CD
FA2D
FBF6
FC5E
FB3D
F9FF
F9E9
FAEA
FBF5
FC24
FB73
FAA0
FA7B
FB19
FBB2
FB86
FAD6
FAB1
FB74
FC03
FB35
F9D1
FA38
FD8E
0205
04BF
0503
04A3
053A
0629
05F2
04C5
0459
0553
0631
0575
03E7
0391
04DA
05F2
0561
040D
03E7
0523
05F4
0527
03DC
03F8
057F
065E
04E2
0191
FE48
FC2B
FB02
FA4C
FA27
FAD3
FBC9
FBF4
FAF5
F9C3
F9AC
FADB
FC19
FC29
FB28
FA58
FA9A
FB75
FBD5
FB79
FB20
FB46
FB62
FAC6
F9F0
FA44
FC62
FF41
0168
02A1
03E6
05A0
06C8
0630
0450
030B
03B9
05B3
070D
0682
049E
0320
0358
04F3
064C
0604
046D
0345
03C5
0536
05E7
055C
04BF
04E0
04A8
026E
FE8F
FB79
FAD6
FB8F
FB78
FA53
F9EA
FB1D
FC56
FBB6
F9E6
F94D
FAC8
FC82
FC7C
FB26
FA7D
FB23
FBC2
FB49
FA90
FAE4
FBDB
FBD3
FA75
F993
FB11
FEA7
0240
0446
04DF
050C
053A
0527
04C0
0470
049D
052A
059F
0593
0508
046B
043D
0489
04DA
04CA
048A
049C
0509
053E
04E8
049C
050C
05B4
04F1
01F0
FDF2
FB2B
FA84
FAF9
FB2E
FAF4
FAFF
FB86
FBD5
FB4F
FA63
FA15
FAD0
FBE8
FC49
FB8D
FA6E
FA27
FB30
FC8A
FCA8
FB37
F9A6
F991
FAE1
FC1C
FC8E
FD6D
001F
03EC
066A
064D
04E0
0432
049E
0502
04CF
04BC
0544
059A
04DF
03C9
03DF
053E
0634
0580
040B
039C
047A
055F
0575
054D
0583
0569
03DB
00FD
FE3D
FC95
FB9A
FA99
F9D5
FA0B
FB17
FBEA
FBCA
FB0B
FA75
FA72
FAF2
FBA8
FC0F
FBA3
FA8C
F9E3
FA99
FC13
FC99
FB79
FA01
F9D8
FAE4
FBCC
FC43
FDA7
00E5
049C
0664
05AD
0460
045F
055B
05BB
0506
0458
049C
054B
0554
04A6
0438
04A7
0571
05A2
04FC
042A
03F3
0485
0560
05C7
0560
046B
0350
01E1
FF86
FC54
F9A6
F908
FA77
FC2F
FC75
FB5E
FA5A
FA61
FB08
FB7B
FB98
FBA5
FB8F
FB1C
FA97
FAAC
FB6C
FC04
FBC5
FB03
FA97
FAB4
FAE0
FB13
FC21
FE9E
01CF
0441
0545
055E
054B
0534
04E5
046D
042B
0458
04CC
053A
0554
04E3
0411
03A6
0459
05B5
0637
0513
0375
0352
0506
06C2
06A0
04AE
0268
009F
FEC7
FC72
FA72
F9E7
FAA6
FB73
FB8A
FB50
FB59
FB81
FB5A
FB0E
FB2D
FBB3
FBE6
FB5B
FA9B
FA78
FB07
FBAC
FBE3
FB96
FAEC
FA35
FA0C
FB09
FD1D
FF80
018D
035D
0531
0680
0655
04C6
035B
037A
04CE
05CC
0591
04A7
0405
03F7
044B
04F2
05CD
062E
055C
03D2
0327
043F
0606
069B
0579
03C9
028E
0153
FF11
FBFF
F9AE
F95C
FA9B
FBEA
FC3E
FBAF
FAFB
FABC
FB0A
FB86
FBAE
FB60
FAFC
FAE7
FB09
FB01
FAD4
FB01
FBA9
FC09
FB4E
F9EC
F96F
FAD3
FD71
FFF3
01E3
03B4
0578
0662
05D4
0472
03A0
0406
0501
058E
0559
04C2
044B
0446
04C7
057D
05CA
0555
0485
0416
0448
04C6
0541
05C5
0621
057F
0331
FFD6
FD0D
FBC3
FB5E
FADF
FA53
FA81
FB72
FC23
FBC7
FACB
FA2F
FA51
FACD
FB4C
FBC4
FBE3
FB29
F9ED
F991
FAEA
FCCC
FD0B
FB13
F8C6
F889
FAD2
FE1C
00D2
02A0
03E9
04D4
054D
0570
0562
0509
046A
0415
04A0
05AE
0623
0576
046F
0429
04B5
0536
0531
04FF
04EA
04AC
0439
045B
0596
06DD
0640
0332
FF58
FCBF
FBB9
FB27
FA6E
FA30
FAEC
FBDD
FBE3
FB07
FA55
FA69
FAE9
FB4B
FB7A
FB87
FB41
FAA8
FA5D
FAF9
FBFC
FC2F
FB35
FA1F
FA07
FAC0
FB8A
FC8E
FEB9
0213
0517
0635
0590
04A3
046D
04A7
04BF
04CD
0519
055E
0520
048D
044F
04A1
0514
0542
053C
0521
04BF
041B
03F4
04FA
0686
06CD
04D5
01A2
FF06
FDA2
FCB5
FB96
FA9D
FA6E
FAF9
FB98
FBD6
FBA5
FB14
FA5C
FA27
FB08
FC69
FCC3
FB65
F9A4
F970
FB04
FCA4
FCBB
FB7F
FA3A
F9B1
F9E1
FAFD
FD74
00D0
0374
044C
041C
046B
056B
05D9
04F2
03AC
0384
04A5
05CF
05F8
053E
0456
03C0
03D1
04B6
05E8
0626
04D6
0324
02FD
04C5
06B2
06CA
04E5
0248
FFCE
FD60
FB2B
FA25
FAB9
FBCB
FBE1
FB07
FA94
FB2F
FBEB
FBB1
FACF
FA71
FAFB
FBAB
FBD4
FBA0
FB66
FB0C
FAA1
FACA
FBC7
FC84
FBB6
F9F7
F9C2
FCB0
0153
049B
052F
0472
0446
04CF
0511
04C1
0488
04BA
04DE
04A9
048F
04EC
0541
04EA
0444
0448
0508
0568
04B6
03BC
03B1
048C
0537
050F
044A
02F8
008E
FD1D
FA33
F985
FAD1
FBFF
FBA7
FA9D
FA78
FB4D
FBCC
FB50
FAB0
FAE4
FBA7
FC03
FBBD
FB6B
FB59
FB33
FAE3
FB05
FBE0
FC99
FC22
FAC0
F9E9
FA96
FC61
FE69
007F
02D6
04FA
05F2
0586
04B1
047B
04D5
050A
04EC
04E8
051F
051D
049D
0414
0413
0479
04BA
04B7
04C8
04F2
04BA
040F
03C6
048D
05C0
05FE
04D2
0326
01C2
002A
FD92
FA9B
F91D
F9EE
FBA9
FC39
FB4A
FA5F
FAAA
FB9D
FBE7
FB4D
FACD
FB25
FBE1
FC13
FB90
FAFE
FAE3
FB1B
FB4B
FB6A
FB96
FBB5
FB73
FAD5
FA7F
FB54
FDB8
011B
043F
05F9
05FD
0504
0438
0442
04DE
0555
0540
04D0
0471
045A
0486
04D9
0521
0516
0499
040E
0416
04D3
0582
053B
0421
0378
0442
05E1
067D
04D3
016F
FDFE
FBBA
FAAF
FA68
FAA1
FB31
FBA5
FB84
FAFC
FAC1
FB24
FB9A
FB76
FAE3
FAB0
FB3C
FBF0
FC08
FB82
FAFC
FADC
FAFF
FB30
FB69
FB82
FB22
FA67
FA50
FBE9
FF00
022B
0431
051A
0594
05C4
0552
0474
0413
04A4
0563
0553
0498
042E
0479
04CF
049D
0455
04A9
054F
055D
04BB
0464
04E9
0582
0538
0470
0457
04E6
047D
01DF
FDF4
FAE7
F9D8
FA19
FA9C
FB20
FBA9
FBC5
FB1F
FA61
FA9B
FBC3
FC8C
FC07
FADC
FA6C
FB13
FBE4
FBF5
FB56
FAA2
FA47
FA85
FB6D
FC69
FC54
FAE4
F9B8
FB13
FF34
03A7
05C8
0578
04B9
04E9
056A
0535
0494
047E
04F4
0508
0470
0402
0465
050D
050C
0472
042A
049B
052C
054A
0518
04D8
0463
03CC
03DA
04F6
05E2
049B
00CE
FCAD
FAB2
FAF9
FB94
FB32
FA70
FA66
FB04
FB73
FB7B
FB7E
FB7D
FB1C
FA97
FACF
FBE7
FCA4
FBE1
FA4F
F9C9
FAF2
FC64
FCA2
FBDA
FB29
FAE1
FAA5
FAD1
FC83
FFDB
0327
04A1
047A
0461
051D
05B9
0548
0468
0453
0510
0593
0552
04D4
04A4
0492
0459
0448
04B8
052F
04F2
0440
041B
04B6
050B
0485
041F
04D5
059F
043D
003E
FC0F
FA5C
FB0F
FBE2
FB7D
FAC0
FADC
FB6E
FB5E
FABF
FA9E
FB41
FBB9
FB5F
FAD1
FAF0
FB86
FBB5
FB5B
FB2C
FB6C
FB89
FB3B
FB20
FB92
FBBA
FAD7
FA0F
FBA4
0001
0492
065B
0543
03D9
0414
054A
05B8
04F9
0423
040D
0489
0512
0574
0583
04FE
0423
03CF
047A
0560
0556
0470
03F4
0487
0545
0530
04B8
04D5
050E
03A1
FFFF
FC13
FA4C
FACB
FB8A
FB1A
FA47
FA7F
FBA5
FC52
FBCF
FAE4
FA9C
FB10
FBA2
FBE4
FBCE
FB72
FAF6
FAC2
FB19
FB97
FB8D
FB0F
FAF6
FB8A
FBE2
FB49
FACA
FC4F
000F
03D4
0556
04CA
044F
0509
05EB
0590
0458
03D1
0489
0576
057B
04B3
040F
0418
049B
0528
0569
0529
0484
041E
047F
052D
050D
0405
0379
0473
05AD
0492
006B
FBAF
F986
FA6A
FC09
FC47
FB54
FA9B
FAA5
FADB
FADE
FB05
FB82
FBDA
FBA1
FB28
FB01
FB24
FB1C
FAE5
FAF7
FB64
FBA3
FB77
FB6C
FBDB
FC14
FB65
FAB6
FC11
000D
0479
0667
0562
03BE
03B2
04F8
05CA
055C
0492
0472
04E7
0532
0503
04A6
0472
0481
04CA
052B
0549
04E5
0456
043E
049B
04BC
045D
043A
04D5
0511
0315
FEDA
FAEB
F9DF
FB5F
FCA5
FBE7
FA48
F9F1
FB25
FC2D
FBC7
FAAA
FA40
FAD6
FB86
FBA1
FB63
FB4E
FB74
FB95
FB91
FB66
FB14
FAD1
FB04
FBA5
FBF8
FB83
FB34
FCCB
00B3
04EA
06CB
05D1
0409
03A2
04A8
058F
0564
04B6
0481
04E8
0551
0549
04EC
048D
045C
0462
048E
04AB
0492
0473
04A1
0501
050F
04A5
045B
049E
04A3
02F4
FF4D
FB6F
F990
FA1E
FB79
FBEC
FB5A
FAD0
FAEC
FB50
FB68
FB28
FAE6
FADB
FB00
FB34
FB5A
FB5C
FB4B
FB5B
FB9F
FBC6
FB80
FB09
FAF4
FB4D
FB6B
FB0F
FB45
FD6E
0152
04CD
05E3
04E7
0404
04AC
0616
0680
0574
0428
03E8
04A0
053E
050C
0462
0417
0482
052D
0569
0506
0476
044C
0491
04D0
04BD
04B1
051C
0589
04B7
01F4
FE35
FB60
FA82
FAF5
FB56
FB01
FA62
FA1D
FA55
FAC5
FB2D
FB6E
FB7B
FB6F
FB86
FBBF
FBC3
FB58
FAD6
FACF
FB43
FB8E
FB56
FB10
FB4B
FBA5
FB44
FA5F
FAA3
FD6A
01D7
0563
0659
055A
0451
0462
052A
05BB
05B3
0549
04D0
047B
046E
049E
04C9
04BE
049B
0494
04A4
04AD
04C4
050B
0544
04F2
0429
03D6
049B
0595
04E1
01C0
FDB9
FB17
FAA5
FB3F
FB80
FB22
FAB8
FA9F
FABC
FAFD
FB73
FBE0
FBC6
FB1F
FA99
FAC2
FB52
FB9E
FB85
FB6B
FB73
FB55
FB0E
FB15
FB92
FBC5
FB06
FA37
FB3F
FEC1
02E2
0524
0502
0430
044E
052F
059D
0525
0480
0465
04B3
04E8
04DE
04B9
048D
0466
0474
04C3
04FD
04D3
0485
0491
04E9
04EF
0482
046B
0534
05D6
047B
00C3
FCA8
FA80
FA9A
FB5F
FB7E
FB2E
FB35
FB94
FBAB
FB50
FB02
FB18
FB4E
FB59
FB63
FB98
FBB1
FB6B
FB11
FB1A
FB59
FB3D
FACA
FABE
FB5E
FBCC
FB38
FA80
FB9F
FF33
0353
0589
056F
04B1
04B0
0523
0516
0484
043B
0491
04EF
04CE
0477
0476
04C9
0505
04F5
04BF
047F
0446
044C
04B5
052B
051A
0498
0479
051F
0570
03CD
0033
FC9E
FAFB
FB24
FB7A
FB13
FA88
FAB2
FB5D
FBC0
FBA7
FB8E
FBB5
FBBE
FB5F
FAF0
FADA
FB04
FB17
FB19
FB42
FB7D
FB83
FB76
FBBA
FC21
FBD4
FAAC
FA25
FC16
004B
0436
0591
04BC
03EA
0461
0559
0586
04E4
0468
0486
04B9
0484
042A
0426
0471
04B4
04D1
04DE
04D0
049D
0484
04C5
050F
04D5
043E
0440
0530
05AE
03CF
FF93
FB6A
F9C6
FA9A
FBCB
FBC8
FAF4
FA87
FADB
FB51
FB6C
FB5B
FB6E
FB91
FB8F
FB77
FB6B
FB5B
FB39
FB34
FB6A
FB9C
FB7B
FB39
FB3F
FB73
FB36
FA84
FA96
FCBD
0096
0413
058A
054C
04D5
04F2
0539
0528
04EF
04EF
0508
04DC
0481
046B
04A8
04C4
0489
0459
048B
04D7
04D8
04B9
04E2
0523
04ED
0456
0445
0509
0550
035D
FF57
FB97
FA3A
FAF0
FBBB
FB73
FABC
FAA8
FB2A
FB6E
FB28
FADF
FAFF
FB3E
FB29
FAE1
FAE1
FB46
FBB6
FBDE
FBC0
FB7F
FB3D
FB20
FB39
FB4D
FB0C
FAB4
FB40
FD84
0107
041E
0571
0525
046E
043C
0494
0503
0535
0521
04E4
04B1
04B3
04DF
04FA
04EB
04E9
0518
0529
04BA
041C
041A
04D2
054D
04BE
03D2
03F3
0525
0575
031B
FED4
FB53
FA5D
FB1C
FBA3
FB49
FAEB
FB30
FBA1
FB88
FB12
FAF3
FB4C
FB88
FB44
FADB
FACA
FB02
FB26
FB32
FB66
FBAB
FB94
FB10
FABD
FB24
FBE6
FC0A
FB44
FA8F
FB55
FDF4
0156
03F3
0512
0514
04C8
04AA
04BC
04DB
0509
0545
055A
0510
048C
044D
0499
0516
0523
04AE
0455
0497
051A
051B
0485
0417
045B
04DA
04D4
0472
0494
0545
050F
0284
FE4E
FAEA
FA25
FB49
FC35
FBD3
FAE8
FA99
FAEF
FB24
FAF1
FACE
FB0B
FB51
FB45
FB2C
FB74
FBE6
FBE5
FB5F
FB06
FB55
FBD1
FBB0
FB0A
FACF
FB69
FBFF
FB89
FA77
FAA0
FD45
0171
04C3
05B5
04EC
0439
0495
056A
05A9
0529
04A7
04AF
04FA
04F4
0491
0440
043F
0454
044D
045D
04B8
050D
04D4
042E
03E7
0461
04F3
04CE
0446
0474
0575
05A8
035C
FF10
FB4F
FA18
FAE9
FBB6
FB66
FAAD
FAA0
FB3A
FBA6
FB8B
FB67
FBA6
FBF5
FBCD
FB4B
FB08
FB41
FB8A
FB7C
FB4B
FB63
FBB1
FBB7
FB55
FB1B
FB7B
FBF3
FB92
FA72
FA31
FC65
009B
046A
05BE
04E0
03DE
0425
0534
05AC
052C
0489
0475
04A6
047E
041B
041E
04AB
0526
0517
04C8
04C1
04F0
04D4
0465
0442
04B6
051D
04BB
03F2
03F5
050B
05AE
0407
0027
FC3F
FA72
FAC3
FB7E
FB59
FAA9
FA75
FAF4
FB70
FB66
FB25
FB30
FB73
FB6F
FB12
FAD6
FB0D
FB64
FB64
FB23
FB1B
FB62
FB7D
FB2A
FAEB
FB54
FC06
FBF6
FAF1
FA6F
FC34
0031
0434
0601
057B
046B
0453
0504
0564
0510
04AD
04D0
052A
0519
04A3
0467
04B1
0512
050A
04C2
04BD
0500
0513
04C3
0482
04AE
04E6
0489
03D5
03D1
04CE
0574
03EF
0024
FC2B
FA41
FA9B
FB90
FBAE
FB19
FAC8
FB0F
FB62
FB50
FB1D
FB3A
FB81
FB74
FB03
FAAA
FAC1
FB0A
FB21
FB12
FB3F
FBA7
FBCC
FB63
FAE6
FB0B
FBB4
FBEC
FB3E
FAB7
FC0B
FF95
0397
05D2
05B4
049F
0425
0470
04AC
0481
0474
04E4
0559
0538
04BC
04AC
0534
059C
054C
04A5
0469
04A8
04C0
0476
0458
04CF
054E
0506
0433
03FA
04C9
055F
03FA
0071
FC9E
FA97
FABC
FBB4
FC17
FBB1
FB2F
FB09
FB13
FAFC
FACF
FAD1
FB04
FB1B
FAEE
FAC4
FAEC
FB44
FB5E
FB28
FB13
FB65
FBC3
FBAB
FB47
FB4C
FBD6
FC04
FB2F
FA56
FB72
FF1E
036E
05BF
056D
0432
03EC
04AC
0543
051F
04D7
04FE
053F
050E
049F
049F
051F
056A
050C
047F
0479
04E4
050B
04A8
0451
048C
04FB
04DE
0445
041D
04D4
0561
0423
00CE
FCF7
FAA3
FA63
FB1F
FB8A
FB65
FB3A
FB56
FB6A
FB2B
FAD3
FAC7
FAFF
FB16
FAEA
FAD2
FB16
FB76
FB79
FB25
FB05
FB66
FBD3
FBB0
FB1D
FAE9
FB69
FBDF
FB76
FAB6
FB5A
FE62
0295
057B
05DA
04CC
0436
04A1
0515
04D9
0470
04AA
0552
0584
0509
04AA
04FC
057D
0559
04B2
046E
04DF
054A
050D
0493
049D
04FF
04E6
0441
0416
0501
05E5
04D1
0151
FD2D
FAAE
FA72
FB47
FBC9
FBA2
FB46
FB0E
FAED
FAC9
FAB5
FACF
FB03
FB18
FAF8
FACF
FACF
FAF5
FB0D
FAFD
FAEF
FB16
FB58
FB5D
FB0F
FAD9
FB12
FB5A
FB0D
FA82
FB3C
FE40
0279
0568
05B2
047E
03F9
04CF
05C5
05A8
04D8
0479
04CE
0514
04DA
04A0
04F6
0589
05A1
0532
04EC
0526
055E
050E
048D
0499
0529
0561
04CC
0422
0455
0513
04C9
0258
FE88
FB5E
FA32
FA96
FB36
FB51
FB20
FB18
FB3A
FB46
FB32
FB33
FB4F
FB4D
FB12
FAD8
FADC
FAFE
FAED
FAAB
FA9C
FAF6
FB5F
FB60
FB11
FB00
FB63
FBA9
FB38
FA89
FB11
FDC7
01D2
0504
05E2
04FB
041B
0454
0514
053B
049B
0413
044C
04DF
0503
04AD
0487
04EB
0566
056F
0526
0504
0513
04F3
049F
0493
0500
0554
04FC
0469
0496
0567
053A
02AF
FE82
FB17
FA10
FAD8
FBAA
FB8F
FAFF
FAD0
FB22
FB80
FB9B
FB87
FB65
FB38
FB0D
FB03
FB14
FB0B
FAD0
FAA2
FAD4
FB4F
FB92
FB3F
FAA1
FA6D
FAF0
FB97
FB94
FB01
FB22
FD33
00F3
0486
0620
05AF
04B5
0480
04F5
0529
04C3
0453
0465
04C7
04F0
04D0
04D0
051F
056C
0563
051F
04F0
04DB
04B1
048C
04BF
0544
0586
051B
0478
0475
050F
04FA
02E2
FF1A
FB96
FA16
FA7C
FB3A
FB2A
FA9E
FA8D
FB2F
FBCA
FBC0
FB4D
FB0F
FB26
FB2D
FAEB
FAA3
FA96
FAA7
FAA6
FAB2
FAFC
FB47
FB2C
FACA
FAD0
FB86
FC2B
FBC5
FAA0
FA6E
FC94
007E
040E
05A5
0575
04E4
04EE
0564
0593
053A
04C8
04B7
04F7
051B
04F1
04B7
04BB
04F3
050E
04EC
04C7
04DE
051A
0539
0536
0531
0516
04B7
0455
0490
0561
0580
0379
FF7F
FBA9
FA00
FA79
FB5A
FB5F
FAE7
FAE3
FB52
FB69
FAEA
FA80
FAC3
FB5F
FB96
FB42
FAE9
FAF0
FB27
FB3C
FB3E
FB5E
FB70
FB19
FA7E
FA4C
FADF
FBA2
FBAE
FB04
FAEC
FCBC
004C
03DA
05A2
058A
04EC
04F3
0576
058C
04EF
0452
0460
04D9
0502
04B3
047F
04C4
051F
0508
049F
0474
04B5
04F8
04F3
04E3
050D
052C
04D3
0448
045A
0521
0555
0376
FFAB
FBED
FA29
FA6B
FB30
FB3E
FAC6
FAAB
FB22
FB83
FB55
FAF7
FB08
FB76
FB95
FB20
FAA0
FAB5
FB43
FBAB
FBA7
FB83
FB83
FB77
FB2D
FAF9
FB4F
FBD9
FBAC
FAAB
FA44
FC23
002C
0434
060D
0596
047F
044C
04EE
055F
0521
04B3
04AC
04F5
0507
04C0
0487
04B8
0524
0555
0523
04DB
04BC
04A5
046A
0448
0496
0515
0517
047D
041F
04AB
0546
0418
007B
FC39
F9F1
FA51
FB94
FBCD
FB00
FA89
FB03
FBA4
FB94
FB0E
FAD4
FB0F
FB3C
FB1D
FB08
FB37
FB56
FB14
FAC2
FAE3
FB5C
FB91
FB4D
FB14
FB54
FBAA
FB61
FA8F
FA70
FC46
FFF0
03BF
05D9
05C2
04A1
0408
047F
0541
0556
04C3
0462
04A7
0519
0517
04C0
04A6
04EF
052A
050B
04DC
04EA
04F7
04A5
0442
0470
0510
052B
0460
03B9
0450
0567
04C9
0162
FCE6
FA2B
FA34
FB6B
FBCB
FB12
FA6E
FAA0
FB34
FB6E
FB4C
FB44
FB70
FB7A
FB2F
FAD5
FAC8
FB03
FB41
FB5A
FB55
FB3A
FB10
FB00
FB42
FBBD
FBF1
FB79
FAB2
FAA7
FC3A
FF48
02A3
04F8
05BD
0569
04E3
04B8
04D3
04D6
04A5
047E
0498
04D2
04DE
04B1
049A
04D7
053E
0570
0550
0511
04D7
049E
0470
0478
04A4
048F
040E
03B9
0448
0543
04EC
020B
FDBA
FA9C
FA1D
FB18
FB87
FAE8
FA61
FAC6
FB7F
FB91
FB12
FAE3
FB4F
FBB0
FB87
FB2D
FB22
FB3D
FB0F
FAB9
FABE
FB28
FB72
FB51
FB21
FB4F
FBB8
FBE6
FBBC
FB75
FB2E
FAFC
FB72
FD66
00B6
03E7
0578
056B
04F1
04DF
0504
04F2
04CB
04E2
0513
04F3
0496
0483
04D4
04FF
04B3
0461
0480
04CE
04C0
046A
0452
048C
04A0
0460
0448
04AE
0517
04E7
047B
04A5
0513
0425
0103
FD18
FABA
FA8F
FB28
FB16
FA8E
FA9A
FB5A
FBE7
FBB5
FB40
FB2D
FB5B
FB52
FB1F
FB35
FB9D
FBE3
FBCB
FB95
FB88
FB8C
FB78
FB6D
FB97
FBC3
FBA8
FB6D
FB7D
FBC0
FB91
FAE7
FB02
FD39
0128
04A6
05E7
0536
0450
0453
04DE
0518
04E0
04AB
04B0
04C0
04C4
04E1
0513
050E
04B3
045A
045D
0490
0482
0430
0407
0431
045E
0457
0462
04AC
04D4
047E
041F
0475
0519
0459
012E
FCF7
FA57
FA5A
FB7E
FBD3
FB36
FAD7
FB31
FB84
FB3D
FADD
FB18
FBB6
FBED
FB9C
FB63
FB90
FBB3
FB76
FB38
FB60
FBA4
FB96
FB68
FB8D
FBDB
FBC5
FB5A
FB4B
FBC0
FBDF
FB34
FAF7
FCE9
00D9
045E
0584
04EA
0481
04FA
0569
0519
048A
0470
0496
0469
040B
041D
0499
04C6
0468
0434
04A4
0520
04E6
0442
040A
0452
046C
0423
0416
0498
04FA
0496
040C
047D
0584
0518
01FC
FD9A
FAA1
FA25
FAE6
FB45
FB06
FADF
FB21
FB66
FB6A
FB6E
FBAC
FBE6
FBC8
FB71
FB3C
FB3E
FB4D
FB5E
FB83
FBA5
FB9B
FB81
FB9E
FBE2
FBCF
FB3D
FAD0
FB2C
FBDC
FBB9
FAAB
FA5F
FC8D
00C3
048C
05FB
0571
04AA
0491
04B4
048E
046A
04AB
04F4
04B6
042C
0422
04BA
0526
04CA
0421
0404
0475
04B2
0471
043D
0476
04B3
048C
045D
04AB
0524
050C
0482
0475
04FC
048B
01B2
FD54
FA27
F9C4
FB09
FBD9
FB98
FB3D
FB77
FBD3
FBBE
FB69
FB58
FB88
FB93
FB6E
FB69
FB8E
FB84
FB34
FB0C
FB4B
FB9E
FBB2
FBB6
FBD1
FBA8
FB00
FA7A
FAEC
FBF0
FC19
FAFB
FA56
FC4C
0095
047F
05E7
0557
04B0
04AF
04AD
044D
0423
0492
0501
04C3
0432
0432
04D1
0530
04DD
0477
04A2
0504
04E0
044D
0404
043F
0475
045B
0459
04C7
0529
04E6
045D
047F
052F
04D5
0232
FE2C
FB1A
FA4E
FAFD
FB8C
FB61
FB0D
FB1B
FB67
FB8D
FB80
FB68
FB45
FB04
FAD0
FAE5
FB34
FB70
FB7B
FB7A
FB86
FB86
FB77
FB8C
FBD3
FBF6
FBA5
FB31
FB31
FB88
FB65
FA97
FA6C
FC74
006C
0419
0585
04F1
0425
0435
04A9
04C3
04A4
04CD
051B
0509
04A8
049E
051A
0576
0523
0483
0451
048E
0495
0437
0409
046B
04E0
04D5
0484
047D
04B1
04A4
046B
04A8
0531
049A
01C5
FDAA
FABA
FA42
FB30
FBBD
FB85
FB5A
FBA0
FBC3
FB53
FAC4
FABA
FB14
FB35
FAFC
FADB
FB12
FB51
FB58
FB5F
FB9A
FBC3
FB92
FB45
FB4E
FB90
FB97
FB5B
FB53
FB8D
FB6A
FAB9
FAA1
FC9F
0080
0421
05A8
055B
04D4
04DE
04EF
047D
03FA
0414
04A6
04F7
04D4
04BE
04FD
052A
04E8
0483
047D
04C4
04EB
04DC
04D5
04D9
04A6
044F
045C
04EE
054E
04D7
041A
0439
0509
04B8
01EB
FDB6
FAAA
FA12
FAE7
FB7A
FB65
FB59
FB9D
FBA1
FB0F
FA7D
FA9B
FB39
FBA0
FB8D
FB5B
FB4D
FB43
FB20
FB11
FB34
FB50
FB2F
FB02
FB14
FB43
FB34
FB09
FB44
FBD5
FBE4
FB21
FAD0
FCA8
0098
0464
05E9
054F
0478
049F
0534
0535
04B8
0491
04F9
0549
0502
047A
0448
0482
04D2
0501
0513
04FD
04AF
0469
0490
0506
052F
04C9
0458
045F
048F
045A
040A
047B
0579
053B
024A
FDB0
FA4B
F9C3
FAEC
FB94
FB1A
FA91
FAC2
FB2F
FB21
FAD2
FAEA
FB56
FB63
FAE8
FA95
FAE7
FB78
FBA5
FB74
FB4F
FB48
FB33
FB2D
FB70
FBBF
FB97
FB0F
FAF2
FB88
FBEC
FB4A
FA96
FBE5
FFC1
0402
0610
05AB
04B8
04AE
0531
0544
04D8
04A6
04F0
053B
0530
050D
0517
0525
0514
051A
0552
0555
04D9
044C
044A
04A9
04BA
0462
044A
04BA
04FD
047A
03EE
0487
05C5
0568
021F
FD89
FA9C
FA69
FB5B
FB8C
FAE7
FA84
FACE
FB1D
FAF8
FAC4
FAFD
FB5E
FB58
FAFA
FAC5
FAE0
FAFE
FB04
FB27
FB6B
FB6D
FB09
FABB
FB06
FB9F
FBC8
FB6A
FB33
FB68
FB59
FA8E
FA21
FBE3
0001
0443
0635
05B9
04C7
04DE
058B
0599
04F0
0480
04C1
0524
050C
04BB
04C6
0532
0579
055F
052C
050C
04D6
0485
0471
04B8
04F0
04C2
0488
04B5
0504
04DB
046A
049D
0570
052E
023D
FD91
FA28
F9C6
FB18
FBB5
FB0E
FA78
FACF
FB54
FB16
FA6E
FA5D
FAFA
FB67
FB2B
FACE
FADD
FB1C
FB16
FAEA
FAE8
FAF3
FAD2
FAC7
FB2B
FBAA
FBA1
FB2F
FB29
FBBE
FBEA
FB03
FA59
FC1A
0068
04AC
065B
05AD
04C2
04D0
0537
0520
04C7
04D1
051F
051E
04CB
04B8
0505
052D
04F5
04DA
0533
057E
0533
04B9
04D1
0557
0563
04BD
043D
0484
04F5
04AB
0401
041D
04EA
048F
01AB
FD70
FA89
FA2A
FB0A
FB5C
FAED
FABF
FB3A
FB9B
FB3B
FA8F
FA73
FAF8
FB70
FB73
FB47
FB45
FB56
FB3A
FAFC
FAD5
FACD
FACB
FAE4
FB34
FB81
FB6A
FB13
FB1B
FBA3
FBE6
FB58
FAF0
FC79
004D
0465
064B
05BB
049C
047E
0509
0523
04BE
04A1
04F9
0516
04AB
0464
04DD
0594
0593
04D7
0459
04A0
051F
052E
04FA
04FB
0517
04EF
04A4
0496
04A2
0459
03F9
0451
0540
050E
023C
FDC3
FA7A
F9FF
FB1B
FBAE
FB41
FAE9
FB31
FB72
FB18
FA9A
FAAB
FB27
FB62
FB3D
FB3B
FB84
FB9A
FB2D
FAAC
FA94
FAC2
FADD
FB03
FB5E
FB8C
FB1B
FA76
FA90
FB76
FC02
FB7A
FB01
FC7C
0019
03C5
057E
0561
04F8
0508
0512
04A9
0451
04A8
0564
05AC
0541
04B3
0484
0491
0486
0473
0495
04DF
050C
0513
0510
04F6
04AB
0476
04D8
05AF
0610
0557
043E
0414
04DB
04C5
023E
FE05
FAAA
F9D5
FABB
FB73
FB41
FAE8
FB12
FB55
FB0D
FA77
FA57
FACE
FB3C
FB38
FB17
FB48
FB9C
FB9F
FB5E
FB4C
FB7F
FB87
FB2A
FAD1
FAE2
FB25
FB2A
FAFC
FAF2
FB0C
FB0F
FB53
FCC2
FFB4
0314
053F
05AA
0543
0518
053C
053F
0517
0510
0527
0512
04D7
04D8
0535
058D
0585
053C
0500
04CD
0479
0433
045E
04D9
0507
04BE
049B
0507
056D
050D
044A
044F
0536
0555
0307
FED1
FB22
F9CB
FA54
FB04
FAFB
FAB6
FAD5
FB2A
FB30
FAE3
FAB0
FACC
FAF9
FAEF
FAC4
FAB9
FAD3
FADF
FAD2
FAE3
FB38
FB9B
FBB7
FB85
FB53
FB64
FB97
FB9F
FB6A
FB37
FB30
FB23
FAD2
FA8B
FB27
FD48
0089
03A3
0565
05A1
051F
04C9
04E0
04FF
04D7
04A9
04E6
057F
05D9
058D
04EC
049A
04C6
050B
050C
04E3
04C2
0489
0410
03B1
03FB
04CD
054C
0501
048A
04AD
0526
0511
0461
042D
050B
05BD
0455
0098
FC96
FA81
FA86
FB2F
FB5E
FB33
FB2D
FB41
FB17
FAB9
FA8D
FABE
FB07
FB25
FB2C
FB52
FB88
FB90
FB61
FB3E
FB66
FBC9
FC1B
FC10
FBAA
FB44
FB32
FB5D
FB5B
FB07
FABD
FAD1
FAFF
FACC
FA80
FB52
FE2C
0249
058A
0665
055E
0447
0450
050F
056F
0511
048E
0490
0505
0557
0535
04E3
04C4
04D9
04DF
04C4
04AE
049A
045B
03F9
03D7
042D
0499
0492
043C
0450
050A
059C
053F
047E
049F
05A5
05B3
0326
FECD
FB4D
FA54
FB10
FB8D
FB04
FA48
FA48
FADE
FB46
FB37
FB0B
FB15
FB49
FB75
FB7A
FB50
FB06
FAC0
FA9D
FAA6
FAE2
FB56
FBD5
FC08
FBD0
FB86
FB96
FBE2
FBDE
FB60
FAF5
FB17
FB4F
FAF3
FA99
FBEE
FF8D
03AE
05DA
0597
04AF
04D3
05C6
0630
059B
04DD
04B7
04EF
04F3
04CD
04D5
04FA
04DB
0488
047B
04DF
0546
0545
0504
04F1
051B
0513
0487
03CD
039B
0432
0503
053C
04BC
043F
047A
04F8
0439
0152
FD5B
FAA7
FA63
FB6E
FBCE
FAF2
F9F0
F9D8
FA7A
FAF5
FAFC
FAFC
FB3D
FB6F
FB3C
FADB
FABF
FAEF
FB15
FB11
FB16
FB51
FB9D
FBC1
FBB5
FB9B
FB87
FB5D
FB02
FAAE
FAD8
FBA1
FC68
FC57
FB91
FB88
FDAA
0191
04FD
05F5
04D9
03CE
0437
0565
05EC
0589
0521
0541
0582
055D
04FB
04D4
04E9
04DE
04A5
04A2
04F4
0524
04C1
0412
03BC
03F2
0451
0479
047B
048E
04AA
048C
0428
03ED
045D
053B
0542
032B
FF33
FB59
F9AA
FA52
FB95
FBCC
FB0C
FA8D
FAD1
FB24
FAE8
FA88
FAAD
FB24
FB34
FACB
FA97
FAFD
FB95
FBD4
FBCC
FBDE
FBFE
FBC5
FB3B
FB04
FB7E
FC24
FC38
FBC2
FB70
FBA1
FBEF
FBBC
FB08
FAB5
FBFB
FF3E
034D
0610
065B
0511
042A
049F
0598
05CB
052A
04B5
04DE
0502
04A5
044A
0490
051B
0523
04B1
0490
0502
0552
04E2
041E
03E0
043E
048B
047D
0483
04D3
04CE
0402
032B
0378
04E1
05CC
04A2
015E
FD92
FB0D
FA80
FB2D
FBC0
FB77
FAA9
FA39
FA8D
FB1E
FB39
FAEA
FAD5
FB38
FB91
FB77
FB36
FB3C
FB5E
FB33
FADA
FADA
FB48
FB93
FB66
FB33
FB87
FC1A
FC20
FB82
FB21
FB8F
FC1E
FBCF
FAE8
FAF5
FD0F
0096
03C4
0551
0566
050E
050B
0547
0545
04E8
049A
04C0
0537
057B
0544
04D7
04A7
04C4
04DE
04CF
04C9
04E8
04F9
04CD
0492
0488
049C
048D
0467
046F
04A0
0491
041D
03DA
047A
05AA
05F4
0415
0061
FC99
FA68
FA22
FAD7
FB5E
FB47
FAF9
FAF7
FB2F
FB27
FAC1
FA79
FAB7
FB3F
FB7D
FB50
FB1F
FB30
FB3F
FB04
FAC7
FAFD
FB76
FB86
FB17
FAEB
FB71
FBFB
FBAC
FAD1
FA8C
FB29
FB98
FAFB
FA39
FB37
FE90
02A5
0544
05C8
0543
04F0
0513
0540
052F
0504
0505
0540
056E
0540
04C2
0459
0458
04AA
04F2
0504
0504
051A
052B
050C
04DA
04D0
04DC
04B6
0476
0490
050C
0548
04DD
046A
04CD
05A4
0547
029C
FE94
FB61
FA40
FA87
FADD
FAC2
FA9B
FAAF
FAC8
FABB
FABA
FAFE
FB66
FBA0
FB84
FB35
FAE9
FAB6
FA97
FA90
FAB3
FB01
FB53
FB70
FB4A
FB1C
FB35
FB89
FBA3
FB41
FAD8
FB12
FBB9
FBCB
FAF5
FA88
FC47
002F
041F
05F3
05A7
04F8
052B
05D3
05E4
0545
04C4
04E1
053F
0554
051F
04FF
0517
052E
0514
04E2
04CD
04DB
04E4
04D8
04D0
04E8
050C
051A
050F
0506
0507
04DD
0458
03BF
03C6
04AA
056E
046F
0118
FCDA
F9F7
F971
FA52
FB03
FAF6
FABB
FAD1
FAFA
FACF
FA79
FA74
FAD4
FB2D
FB37
FB1E
FB1E
FB19
FAD7
FA82
FA97
FB34
FBCA
FBB8
FB1A
FAB6
FB00
FB88
FB97
FB38
FB2A
FBBA
FC1F
FB71
FA44
FA94
FDAD
0257
05BD
0647
050E
045A
050D
0619
0639
0580
04E8
04EB
0514
04E9
049C
04A4
04FA
052E
0512
04EA
04F1
04FD
04CC
0477
0458
0491
04D3
04CA
0491
0492
04E2
0512
04C4
044E
0465
0507
0500
0306
FF4E
FBC0
FA30
FA94
FB50
FB27
FA72
FA34
FAA1
FB0E
FB0F
FB02
FB54
FBB9
FBA0
FB1B
FAD4
FB11
FB4B
FB08
FAA6
FAD7
FB89
FBEB
FB88
FAF2
FAF4
FB7A
FBB1
FB43
FADF
FB46
FC18
FC20
FB02
FA21
FB68
FF2A
038B
062E
0657
054A
04AB
04E3
053A
051E
04D0
04C8
04FB
0503
04C2
0483
047B
0487
0484
049D
04FA
0554
0538
04B9
0481
04F9
05A5
05AB
04E9
041D
03FD
0466
04B8
04C7
0502
059A
05C3
043F
00CA
FCC3
FA2A
F9DC
FAEB
FBA8
FB51
FA8B
FA5A
FAE0
FB66
FB6D
FB48
FB7B
FBE2
FBDA
FB2F
FA7E
FA7B
FB12
FB8C
FB75
FB0E
FADA
FAF9
FB2A
FB39
FB28
FAF8
FAAF
FA87
FAD5
FB87
FBEB
FB70
FA93
FAD3
FD40
0136
04BD
0648
0603
054B
0527
0575
058B
0534
04DC
04D4
04E7
04BA
0461
0442
047C
04BA
04B8
04B4
0509
058B
059E
050C
046C
0476
0515
0582
054B
04DF
04D0
04FA
04CA
044F
0453
0524
0595
03F1
0006
FBC6
F986
F9C2
FAF7
FB7E
FB23
FAC7
FAF1
FB40
FB33
FAEC
FAE1
FB27
FB5D
FB44
FB06
FAE2
FAD1
FAB2
FA9F
FAD2
FB39
FB6E
FB3A
FAE2
FAD3
FB14
FB4B
FB47
FB42
FB7E
FBCD
FBB6
FB2E
FAFA
FC27
FEFE
0283
0522
05F2
0565
04B6
04B5
0528
0559
0515
04CC
04DF
0519
0509
04B2
0482
04B4
0505
051E
0513
052B
0554
0533
04BB
0466
0493
04FC
050B
04A8
044D
0453
0487
0499
04AF
0512
055B
0472
01BA
FE0A
FB20
FA09
FA58
FAE1
FB00
FAEF
FB15
FB60
FB71
FB36
FB07
FB2A
FB75
FB8A
FB54
FB16
FB03
FAFD
FAD4
FAA8
FACE
FB4D
FBB0
FB8A
FB09
FAC4
FAF9
FB48
FB52
FB43
FB74
FBAD
FB51
FA7E
FA9A
FD08
015E
0550
06CC
05EB
048E
043B
04CC
053B
0515
04C3
04AC
04A9
0481
0461
048F
04E0
04EB
04AB
0490
04D5
051F
0500
04A3
0492
04E6
0520
04E1
0475
0459
0489
049F
0486
0498
04F4
0523
04CA
045D
0491
0512
0469
019F
FDB0
FAD1
FA3B
FB1A
FBB7
FB64
FAD0
FAD0
FB4E
FB9F
FB79
FB2C
FB14
FB22
FB19
FAED
FAC7
FAC1
FAD4
FAF7
FB28
FB4D
FB3F
FB01
FAD7
FAFC
FB5A
FB9B
FB99
FB78
FB58
FB21
FACC
FAB0
FB31
FC04
FC39
FB61
FA8B
FB89
FEF0
0317
058E
0588
0471
040A
048F
04FE
04CC
048A
04D6
0554
0542
04B0
0477
04F8
0588
0567
04D3
049B
04EE
0531
04F8
04A5
04BB
0510
0518
04D0
04B5
04E5
04DE
0463
040F
0483
054F
056E
04CA
0481
0531
0597
03C3
FFA0
FB88
F9E5
FAB4
FBE5
FBE9
FB23
FACA
FB24
FB6D
FB22
FAAB
FA97
FACA
FACB
FA9A
FAAF
FB29
FB80
FB3B
FAA8
FA7D
FAE9
FB5F
FB5F
FB0E
FAE7
FB07
FB2A
FB2F
FB47
FB81
FB8F
FB40
FAF3
FB25
FB9A
FB91
FAFB
FB0F
FD1A
00C7
0420
057B
0516
0480
04B3
0545
0566
050F
04D9
04FC
0511
04D0
048F
04C3
054B
0594
0566
051C
051C
054A
0547
04FD
04B5
049C
0491
0475
0470
04B1
0513
053E
0521
04F6
04DD
04A7
044C
0441
04E2
0583
049C
0166
FD23
FA36
F9DB
FB0D
FBDF
FB92
FAE9
FAC5
FB0C
FB27
FB08
FB20
FB7C
FB95
FB26
FAA8
FAA4
FAEE
FAF1
FAA2
FA91
FB00
FB6E
FB4F
FADF
FAC0
FB02
FB0E
FAA3
FA54
FAAE
FB56
FB90
FB58
FB57
FBB6
FBB2
FADC
FA4B
FBC9
FF9E
03CF
05F8
05AF
0495
044A
04D4
0534
04F4
0497
04B2
051E
054E
0517
04D0
04C2
04D5
04DB
04E4
0509
0524
04FF
04BE
04CB
0537
058C
0559
04D9
04A2
04DA
0507
04CF
0484
049F
04EB
04CE
0456
0453
0506
0534
0342
FF51
FB8C
FA07
FAA9
FB97
FB81
FAD9
FABA
FB4C
FBB3
FB65
FAC8
FA8D
FAC4
FAFF
FAFA
FADE
FAE0
FAF6
FB03
FB0A
FB1D
FB28
FB17
FB09
FB30
FB6D
FB5F
FAEA
FA83
FAA5
FB2E
FB80
FB56
FB21
FB56
FBA1
FB4A
FA89
FAE0
FD8F
01CE
0533
0610
050F
042B
0469
051F
0552
050D
04FC
0539
0532
04B2
0450
0490
051C
0548
050E
04F8
0535
0551
04FD
0492
0490
04D2
04D7
0495
048A
04DF
050A
04AA
043D
0475
0519
053F
04B0
045A
04EF
0588
045F
00FB
FD13
FAD7
FAB9
FB56
FB54
FAC4
FA86
FAE5
FB50
FB42
FAF3
FAE4
FB28
FB5B
FB3D
FB02
FAF3
FB0E
FB29
FB3A
FB56
FB68
FB4A
FB0F
FB09
FB4B
FB75
FB2E
FAB9
FAB4
FB3E
FBB6
FB8F
FB1D
FB1E
FB8D
FB8C
FABF
FA51
FBF1
FFC5
03E6
061B
05F8
04EA
0470
04B9
050F
050A
04EA
04F2
04F9
04C6
0488
0498
04F0
0526
04F8
04A1
047A
048B
0495
0483
0482
04A4
04BC
04A8
049A
04CA
0508
04EB
0482
045F
04C2
051F
04D0
042C
043E
0522
0546
02FE
FEBF
FB11
F9F5
FAE4
FBC1
FB6C
FAA9
FA9E
FB33
FB7A
FB20
FACE
FB0A
FB7D
FB89
FB38
FB08
FB1B
FB1F
FAF2
FAE4
FB27
FB71
FB66
FB39
FB57
FBB1
FBB6
FB39
FAD6
FB19
FB9F
FB98
FB00
FAC3
FB62
FC09
FBA6
FAAD
FB11
FE0E
0273
05A0
0632
052B
046F
04AC
051D
04FF
049A
049A
050F
0566
054B
0503
04E6
04DE
04AF
047B
0498
0502
054B
0530
04F2
04E8
04FA
04D4
047E
0461
04A0
04D2
0495
0433
0441
04BB
04F7
04AB
0479
04FC
0580
0459
00DE
FC95
F9EC
F9D0
FAF9
FB9F
FB55
FAF4
FB15
FB55
FB24
FAAD
FA8A
FADA
FB22
FB14
FAF9
FB24
FB63
FB4E
FAF4
FACB
FAF9
FB1B
FAE1
FA98
FAB8
FB2F
FB78
FB61
FB46
FB6B
FB84
FB40
FAF8
FB41
FBE2
FBE2
FAF9
FA7C
FC2A
0008
03FC
05E2
0599
04BB
0493
04FE
0530
04FB
04DC
0513
0552
054A
0523
052B
054D
0538
04E8
04AE
04B9
04DC
04E5
04EC
050E
0520
04E5
0488
0480
04E6
0538
04FD
047D
0461
04BB
04E2
0475
0419
04A9
05B7
0587
02DF
FEA8
FB3D
FA29
FACF
FB74
FB3B
FAAF
FAA2
FB0B
FB3D
FAE8
FA6D
FA4B
FA88
FAD6
FB10
FB45
FB74
FB7C
FB54
FB2C
FB21
FB11
FAD9
FAA5
FAC3
FB2B
FB77
FB6D
FB4E
FB70
FBAA
FB89
FB16
FAE7
FB4A
FB9F
FB2B
FA6E
FB13
FE17
0252
055A
05F3
0519
0494
04F2
055D
0525
04B5
04D0
0566
05AF
054A
04B5
0484
04A1
0499
0463
0463
04C8
0538
054F
051C
04EA
04CD
04A4
047D
048D
04C4
04C9
0488
0470
04D7
054B
0514
0453
041B
04F6
05B1
0459
0082
FC22
F9BB
F9EE
FB2B
FBAE
FB33
FAA9
FAB8
FB18
FB3B
FB0D
FAE5
FAF8
FB33
FB72
FBA2
FBA9
FB77
FB34
FB2A
FB62
FB7E
FB3B
FADE
FAF0
FB7C
FBED
FBC8
FB4E
FB1E
FB56
FB80
FB53
FB31
FB7B
FBCF
FB68
FA72
FA65
FCA3
00B9
0483
062B
05C7
04E5
04B9
0527
056A
0534
04D3
0495
0474
0459
045C
048A
04B1
049E
0477
0490
04E6
0511
04D6
047E
0470
0498
048D
043D
041E
0479
04E6
04D6
046A
0458
04DB
0541
04EF
0462
048F
054B
04EF
022E
FDE6
FA8C
F9B2
FA97
FB5C
FB2B
FAB3
FAC3
FB31
FB50
FB03
FAD7
FB21
FB94
FBBF
FBA3
FB85
FB75
FB50
FB21
FB18
FB2F
FB25
FAF0
FAF2
FB6C
FBFC
FBFF
FB75
FB11
FB46
FBAB
FBA2
FB4E
FB5E
FBE0
FBED
FAF7
FA07
FB03
FE84
02E0
05B5
062B
0569
04F3
0527
056C
0558
051D
0504
04ED
04A1
0449
0446
04A4
04FC
04F5
04A3
045C
0450
0471
049F
04C6
04CE
04AF
0494
04B9
050E
0525
04B9
042C
0423
04A6
04F4
0482
03E3
0426
0540
0593
0389
FF8D
FBE4
FA71
FAE8
FB84
FB36
FA8D
FA87
FB1A
FB66
FB0C
FAA8
FAE4
FB82
FBC6
FB80
FB39
FB4C
FB6C
FB37
FAE1
FAEB
FB51
FB7E
FB30
FAE0
FB17
FB9C
FBC2
FB64
FB14
FB39
FB7F
FB78
FB64
FBC2
FC47
FC07
FAFA
FAB5
FCDF
0105
04AB
05DB
0513
0450
0496
0528
050E
0483
046E
04EA
0533
04E2
048C
04CD
054B
053B
0499
0438
0493
0522
0525
04B7
048A
04CB
04EC
049C
0459
04AD
0538
0527
046D
03F0
0443
04C9
049E
03F7
03DD
0474
0446
01E8
FDFE
FADB
FA13
FAF5
FBAC
FB71
FB02
FB34
FBBE
FBC7
FB2A
FA9F
FAB9
FB3C
FB91
FB89
FB5F
FB42
FB2B
FB22
FB48
FB8C
FB97
FB43
FAE7
FAEA
FB3A
FB65
FB4B
FB4D
FBA5
FBEE
FBB7
FB4E
FB6A
FC06
FC20
FB29
FA4F
FB93
FF69
03C7
0616
05CA
049B
044B
04DA
0534
04EB
04A9
04F7
056B
0552
04BC
0458
0476
04B1
049F
0470
0487
04D2
04E6
04A5
0462
045D
0473
0475
0480
04BB
04ED
04BE
0455
043D
049B
04DE
0488
03F7
03E9
0464
04AB
0467
0441
04CB
052B
03B2
0004
FC02
F9FD
FA51
FB51
FB70
FAD5
FA8D
FAE4
FB29
FAE5
FA8B
FAB3
FB2A
FB45
FAEA
FAB2
FB08
FB98
FBD3
FBA7
FB70
FB68
FB6B
FB61
FB69
FB94
FBA9
FB7A
FB3F
FB4A
FB91
FBB5
FB98
FB7B
FB88
FB7E
FB2B
FAE8
FB2E
FBB4
FBA2
FADF
FACE
FCFC
0121
04FC
0682
05DB
04DB
04C8
053E
053C
04B4
047A
04EF
0576
0557
04BB
0464
04A6
0506
04F6
0486
0440
0468
04C5
04F9
04E9
04B8
048D
0479
0481
0499
04A5
0492
0472
045E
0454
0441
0437
0458
048A
047A
041E
0401
04A8
058D
0524
025D
FE17
FAA2
F99E
FA7A
FB4F
FB02
FA35
FA1A
FADF
FB90
FB6A
FAB8
FA5A
FAAA
FB38
FB71
FB45
FB0B
FB01
FB1A
FB30
FB3F
FB54
FB70
FB7D
FB67
FB39
FB14
FB1B
FB47
FB68
FB59
FB39
FB4A
FB90
FBB8
FB86
FB4A
FB89
FC29
FC49
FB5B
FA49
FAF5
FE3D
02B9
05E3
067B
057A
04B7
04EA
0565
055F
04F3
04BE
04EF
0529
0525
0509
0512
0532
0537
051A
04FF
04F6
04E7
04CF
04CC
04E1
04EB
04D8
04CA
04DB
04DF
04A8
0461
0465
04B8
04EA
04BA
0481
04AE
0506
04E3
0449
0426
04FD
05B4
0466
00AD
FC75
FA2D
FA49
FB22
FB1C
FA57
F9F9
FA6F
FB01
FB00
FAAB
FAA7
FB0B
FB58
FB41
FB02
FAE6
FADF
FAC6
FAB1
FACA
FAEE
FADA
FAA0
FAA2
FB01
FB5F
FB63
FB33
FB34
FB69
FB72
FB30
FB00
FB1D
FB36
FAF0
FA9B
FADC
FB95
FBCC
FB0B
FA7D
FBF1
FFAD
03C9
0607
0608
053C
04FD
0542
0550
050B
04FF
0561
05A9
0558
04B6
0474
04C8
053A
0551
0518
04E4
04DD
04EE
0506
0525
053F
053B
051F
050F
050D
04ED
04A7
047C
049C
04CB
04AC
0453
043B
0495
04E9
04CA
049A
0511
05E7
0596
02EA
FEAD
FB27
F9E5
FA5D
FAEA
FABE
FA65
FA89
FAF3
FB03
FAB5
FA9A
FAF3
FB4E
FB32
FACB
FAA5
FAE8
FB38
FB40
FB11
FAE7
FAD3
FACF
FAF0
FB37
FB5F
FB22
FAB5
FAA4
FB19
FB90
FB80
FB1E
FB0C
FB69
FBAB
FB88
FB81
FC10
FCA6
FC39
FAF3
FAA7
FCEF
011A
04A1
05C6
0533
04C1
0531
05B6
057B
04D6
049B
04E6
0517
04E3
04BA
0500
0565
055C
04F1
04B6
04E9
0530
0525
04EB
04DB
04FE
0517
051C
053A
0565
0542
04B4
0429
0418
045C
0471
043E
0429
045C
0468
0404
03C1
0456
053E
04BF
01D3
FDAA
FAAF
FA15
FAE9
FB81
FB5D
FB22
FB41
FB5F
FB1B
FAC1
FACF
FB1C
FB16
FAAA
FA6D
FABF
FB3A
FB40
FAD8
FA99
FAD1
FB28
FB37
FB0E
FAF8
FAFC
FAF6
FAFC
FB49
FBC0
FBF2
FBB8
FB79
FB9D
FBE6
FBD8
FB8C
FBA2
FC27
FC35
FB35
FA32
FB1E
FE99
02E8
0596
05DF
050C
049D
04C4
04DB
04AF
04AD
04FB
0520
04C6
045A
0484
0535
05B2
058C
051C
04F6
0523
0545
052D
0504
04E7
04BF
0485
046B
0488
049D
046C
0429
043A
0490
04A8
0450
0401
0435
049B
0487
0414
042E
0525
05AE
040F
0043
FC5B
FA75
FAA9
FB65
FB72
FB03
FADC
FB0C
FB18
FAE5
FAE7
FB4B
FB96
FB51
FAC6
FA9B
FAED
FB38
FB24
FAEF
FAF4
FB16
FB05
FAD4
FAE6
FB45
FB7B
FB41
FAFA
FB21
FB8C
FBAD
FB6C
FB4B
FB99
FBEB
FBCB
FB7E
FBA0
FC03
FBC2
FAB9
FA5C
FC4A
0036
03E0
055F
04FA
0462
0494
0510
051A
04D7
04DB
051D
050E
049B
0461
04C1
0541
0537
04BA
0479
04B8
0500
04F0
04D2
0514
0580
057D
04F8
048B
049D
04D6
04B2
044F
0435
0478
0499
0460
0441
049D
050E
04F3
0483
0493
0526
04E0
027C
FE97
FB58
FA39
FAB8
FB58
FB73
FB6D
FB8B
FB6B
FAD1
FA55
FAA9
FB8A
FBFA
FB8E
FAF7
FAF9
FB63
FB71
FAF4
FA81
FA8A
FAC7
FACE
FAC2
FB0D
FB9A
FBD6
FB8B
FB35
FB4A
FB91
FB82
FB22
FAF6
FB30
FB68
FB4C
FB2C
FB61
FB8D
FB1A
FA79
FB2F
FE24
0238
052F
05ED
055E
04FB
051F
051F
04AA
0447
046D
04C3
04B2
045D
0466
04EE
0553
0519
049B
0486
04E3
0521
04F9
04CA
04F3
0539
0529
04D2
04A9
04D1
04E6
04A4
0453
045C
04A8
04D1
04CC
04E9
052C
051F
04A1
045D
04E8
0585
0484
0138
FD16
FA6E
FA19
FAE7
FB4C
FB05
FAD3
FB1D
FB78
FB78
FB4D
FB53
FB6D
FB3D
FAD6
FAB2
FAF8
FB38
FB0E
FABB
FAC4
FB2A
FB71
FB5A
FB37
FB5D
FBA0
FB9C
FB5A
FB3E
FB5F
FB64
FB1A
FAD8
FAFB
FB49
FB45
FB00
FB0D
FB89
FBBD
FB2B
FAAF
FBE1
FF24
02E3
0517
0552
04D1
04C4
0517
0523
04DA
04D3
0545
05AD
058E
0523
04F4
0511
0518
04E2
04B5
04C7
04E1
04C3
048E
0495
04D0
04EC
04CE
04BF
04E5
04EC
0488
040D
0414
04A4
0517
04FE
04B6
04C7
0509
04E4
0469
046C
0529
0560
037E
FFA6
FBF6
FA6C
FAE8
FBA8
FB6A
FA91
FA23
FA5B
FAA8
FAB5
FAC7
FB18
FB5D
FB39
FAD5
FAAF
FAEF
FB3E
FB50
FB39
FB2A
FB1B
FB01
FB08
FB58
FBAC
FB97
FB1F
FAD4
FB09
FB59
FB3E
FAE6
FAFE
FB9C
FBFB
FB8C
FADC
FAE0
FB84
FBB3
FB0D
FAE5
FCEC
00F0
04B6
063E
05B8
04E7
04ED
055E
055B
04E3
04A2
04E2
0536
053A
0514
050E
0519
04F1
04AC
04A5
04F6
0549
054B
0511
04DA
04B1
0482
046E
04A9
050D
0524
04CE
0489
04CA
0548
0555
04DD
0485
04B9
04F8
0499
03EB
03E4
048E
046F
0222
FE40
FB0C
FA1D
FAD6
FB78
FB36
FABB
FAD4
FB50
FB78
FB28
FAE4
FAFE
FB2E
FB19
FAD8
FAC5
FAEA
FB08
FB06
FB17
FB53
FB82
FB69
FB23
FAFB
FB06
FB19
FB1A
FB1D
FB24
FB0E
FADF
FADB
FB27
FB6E
FB3B
FABB
FA9F
FB22
FB88
FB19
FA7D
FB72
FECB
0319
05DC
060B
04F1
0474
04FD
0581
0532
047F
043E
0483
04B3
048A
0470
04BB
0518
0503
048C
0448
0490
0515
0553
0524
04C1
0463
0428
0424
0461
04B9
04F1
0506
0528
0558
054A
04E2
0482
049A
04F6
04F9
0496
0490
0553
05D8
046C
00C7
FCCF
FAC6
FAEF
FB8C
FB27
FA33
FA18
FB23
FC20
FBF6
FB01
FA7F
FAEF
FBA4
FBCB
FB69
FB16
FB1C
FB3A
FB29
FB04
FB0E
FB4B
FB89
FBA3
FB96
FB6C
FB3C
FB2C
FB53
FB83
FB6B
FB0F
FADE
FB33
FBCC
FC0F
FBCD
FB6D
FB4C
FB39
FAE5
FA8D
FABE
FB5C
FB87
FADB
FA7C
FC22
FFF3
03E3
05A8
0517
040A
0421
051E
05B7
056F
0500
0525
05A0
05B6
0540
04BF
0499
04AD
04B3
04A9
04AE
04B2
0493
0469
0473
04B2
04DE
04D0
04B4
04BC
04C5
0496
0458
046F
04E9
054B
0532
04D9
04CB
0523
056F
055C
0518
04F0
04C9
046F
042C
048B
054C
0511
02AB
FEB4
FB58
FA43
FB06
FBD0
FB85
FAA6
FA45
FA98
FAF2
FAE3
FAB4
FAD7
FB32
FB5C
FB42
FB38
FB6B
FBA7
FBAF
FB9C
FB9A
FB96
FB5C
FB01
FADF
FB0B
FB28
FAF0
FAA1
FAAE
FB19
FB6B
FB54
FB0F
FAFA
FB1D
FB41
FB63
FBA1
FBD5
FBA1
FB0E
FAB4
FAEF
FB35
FACA
FA18
FAC1
FDD6
0248
05A8
0680
059D
04D2
04F0
055A
0547
04D6
04A2
04D1
04FB
04D8
04A6
04B3
04E8
04FD
04F2
0504
0538
0545
0500
04AA
049E
04D6
04FB
04E2
04C0
04C6
04D8
04C7
04A7
04B8
04EF
04F6
04A0
043A
0428
0467
04A5
04CD
050C
055E
0566
0504
04BE
0508
0541
03FC
00AA
FCAE
FA39
FA1E
FB27
FBAB
FB50
FAE8
FB00
FB3B
FB0B
FA95
FA68
FAAE
FB09
FB30
FB49
FB82
FBAC
FB7F
FB19
FAE1
FAFA
FB20
FB1A
FB0A
FB29
FB68
FB83
FB6C
FB5A
FB69
FB6F
FB3E
FAF9
FAE8
FB12
FB3B
FB40
FB3E
FB51
FB59
FB3B
FB29
FB5A
FB91
FB48
FA97
FA9F
FC96
0047
03E7
05B3
0591
04E3
04D9
0554
058D
0549
0506
0521
0554
0537
04E5
04CE
0507
0531
0506
04BA
049D
04AE
04B3
04A8
04B7
04E3
04F7
04E1
04DA
050A
0537
0517
04C3
04A3
04D5
0500
04DD
049B
0490
04AE
04AB
0490
04AD
0500
050C
0498
0448
04D2
05B6
054A
0283
FE67
FB35
FA2D
FA8B
FACD
FA71
FA21
FA72
FB0E
FB47
FB01
FAB6
FAB9
FAE4
FAF8
FB02
FB28
FB54
FB50
FB28
FB1A
FB38
FB46
FB1A
FAE4
FAEB
FB1D
FB2C
FB03
FAF4
FB2D
FB68
FB44
FAE2
FAC8
FB25
FB92
FBAE
FB9E
FBAE
FBB8
FB59
FABC
FA9C
FB31
FBA2
FB1B
FA58
FB3F
FEA8
0301
05C9
0622
0561
0526
058F
05A8
0515
0486
049B
050C
0536
0511
050E
0546
0557
0511
04D2
04F4
053F
053E
04ED
04B6
04C9
04D6
049C
0460
0483
04E9
0518
04F0
04D3
0504
0536
0503
0499
0483
04DB
051C
04EA
049E
04BA
050A
04E8
0451
0425
04D5
0549
03C6
0011
FC18
FA12
FA47
FB1C
FB2A
FA9E
FA71
FAD4
FB17
FAD2
FA81
FAB3
FB2C
FB4B
FAFD
FACB
FB05
FB54
FB4F
FB19
FB17
FB4B
FB55
FB21
FB09
FB40
FB72
FB45
FAEC
FADC
FB11
FB1A
FAD1
FAA7
FAF9
FB79
FB97
FB5F
FB5C
FBB6
FBE0
FB86
FB2D
FB77
FC04
FBCE
FAD4
FAAB
FCDF
00EC
0480
05D5
055D
04CB
0504
0577
055D
04E0
04B3
04FC
053A
0518
04E1
04FC
0548
0552
0505
04C1
04CC
04FA
0501
04ED
04F5
0516
0512
04E2
04CB
04F1
0514
04F3
04BA
04C2
04FF
0503
04A7
0454
046C
04AB
048A
0421
0418
04A1
0511
04D6
0479
04E0
05AE
0521
0219
FDC4
FAAA
FA0C
FACE
FB24
FAA8
FA4C
FAAF
FB4C
FB67
FB15
FAF4
FB33
FB6C
FB55
FB2A
FB32
FB42
FB0F
FAB5
FA9D
FAE0
FB28
FB31
FB23
FB42
FB7C
FB8B
FB69
FB59
FB78
FB89
FB5F
FB2F
FB46
FB8D
FB9D
FB5C
FB34
FB6D
FBB5
FB8E
FB1D
FB09
FB78
FBAC
FB17
FA8B
FBBC
FF34
0352
05BE
05C6
04D6
0495
0529
0598
055C
04F3
04EE
051E
0506
04B6
04AD
0507
0545
050F
04B8
04BD
050A
051B
04BE
044D
042B
0452
0489
04BF
04F6
050B
04D6
0487
0481
04CC
04FC
04C6
0474
046D
0498
048F
045D
0486
052B
05A1
0545
0488
0484
0555
0578
0354
FF3E
FB6B
F9C4
FA23
FAEC
FB02
FAA9
FAA6
FB0C
FB4C
FB16
FAC6
FAC5
FAFE
FB15
FAF9
FAF6
FB36
FB83
FB98
FB7A
FB60
FB5C
FB56
FB42
FB34
FB34
FB2F
FB25
FB3B
FB71
FB7E
FB29
FABF
FAD1
FB6B
FBF1
FBE9
FBA4
FBB6
FC05
FBE3
FB2C
FAB1
FB18
FBBE
FB78
FA79
FAA5
FD6B
01C7
051B
05E7
051C
0495
04EB
054F
0518
04A2
0490
04C9
04C4
0473
0452
04A0
050C
0536
0537
0553
057B
0563
050D
04D0
04D7
04E0
04B1
047F
04A1
04FA
0510
04C2
047E
049E
04DD
04B9
0443
041B
048F
0521
0531
04DC
04B6
04DA
04B7
0422
03E6
04BD
05CE
0514
019D
FD06
FA08
F9BF
FAD2
FB5A
FAF8
FAAC
FB10
FB92
FB88
FB2C
FB27
FB7B
FB85
FB0B
FA96
FAAA
FB0A
FB22
FAE7
FAD6
FB25
FB74
FB67
FB31
FB33
FB5A
FB50
FB15
FB09
FB4F
FB84
FB58
FB0E
FB16
FB55
FB4B
FAE1
FAA2
FAEC
FB54
FB4B
FB02
FB2A
FBC7
FBFA
FB51
FAEB
FC7B
002B
0407
05E9
059C
04BF
04AD
052E
0548
04C0
044B
0472
04E6
0512
04EC
04DD
0509
0522
04F0
04AE
04B8
050C
0553
055B
0539
0504
04BD
0472
045F
0496
04DA
04E3
04CB
04E5
0530
0543
04E9
0483
0491
04F4
051A
04CF
048F
04B9
04F4
04BB
0453
0489
054C
0528
02BD
FEA1
FB20
F9F6
FAA8
FB6B
FB43
FABE
FABC
FB35
FB80
FB5E
FB33
FB47
FB5A
FB1B
FAB6
FA91
FAB9
FADE
FADE
FAEB
FB1F
FB44
FB2E
FB15
FB48
FBA0
FBA4
FB3C
FAE7
FB07
FB52
FB42
FAE8
FAE3
FB72
FC0A
FC0B
FB9B
FB59
FB71
FB79
FB40
FB3D
FBB5
FC09
FB75
FA80
FAF3
FDE2
0226
054E
060D
0546
04AC
04DB
052E
0513
04CA
04D1
0518
0530
04F6
04BE
04C3
04DB
04C9
04A6
04B3
04ED
0513
050A
0506
0526
0534
04F3
0482
0448
046C
04AB
04B4
0497
049C
04CB
04DE
04AD
0472
0479
04B4
04D9
04D2
04CA
04C5
0490
0430
0425
04B7
0520
03F1
00B3
FCD5
FA7D
FA6B
FB65
FBD3
FB6A
FAFA
FB09
FB41
FB2C
FAEB
FAE7
FB1D
FB30
FB08
FAF7
FB26
FB51
FB36
FB06
FB11
FB40
FB3F
FB0B
FAFD
FB3F
FB8C
FB9A
FB84
FB8C
FBA6
FB8D
FB46
FB32
FB81
FBD5
FBCA
FB81
FB5D
FB60
FB34
FAD8
FAD0
FB64
FC02
FBD3
FB01
FAF4
FCF9
00B2
043C
05E8
05A7
04C9
0480
04E3
0546
0534
04E5
04C5
04DB
04E4
04CD
04CA
04F2
0507
04D7
048D
0479
049B
04AB
0491
0488
04BB
04EF
04D8
0494
0482
04A3
0497
0446
0420
0470
04D5
04C8
046E
0460
04BA
04DD
0466
03D7
03E4
045F
047E
0430
0448
04F8
04DD
0275
FE43
FAB1
F99C
FA86
FB7E
FB5F
FAA5
FA4F
FA91
FAEE
FB1B
FB36
FB5F
FB7B
FB74
FB5B
FB45
FB32
FB20
FB1A
FB23
FB2B
FB28
FB23
FB2D
FB47
FB64
FB78
FB7C
FB71
FB5F
FB5D
FB76
FB92
FB93
FB87
FB93
FBA0
FB74
FB1E
FB01
FB42
FB84
FB78
FB5E
FBAA
FC36
FC55
FBDA
FB81
FBE9
FC7A
FC1C
FB0E
FB27
FDBA
01C5
04E0
05CA
055C
0512
0556
058D
054A
04DF
04C1
04EC
0517
0520
050D
04D9
0494
047B
04B1
04FD
0514
0500
04FA
0508
0503
04E8
04E5
050A
0521
0505
04E5
04FF
0538
0534
04E0
048F
0476
0468
0444
043E
0476
04A8
0492
0465
0472
0496
046D
0408
03F6
0460
04A4
0447
03ED
048B
05A2
0533
0214
FDB4
FABE
FA4C
FB1C
FB72
FAF6
FA7C
FA8E
FAD7
FAD8
FA9C
FA7C
FA92
FABE
FAF4
FB37
FB6A
FB6A
FB41
FB0E
FAD8
FAAA
FAAE
FAEC
FB24
FB13
FAD5
FAC1
FAE9
FB07
FAEF
FADE
FB1F
FB89
FBB4
FB9D
FBA9
FBF2
FC0E
FBC3
FB6E
FB6E
FB8E
FB75
FB49
FB6B
FBB2
FB96
FB25
FB2C
FBFF
FC9D
FBF0
FABB
FB45
FEA1
0311
05D2
060A
052E
04D9
0525
054C
0510
04E8
051E
0563
055F
0537
0535
054F
054E
0531
051D
0517
0511
0519
053A
054F
0534
0509
04FE
04FE
04D5
048F
0473
0499
04AE
046E
041B
0425
047C
0498
0454
0422
0457
04A6
04B4
04AA
04D4
0500
04C9
0459
0443
0489
0470
03B0
033D
040E
054E
04CA
0193
FD6B
FAE6
FAAB
FB39
FB28
FA96
FA5F
FAA9
FAE0
FAB3
FA7A
FA95
FADB
FAFE
FB08
FB31
FB70
FB88
FB6F
FB4E
FB3D
FB35
FB39
FB44
FB3E
FB1F
FB10
FB33
FB64
FB64
FB3D
FB3E
FB80
FBB2
FB87
FB3C
FB49
FBA0
FBC4
FB94
FB87
FBD1
FBFB
FBA5
FB41
FB6C
FBE5
FBE1
FB58
FB32
FBD7
FC49
FB88
FA82
FB7B
FF33
0393
05E6
05BD
04DC
04C2
0537
055B
0517
04F8
052A
0540
0506
04D5
04F9
052C
050E
04C1
04A7
04C9
04E2
04E0
04EC
0511
0527
051A
04FB
04D9
04A8
046E
0453
046C
0495
049B
0481
0470
0464
043A
0405
040E
0452
0480
047D
0499
04EF
050A
0495
0407
041C
04AC
04C6
0420
03BB
0479
0562
0459
00C2
FCA0
FA75
FAA5
FB80
FB98
FB10
FAC4
FAEB
FB10
FAF5
FAD5
FAE8
FB09
FB09
FAFF
FB0D
FB1B
FB09
FAF2
FAFC
FB15
FB22
FB35
FB60
FB74
FB43
FB02
FB0D
FB61
FB99
FB7D
FB55
FB7C
FBCF
FBE1
FBAB
FB94
FBBB
FBC5
FB7E
FB35
FB30
FB33
FAFB
FAD7
FB37
FBD4
FBF2
FB7D
FB41
FBAA
FBE6
FB18
FA27
FB3B
FF08
0376
05C6
0585
049D
04B6
0589
05E7
0586
0522
0534
055C
0528
04CD
04C1
04FC
0516
04F7
04EA
051B
0557
055A
051A
04C0
0483
0483
04B3
04E1
04E9
04DB
04D7
04D5
04B4
047B
046B
04A5
04E7
04DE
04AF
04C2
050C
0514
04BD
048B
04CB
04FE
04A2
041C
043B
04E6
0516
0470
040B
04DD
05C9
0475
0055
FBCA
F99B
F9F7
FADB
FADA
FA6E
FA8C
FB0F
FB27
FABA
FA80
FAD0
FB29
FB14
FAE0
FB0B
FB6E
FB89
FB58
FB47
FB71
FB83
FB4B
FB0A
FB04
FB21
FB1E
FAF6
FAEA
FB14
FB4A
FB59
FB4E
FB4E
FB64
FB87
FBAB
FBAD
FB71
FB26
FB1D
FB4C
FB4D
FB0D
FB0E
FB9B
FC29
FBFB
FB4C
FB26
FBD7
FC4C
FB9B
FACF
FC10
FFDB
03FB
05F5
05B1
0509
0535
05A8
0572
04BC
045F
049C
04EA
04E5
04CC
04E3
04FA
04CF
0496
049B
04C1
04C2
04B1
04D6
0520
053B
051E
0514
053D
0548
04E6
0450
0406
0432
0480
04A4
04AD
04BE
04C5
04B3
04A3
049B
047A
0454
0475
04D7
04EE
046C
03E5
041F
04E3
0527
0495
0442
0510
05DC
046A
0050
FBFE
FA1E
FAB5
FBA4
FB80
FADF
FAD2
FB44
FB5A
FADF
FA83
FABD
FB2F
FB56
FB43
FB4E
FB6A
FB52
FB0D
FADE
FAD7
FADF
FB02
FB53
FB9E
FB89
FB1A
FAC0
FACE
FB17
FB41
FB4B
FB78
FBC8
FBE1
FBA0
FB54
FB4A
FB6A
FB75
FB63
FB35
FADF
FA8F
FABA
FB70
FC00
FBC7
FB27
FB22
FBD0
FC04
FB0B
FA48
FBF5
003C
0489
0653
05C3
04EB
04F5
0536
04D4
042C
0428
04D1
055B
0554
0521
0532
0556
0537
04F7
04EE
050F
050B
04E4
04DA
04F4
04F9
04D1
04A6
0495
048D
048B
04AE
04FB
052F
0507
04B0
0492
04C3
04E2
04B1
046D
0462
0488
04BC
04FB
0522
04E2
0444
03EB
0450
04F8
04FA
0464
044F
052D
0589
0379
FF3C
FB70
FA3C
FB0D
FBC0
FB60
FAC4
FAD3
FB3C
FB35
FABB
FA6A
FA80
FA9D
FA8A
FA91
FAE2
FB1E
FAF1
FAA8
FAC7
FB36
FB72
FB4D
FB21
FB32
FB57
FB4A
FB0F
FADD
FAD4
FAE6
FB06
FB30
FB47
FB28
FAF0
FAEC
FB37
FB8F
FBB3
FBA6
FB7E
FB3D
FB0A
FB2F
FB9E
FBD2
FB82
FB27
FB5E
FBD2
FB80
FA5A
FA12
FC6F
00F1
04F2
0665
05CD
0512
051C
0550
050C
0499
0490
04E8
052C
052B
0518
050B
04E5
04B5
04CB
0531
0574
054A
050A
052A
057E
057D
0509
049F
04A8
0505
054E
0554
052E
04F6
04B8
0493
04AA
04DE
04E2
0499
0449
043A
046A
04B1
04F4
0506
04BA
043C
0417
0486
0506
04F9
0499
04BA
055F
051E
02A0
FE8C
FB41
FA5C
FB24
FBBC
FB5C
FABD
FAB1
FB14
FB4A
FB22
FAEC
FAE4
FAF7
FB06
FB0C
FB01
FAD2
FAA5
FAC7
FB37
FB7D
FB3D
FABF
FA9B
FAF4
FB60
FB7F
FB60
FB44
FB41
FB42
FB41
FB51
FB72
FB87
FB83
FB81
FBA0
FBCE
FBDE
FBB3
FB4E
FADA
FAAD
FAFE
FB8B
FBC6
FB8B
FB4E
FB66
FB66
FABA
F9DB
FA64
FD5D
01BD
0515
05F5
0522
0464
0489
050C
053B
0517
0509
053C
0580
059B
057A
052C
04DC
04C3
04F9
053A
052E
04E6
04CF
0518
055C
052B
04AD
046E
049F
04E5
04DF
04A2
0477
046C
0452
0426
0425
046C
04BB
04BD
0476
0440
045A
04B0
04FD
0510
04F6
04F4
0535
057D
0559
04C9
0478
0500
05D5
0563
029A
FE5E
FAF2
F9D3
FA70
FB1C
FAF5
FA7A
FA72
FADD
FB19
FAD5
FA6F
FA6C
FAD3
FB31
FB2A
FAD7
FA9F
FABF
FB1A
FB5A
FB50
FB20
FB12
FB3B
FB68
FB66
FB3E
FB0F
FAE8
FAC8
FAC8
FB08
FB79
FBD7
FBEA
FBB9
FB7D
FB62
FB61
FB59
FB33
FB00
FAF3
FB3A
FBAE
FBD7
FB70
FAEF
FB1F
FBFE
FC78
FBB3
FA80
FAE4
FDE4
0224
052C
05ED
057F
0563
05B9
05A0
04D4
042A
0466
053C
05C5
05AA
055B
054C
055E
053F
04FA
04D8
04EA
04F9
04E9
04E5
0505
051E
04FC
04B1
0480
0486
049E
04A6
04A6
04AC
04A7
048A
0477
0498
04CC
04BC
0460
0428
046F
04DE
04CB
0435
03FA
04AE
0570
0479
0124
FCFF
FA6D
FA44
FB26
FB55
FA98
FA0A
FA61
FB14
FB3D
FAD2
FA88
FAC3
FB20
FB2A
FAFB
FAFA
FB35
FB5E
FB51
FB43
FB60
FB82
FB74
FB48
FB3A
FB52
FB57
FB2A
FAF1
FADA
FADE
FAE4
FAEF
FB08
FB10
FAEF
FAD5
FB11
FB8D
FBC7
FB80
FB2E
FB72
FC12
FC1F
FB4C
FAD5
FC68
0029
042D
0648
0620
052C
04DB
0532
0552
04DF
0462
046C
04DA
051F
0505
04D1
04D3
0505
053B
055E
0562
0536
04DA
0480
0464
048A
04BB
04D6
04E5
04F9
0503
04FC
0502
0525
053B
0512
04D6
04EE
055E
0598
0535
049E
0498
0529
0576
04EE
043C
0478
0568
0549
02B5
FE6D
FAD0
F983
FA11
FAE7
FB1E
FB07
FB35
FB99
FBBF
FB7E
FB1E
FAEC
FAF5
FB26
FB69
FB94
FB7A
FB27
FAF3
FB1D
FB78
FB99
FB62
FB25
FB2A
FB54
FB59
FB37
FB26
FB2C
FB0C
FABB
FA9F
FB07
FB95
FB99
FB07
FA9D
FAE7
FB6D
FB54
FAAF
FA7F
FB3D
FBF6
FB80
FA67
FAC2
FDCC
022D
053F
05CE
0509
04BA
0545
05C6
05A8
054B
0532
0536
04F7
0495
0475
0493
048A
0442
0426
0476
04D4
04C5
046F
0462
04BF
0503
04D7
0492
04AB
0500
0514
04E0
04D8
0523
053F
04C8
042B
0425
04B7
0515
04CB
046A
04A5
0536
0537
0490
0447
0508
05C9
04A4
010E
FCC7
FA31
F9FE
FAE2
FB5B
FB34
FB26
FB81
FBC5
FB86
FB0E
FAEC
FB28
FB4E
FB27
FB02
FB2F
FB81
FB95
FB61
FB3B
FB4D
FB65
FB5B
FB53
FB77
FB9A
FB7F
FB41
FB37
FB6A
FB81
FB51
FB29
FB5C
FBA7
FB89
FB0E
FAD6
FB2A
FB90
FB88
FB59
FB91
FBED
FB95
FA8C
FA58
FC86
00A5
046A
05F7
0595
04E0
04D2
0511
04FC
04A5
0480
04A3
04B5
0487
044C
0446
046B
0492
04B3
04D7
04EF
04EE
04F4
0522
0557
054B
04F8
04B3
04BD
04E4
04CF
047E
0455
048E
04E6
04F1
04A9
0465
0456
0451
0436
0444
04B0
0528
050B
0458
03F5
04A1
05AF
0549
0262
FE21
FAED
FA14
FAC0
FB4B
FB18
FAC8
FAEC
FB3C
FB31
FAEB
FAF0
FB4A
FB75
FB2D
FADF
FB07
FB7E
FBC1
FBB0
FB95
FB8D
FB5C
FAED
FA9F
FAC6
FB1E
FB26
FAE1
FAD8
FB45
FBB8
FBB8
FB73
FB56
FB5A
FB24
FACA
FAD9
FB77
FBF6
FBBB
FB37
FB5F
FC31
FC6D
FB51
FA13
FAE3
FE68
02CF
0596
05F6
052D
04B7
04D3
04E0
049B
0473
04C4
053D
0553
04FD
04B6
04CA
04FE
04F7
04BF
04B8
050A
056E
0585
054E
0515
0509
0516
051A
051B
0521
051E
0506
04E9
04D9
04C3
0495
046C
047F
04BD
04CD
0491
046B
04BA
0531
0524
0495
0460
04F5
0547
03B0
FFFE
FC0C
F9FF
FA27
FB0A
FB4E
FB02
FAE5
FB1F
FB2A
FACE
FA80
FAB1
FB2E
FB75
FB60
FB38
FB39
FB43
FB26
FAEE
FAC4
FAB7
FABD
FAD4
FAF8
FB05
FAE0
FAAF
FAB1
FAEE
FB29
FB3A
FB43
FB6C
FB8D
FB5E
FAF7
FACF
FB20
FB80
FB5F
FAD7
FA9F
FB10
FB92
FB61
FAC3
FB1F
FD88
015B
04A8
0601
05AD
050C
04FC
0544
0557
0533
0538
0572
0575
0505
0476
0447
0482
04C3
04D6
04E4
0512
052A
04EF
0483
044C
046D
04B3
04E4
0502
051D
0529
051D
0519
0538
0547
04FB
0473
042F
0462
04A6
0491
045A
0484
04FB
0514
0493
043C
04CF
05A1
04EB
01D0
FDA9
FACF
FA3E
FAE2
FB27
FAB7
FA5E
FAAA
FB35
FB58
FB0E
FAD2
FAE6
FB12
FB1C
FB23
FB54
FB90
FB8B
FB40
FB01
FB11
FB54
FB7D
FB6D
FB48
FB34
FB2C
FB21
FB20
FB39
FB61
FB79
FB79
FB6A
FB46
FB05
FACF
FAE5
FB4D
FBAA
FBA8
FB7C
FBA0
FC0B
FC08
FB37
FA90
FBC0
FF45
0380
061B
063F
0523
0474
04A2
04F6
04E0
049F
0499
04B2
0492
0449
0440
0496
04E4
04D1
048B
047B
04B9
04F6
04FB
04E6
04E8
04F5
04EB
04CF
04CB
04E8
0506
0513
051B
051E
0505
04D2
04B3
04BE
04B8
0465
03F2
03E0
044F
04B6
0496
0449
0499
0579
058A
036D
FF84
FBE1
FA53
FAB7
FB7D
FB7D
FAF8
FABE
FB00
FB3A
FB1E
FAF6
FB1F
FB73
FB8E
FB5D
FB31
FB38
FB4D
FB46
FB3A
FB52
FB6D
FB4F
FAFC
FAC8
FAE1
FB13
FB1A
FB01
FAFD
FB1A
FB33
FB41
FB63
FB96
FB95
FB45
FAFB
FB12
FB58
FB3E
FABB
FA7F
FB04
FBAF
FB82
FAB0
FAE6
FD83
01C0
052C
0625
0553
0496
04D8
056A
055D
04C1
0457
0472
04AF
04B1
049C
04B6
04E3
04DE
04BA
04D1
052E
0568
0530
04BF
048D
04B5
04EA
0500
051C
0553
056C
0533
04DF
04D5
0516
053D
0512
04DA
04E2
0502
04E2
049E
04A7
0507
052D
04C8
046D
04C9
0556
0475
0149
FD12
FA2E
F9C0
FAC4
FB76
FB45
FAEA
FB14
FB86
FBA3
FB50
FAF5
FADA
FAE8
FAF9
FB22
FB6B
FB9D
FB82
FB36
FB03
FAF3
FACC
FA81
FA5A
FA90
FAEB
FB00
FAC5
FA9C
FACA
FB18
FB23
FAE5
FAB1
FABA
FAEA
FB1F
FB60
FBA5
FBAE
FB61
FB1E
FB5E
FBEA
FBED
FB21
FAAA
FC23
FFBE
03B3
05E2
05DF
0501
04AB
04F3
0524
04EB
04A2
0496
04A1
0499
04A9
04F8
0543
0529
04D0
04CC
054E
05CD
05BA
0547
051A
0567
05BA
05A8
055B
0534
0535
0518
04D7
04BA
04CF
04C3
046E
0425
044B
04A9
04C1
0490
0498
0500
052D
04A7
0406
0451
0557
0557
02D8
FE9A
FB15
F9F7
FAA3
FB4C
FB14
FA94
FA98
FB02
FB31
FB00
FAD7
FAEA
FAEB
FA9F
FA5D
FA9B
FB39
FB99
FB64
FAE6
FA93
FA7D
FA6E
FA65
FA8E
FADE
FB02
FAD6
FAA5
FAC3
FB12
FB37
FB30
FB51
FBAA
FBD7
FBA0
FB6F
FBBE
FC3C
FC19
FB3E
FAA3
FB11
FBEB
FBF6
FB45
FB95
FE3C
023D
0520
0599
04B8
0458
04FB
05AE
059E
050E
04A7
048B
047E
048B
04FB
05AF
0617
05E7
0578
054A
0564
056E
054A
0524
0509
04C7
0460
0439
0499
051B
051F
04A2
044D
048A
04FD
0515
04E2
04E9
0538
0535
0491
03E5
03FB
04A7
04F5
048A
0437
04BE
0559
0447
00EF
FCE6
FA6E
FA31
FAE2
FB08
FA8A
FA46
FAA9
FB3B
FB70
FB54
FB30
FB05
FAB1
FA5E
FA6C
FADC
FB44
FB60
FB64
FB8E
FBAF
FB6F
FAF0
FAB5
FAE7
FB10
FAD1
FA85
FABD
FB6C
FBEE
FBF4
FBD9
FBED
FBE1
FB54
FAB0
FAC1
FB6B
FB8F
FAB0
FA2A
FBEB
FFFA
0404
05BC
0537
0471
04C7
05A4
05CD
0523
049C
04D3
0559
0580
053D
04FB
04E4
04C8
0497
0487
04AB
04C4
04A2
047B
0495
04CF
04C3
0469
0431
0468
04CD
04F1
04D5
04CF
04F7
04FE
04C6
04A8
04EE
053A
04FE
046A
0451
04D8
04BA
0284
FE87
FAF6
F9B9
FA81
FB69
FB43
FAA0
FA9D
FB40
FB9D
FB3A
FAAC
FAAD
FB20
FB5C
FB24
FAE0
FAED
FB2B
FB4F
FB54
FB5C
FB57
FB22
FAE0
FAEE
FB59
FBBA
FBB5
FB73
FB52
FB5F
FB5B
FB35
FB27
FB44
FB4D
FB1B
FAF1
FB10
FB25
FAAE
FA13
FAC6
FDBE
020D
056F
067D
05D7
051C
050A
051E
04CB
0463
048B
0538
05BA
05AA
055C
054C
0576
057D
0541
0502
04F0
04E2
04A0
0441
040D
041C
044B
0471
048B
049C
04A2
04A5
04BD
04E0
04D1
047B
042F
0452
04C8
04FC
04AC
0465
04B8
0524
0446
016F
FDC1
FB38
FAAB
FB27
FB4D
FAE1
FAA2
FAF0
FB41
FAFF
FA6E
FA45
FAAB
FB04
FAD2
FA58
FA2F
FA78
FAD2
FAF0
FAEF
FB02
FB23
FB2E
FB25
FB2C
FB51
FB86
FBBD
FBE8
FBD3
FB5C
FAC8
FAA4
FB18
FB8E
FB5F
FABF
FA86
FB09
FB8A
FB4E
FAF3
FC0F
FF44
0328
058E
05BB
04DF
047C
04CD
050E
04D5
0492
04C6
0544
0589
0579
0567
057C
057D
0540
04FF
0506
053A
053E
04F1
0496
0474
0485
04A4
04C9
04ED
04ED
04B7
0488
04AE
050C
051E
04B7
045E
04A7
0553
058E
0520
04CF
052F
0570
03F9
0063
FC57
FA03
F9F3
FAD1
FB2A
FAE4
FACB
FB36
FBAA
FBAF
FB63
FB1A
FAD5
FA71
FA21
FA4D
FAED
FB66
FB49
FAD9
FAAD
FAE5
FB21
FB19
FAF6
FAFB
FB1B
FB24
FB1D
FB33
FB56
FB4C
FB1A
FB1A
FB6B
FBA6
FB66
FAF0
FADE
FB32
FB38
FAB3
FAB1
FC94
0047
03E7
059D
056A
04C8
04C1
0501
04C9
0437
0412
0499
052B
052E
04D8
04BF
04F4
04FF
04AB
045A
0474
04D6
050B
04F3
04D5
04E3
04FA
04F2
04E8
0506
052D
0520
04E4
04BC
04C5
04CD
04B5
04A4
04B6
04B6
0472
044A
04D1
05B8
0589
0312
FF02
FB9A
FA7C
FB27
FBD5
FB94
FB00
FAFD
FB67
FB71
FAE4
FA70
FAA9
FB3A
FB6F
FB29
FAF3
FB2C
FB8F
FBA6
FB6C
FB3A
FB40
FB57
FB57
FB4A
FB42
FB2A
FAF4
FAC1
FABD
FAE3
FB07
FB23
FB52
FB82
FB73
FB22
FAF0
FB21
FB57
FB02
FA75
FB09
FDB8
01B3
04E1
05DE
0541
0499
04A4
04DC
04A3
0440
045C
04F5
055B
0526
04BD
04B2
04F5
0507
04BF
047F
049D
04E4
04E8
049D
045E
046F
04B3
04E4
04EC
04DC
04C7
04BD
04CB
04E8
04E7
04AD
0471
047F
04C3
04D3
048E
046D
04DB
0543
044F
0165
FDA2
FAF7
FA4C
FAD9
FB51
FB40
FB16
FB22
FB1C
FAC0
FA61
FA81
FB12
FB7E
FB6B
FB1F
FB0F
FB44
FB6F
FB66
FB54
FB5B
FB61
FB46
FB18
FAFE
FAF6
FAED
FAEC
FB0E
FB48
FB6C
FB75
FB8F
FBC0
FBBF
FB5F
FB00
FB25
FB9A
FB7C
FA7E
F9D5
FB42
FF0E
035C
05DF
0602
0520
04B0
04DA
04E8
0494
0457
0496
0506
052D
050C
0507
053D
0563
053E
04FE
04EA
04F7
04E5
04B1
0494
04A3
04B5
04AE
04B5
04F2
053D
054A
0516
04EA
04E7
04DC
04A4
0472
047F
04A2
048B
0468
04CA
05A7
05CC
03E2
000F
FC34
FA39
FA4D
FB12
FB4B
FAFC
FAD5
FB1A
FB67
FB66
FB39
FB1D
FB09
FADA
FAAF
FACB
FB23
FB59
FB39
FAF4
FAD6
FAE0
FADE
FACC
FAD9
FB0C
FB29
FB09
FAE5
FB00
FB40
FB4F
FB1C
FAF8
FB22
FB67
FB79
FB6A
FB7A
FB88
FB2B
FA8F
FAD1
FCFD
00AB
0410
05A7
058E
050A
04FB
0529
0514
04D5
04E6
054B
057E
0537
04D3
04CC
0506
0504
04A0
0448
0466
04D5
0527
0532
0521
0514
04F7
04C5
04AD
04CE
04FA
04F2
04C2
04B7
04E4
050F
050C
04FE
050C
050D
04D4
04A7
04F6
0576
04F8
028B
FECA
FB88
FA1D
FA3D
FAA6
FAA7
FA89
FAB5
FB00
FB09
FAE7
FAFF
FB54
FB68
FAF3
FA61
FA55
FAD4
FB49
FB42
FAF1
FAD5
FB1F
FB92
FBDB
FBD2
FB82
FB21
FAFB
FB33
FB88
FB82
FB09
FA91
FA90
FAE0
FB04
FAEC
FB0B
FB8B
FBCE
FB45
FA94
FB54
FE49
0235
04ED
0574
04C2
0461
04CB
0557
0564
0517
04E8
04F3
04FE
04FC
0513
0547
055D
052B
04D9
04A8
04A9
04BF
04D2
04E4
04EE
04ED
04FB
0535
0570
054C
04BF
044D
047D
0518
0553
04D8
043B
043C
04BE
04F7
04A3
0478
0503
0578
0445
00F0
FCF8
FA7D
FA37
FB07
FB7D
FB41
FAF3
FB0A
FB50
FB5D
FB29
FAF3
FAD5
FABD
FAAD
FAC3
FAF7
FB13
FAF7
FAD1
FADE
FB1A
FB48
FB48
FB2B
FB06
FAD6
FAA9
FAB7
FB1D
FB9C
FBCA
FB94
FB53
FB47
FB4A
FB23
FB04
FB43
FBA7
FB7C
FAA8
FA5D
FC20
FFEC
03CE
05A8
0547
044E
043C
04F6
0568
051E
04B4
04CF
053D
055E
050B
04B1
04A7
04CA
04D5
04D2
04EE
051E
0526
04F9
04D2
04DA
04F6
04FF
04FD
04FE
04EC
04B6
048B
04AC
04F8
0502
04A8
045D
0489
04DE
04C1
0455
0478
0562
05C3
03E1
FFC2
FB8F
F989
F9DF
FAE7
FB3A
FAFF
FB0A
FB7D
FBB6
FB64
FAF3
FADA
FAF4
FAE1
FAAA
FAB2
FB07
FB43
FB21
FAE6
FAF2
FB2D
FB38
FB00
FADB
FB03
FB4B
FB71
FB74
FB75
FB61
FB19
FACB
FACF
FB24
FB52
FB1E
FAEC
FB2E
FB97
FB74
FAEB
FB51
FDC7
01A3
04CB
05CB
052E
0490
04BB
0527
051F
04C9
04C1
051F
0563
053A
04F2
04F9
0539
0544
04FB
04B0
04AF
04E4
0507
0504
04F6
04F2
04EE
04E3
04D5
04B5
046E
0419
0405
045D
04E2
0532
053D
053D
0547
0522
04C5
049C
0500
0557
0450
0151
FD7F
FAE0
FA6D
FB3B
FBB7
FB58
FAD7
FAE3
FB39
FB2E
FAB9
FA77
FAC6
FB41
FB5B
FB1B
FAFE
FB3B
FB7A
FB67
FB1F
FAFE
FB17
FB33
FB38
FB43
FB63
FB66
FB30
FAFC
FB1B
FB78
FBAC
FB82
FB3B
FB29
FB46
FB62
FB7A
FB9C
FB8B
FB0A
FA99
FB82
FE80
0282
054F
05B3
04B0
042D
04CF
0596
0584
04E7
04B4
0515
0547
04DF
046A
0495
0520
0543
04D6
0480
04BA
0518
04F9
0477
0446
04AA
0521
0522
04CD
049A
0498
0482
044F
0443
0467
0469
043C
0464
051B
0569
03C7
0006
FBFE
F9E7
FA22
FB20
FB67
FB02
FADC
FB3A
FB7B
FB38
FAE1
FAFD
FB56
FB4C
FAD3
FA84
FABF
FB28
FB46
FB31
FB53
FBA6
FBAD
FB3B
FACA
FADD
FB4A
FB83
FB62
FB48
FB6D
FB87
FB58
FB34
FB88
FC04
FBE0
FB22
FB21
FD3D
0119
04A9
062C
05CD
0518
051C
0590
05B1
055F
051E
052E
0544
0514
04CB
04BA
04D3
04C8
048F
0478
04AF
04F8
0505
04E6
04E1
04FB
04F1
04B7
049A
04C4
04DE
048B
0412
042B
04F4
05A2
057A
04DA
04B2
04F3
0437
0164
FD58
FA53
F9A4
FA6C
FAF2
FA9D
FA34
FA62
FAC2
FAAD
FA50
FA67
FB1A
FBB1
FB96
FB1F
FAF9
FB33
FB4B
FB18
FB09
FB6D
FBDD
FBC5
FB3D
FAE7
FB0F
FB57
FB5B
FB3A
FB39
FB36
FAF2
FAB3
FB08
FBC9
FBFE
FB30
FA88
FBDD
FF83
0396
05D5
05E2
0535
051C
0578
057D
051A
04F2
0546
058E
0551
04E6
04F8
0583
05D9
058D
04F7
04AC
04BB
04C7
04A3
0485
0498
04BC
04C7
04CC
04E7
04EA
049E
043A
043F
04BB
050B
04A8
0400
0406
04D3
0511
0342
FF8E
FBDA
FA05
FA31
FB02
FB46
FAFC
FACF
FAFE
FB2F
FB19
FAF1
FB07
FB46
FB56
FB28
FB03
FB0F
FB19
FAEC
FABB
FAE4
FB60
FBAF
FB71
FAE5
FA9D
FADA
FB55
FBAD
FBBC
FB8D
FB36
FAF1
FB16
FBA1
FBF2
FB73
FAA6
FB22
FDF7
022A
0556
05FA
04EE
0434
04B6
058F
058F
04C7
0440
0487
050D
050C
048A
0425
0439
048F
04D0
04ED
0500
0508
04F8
04E6
04EF
0501
04F3
04D5
04DA
0500
04FC
04B0
046E
0491
04DC
04C2
0445
042A
04E3
0591
0494
015C
FD4F
FA8C
F9F1
FA8C
FAF2
FAB4
FA68
FA96
FB19
FB77
FB85
FB73
FB6C
FB6C
FB72
FB8A
FBAE
FBAF
FB71
FB21
FB08
FB36
FB6C
FB6E
FB43
FB19
FB04
FAFC
FB06
FB34
FB71
FB75
FB28
FADC
FAF4
FB49
FB41
FABB
FAAD
FC6E
0019
0406
062B
060F
0511
04BB
0534
0586
0520
0485
046F
04C9
04EC
04A4
046E
04A6
04F4
04D1
045B
0429
0469
049E
0462
040A
0435
04DD
0552
0521
0499
044E
045F
048B
04B7
04F8
0526
04F3
0483
047F
050F
0512
0309
FF04
FB14
F960
F9FC
FB19
FB38
FA9A
FA66
FAF2
FB83
FB80
FB3A
FB4B
FBA3
FBBC
FB71
FB32
FB54
FB97
FB94
FB57
FB4A
FB91
FBDB
FBD6
FB96
FB62
FB58
FB67
FB7F
FB90
FB78
FB2C
FAF6
FB34
FBBF
FBDA
FB29
FA88
FB82
FEA6
02A7
0569
05FD
0547
04C1
04F8
0566
0568
0504
04A2
0477
046B
0469
0478
048B
047C
0448
042C
0458
04A0
04AA
0468
042E
0444
0488
04AC
049D
048F
0497
0489
0456
0444
0489
04D9
04B4
0433
041D
04D5
0565
042F
00CC
FCD5
FA7B
FA5F
FB34
FB79
FB05
FAB2
FAF7
FB5F
FB6B
FB50
FB83
FBE7
FBEC
FB77
FB1B
FB46
FB9E
FB8D
FB25
FB08
FB76
FBE5
FBCA
FB60
FB49
FBA4
FBEC
FBD0
FBA0
FBB6
FBD7
FB9B
FB38
FB44
FBB6
FBBB
FAFF
FAA7
FC5D
0036
042E
061D
05D4
04E9
04B2
0503
0500
047E
0419
043E
04A5
04E4
04FD
052A
0550
051B
0496
0432
043F
0487
04A4
047F
044F
043A
0437
0446
047E
04C8
04D2
0483
043A
0460
04C1
04B6
041C
03B4
043B
052E
04EE
026C
FE79
FB2B
F9F8
FA8F
FB81
FBC5
FB65
FAF5
FAD1
FAE9
FB14
FB3F
FB5F
FB63
FB51
FB50
FB72
FB90
FB79
FB39
FB15
FB35
FB6F
FB89
FB79
FB67
FB63
FB5F
FB5C
FB81
FBCA
FBE6
FB96
FB2B
FB37
FBC2
FC06
FB73
FAC4
FB98
FEA4
0299
053D
05A1
04D3
046B
04CD
0530
04FC
0496
049F
050A
0546
051A
04E0
04D8
04C7
0470
0411
0412
0466
04A2
04A5
04C6
052E
056A
050A
045D
041F
0477
04BA
0476
041F
0454
04CC
04B4
0411
03F6
04E9
0599
0410
0023
FC0A
FA1A
FA73
FB50
FB5C
FAE3
FACC
FB2E
FB66
FB3B
FB22
FB69
FBAE
FB7F
FB17
FB0D
FB6E
FBA6
FB58
FAE6
FADC
FB36
FB7E
FB77
FB56
FB46
FB21
FAD6
FABE
FB2C
FBCB
FBE1
FB5A
FB05
FB7F
FC30
FBF5
FAE3
FABA
FD10
014F
0502
064B
059D
04CE
04E4
0553
0541
04C9
049D
04E6
050F
04B5
0442
0448
04AF
04E7
04BE
049F
04D3
0509
04CD
0448
041E
048F
0524
054B
0508
04C3
04A8
0496
0489
04B2
04FC
04ED
0454
03D5
0431
04FF
04A2
0204
FE19
FB1D
FA4A
FACC
FB17
FABC
FA78
FAC7
FB2F
FB15
FAB8
FAC0
FB31
FB66
FB21
FAF2
FB54
FBDF
FBD2
FB34
FACE
FB0E
FB7C
FB7B
FB2B
FB13
FB48
FB63
FB4E
FB77
FBF9
FC33
FBAB
FAFC
FB2A
FC13
FC5B
FB4B
FA30
FB30
FEC4
02FE
057C
05B9
050D
04D4
052C
0578
0565
0521
04E5
04B6
0499
04AB
04E5
0507
04EF
04D7
0504
0551
054D
04E0
047C
048B
04D5
04CE
0462
0421
0473
04F3
04E7
044D
03FB
0478
0529
050E
0435
03CC
0481
0534
03FB
006C
FC60
FA2A
FA49
FB45
FB8D
FB07
FA98
FAC2
FB2A
FB49
FB18
FAE1
FAC8
FAC5
FAD8
FB10
FB4C
FB52
FB22
FB05
FB2F
FB6D
FB6F
FB40
FB33
FB5E
FB75
FB43
FB04
FB14
FB5B
FB66
FB20
FB07
FB73
FBE1
FB85
FA9E
FAB2
FD06
00EF
043C
0562
04E7
047A
04F3
05B6
05E2
057F
0534
0541
0546
050B
04E0
0510
055A
0549
04E1
0491
048C
0495
047E
047F
04CC
052B
0536
04F5
04CF
04E1
04CF
0471
0441
04AF
0550
0545
0488
042B
04F7
0608
0567
0234
FDCD
FA93
F9B7
FA74
FB3F
FB4E
FADE
FA80
FA6F
FA97
FAD3
FB07
FB19
FAFD
FACF
FABF
FAD9
FAFB
FB0C
FB1A
FB3D
FB61
FB51
FB0A
FACC
FAD8
FB17
FB3E
FB2C
FB1A
FB39
FB64
FB58
FB2C
FB3A
FB82
FB7A
FAE1
FA87
FBD3
FF2A
0321
05A3
05E7
0505
0494
0507
05A2
05B2
0554
050B
0501
0500
04EB
04EA
050F
0529
050F
04E5
04EB
051E
0536
0511
04D6
04BA
04BB
04C1
04CB
04E1
04E4
04B5
0487
04B8
0540
0581
0508
044E
044E
0514
0536
032B
FF2F
FB56
F994
F9EF
FAE8
FB4C
FB23
FB03
FB0C
FAF6
FAC4
FACB
FB15
FB36
FAF1
FAA6
FACD
FB43
FB7C
FB4E
FB1D
FB2E
FB44
FB11
FAC7
FAD5
FB2F
FB55
FB1B
FAFB
FB4E
FBAE
FB83
FAFB
FAE6
FB7D
FBEE
FB73
FAA3
FB1C
FDBE
0192
04AA
05EA
05B9
052E
04F3
04FF
0504
04DD
04A5
0488
0498
04C8
0505
053B
0559
054D
0520
04F3
04EA
04F7
04EA
04BA
04A8
04F0
0558
0564
04FB
0496
0496
04B8
0482
041A
042E
04D2
04E0
0307
FF71
FBEE
FA3C
FA68
FB1D
FB44
FAF6
FADB
FB24
FB6B
FB5C
FB24
FB21
FB61
FB95
FB79
FB21
FADB
FADF
FB27
FB79
FB99
FB74
FB2D
FAF4
FAE9
FB11
FB4C
FB69
FB4E
FB24
FB2D
FB68
FB73
FB1C
FAFE
FC3B
FF41
02F8
0580
05F9
0542
04DD
0547
05BB
057B
04C6
046B
04AB
0506
0506
04D3
04C9
04D8
04AB
044A
042B
0485
04F1
04EE
0499
0486
04E0
0524
04E4
0474
047E
0502
0541
04D0
0450
049A
0552
04E6
0244
FE49
FB1F
FA22
FAC0
FB63
FB36
FAAA
FA81
FAD2
FB1A
FB0C
FAE4
FAF9
FB42
FB6C
FB4D
FB18
FB0F
FB39
FB64
FB74
FB7F
FBA3
FBD6
FBF1
FBE4
FBC1
FB90
FB46
FAF7
FAE8
FB3C
FB93
FB5C
FAB7
FAD3
FCE9
00B3
0441
05B7
051D
0424
043B
0522
05A3
0533
047A
044C
04A0
04E0
04D3
04D2
0517
0559
053C
04DA
049F
04A7
04A2
045B
0411
0427
048C
04CC
04B0
047C
047D
048E
045B
0409
0430
04FC
0573
0425
00BC
FCB4
FA27
F9EE
FB07
FBE0
FBDA
FB72
FB45
FB5B
FB69
FB60
FB60
FB5E
FB2B
FAE0
FAE5
FB59
FBCA
FBBC
FB56
FB29
FB6C
FBAD
FB78
FAF9
FAC4
FB07
FB57
FB57
FB3E
FB76
FBDC
FBD0
FB1F
FAA1
FBA8
FEA3
0273
0537
05E8
0525
0462
046A
04D7
04F0
04AA
0491
04E6
053A
0511
049B
046B
049B
04B3
046E
0435
0476
04EE
04F8
0483
0432
0474
04E9
04F1
049E
0490
04F5
0533
04D2
0453
0489
0537
04EA
027F
FE9C
FB4A
FA1A
FAC8
FBBE
FBC8
FB13
FA97
FAD4
FB5F
FB94
FB63
FB3A
FB58
FB79
FB53
FB18
FB2B
FB84
FBB1
FB8A
FB78
FBCD
FC2A
FBF3
FB3A
FABA
FADD
FB2C
FB0D
FAB5
FADD
FB88
FBD0
FB42
FAF2
FC86
0026
03FC
05F6
05C2
04CC
0470
04B8
04E0
04A3
0481
04DB
054A
0525
0476
03FA
0436
04D1
0509
04A3
0423
040A
043E
0457
045E
04AD
0539
056B
04F4
0467
0481
0519
053E
0496
040D
0491
0571
04B9
0175
FD1D
FA3C
F9E2
FADD
FB69
FB17
FABA
FAFB
FB83
FBA8
FB62
FB3A
FB74
FBB4
FB95
FB3A
FB1F
FB65
FBAB
FB97
FB4E
FB39
FB6F
FB96
FB6F
FB3A
FB4F
FB8A
FB71
FAF9
FAB4
FB02
FB68
FB30
FAAC
FB49
FE07
020E
0537
0618
053E
044D
0443
04CF
052B
0510
04C7
049D
049A
04A3
04B5
04D3
04E7
04D7
04AB
048F
0499
04A5
0486
0451
044F
04A1
0501
050E
04CE
04B4
0503
0554
051D
048F
047D
0514
0525
033C
FF70
FBB3
F9FE
FA72
FB85
FBD4
FB63
FB09
FB28
FB64
FB57
FB18
FAF3
FB03
FB27
FB48
FB64
FB77
FB6C
FB3D
FB11
FB1A
FB57
FB8F
FB8B
FB57
FB23
FB0C
FAFA
FADD
FAE2
FB3E
FBB9
FBA9
FADC
FA5F
FBC0
FF49
034D
05A9
05D3
0514
04D0
0517
0520
04B0
0456
046D
0497
046F
043C
047B
0505
0538
04E4
0487
0494
04D9
04E6
04B8
04B5
04FB
052C
04FC
04A8
04A5
04FB
053E
051F
04CE
04B9
0504
0525
0426
017E
FDDE
FAF1
F9F5
FAA0
FB7C
FB78
FAD6
FA8D
FAF7
FB86
FBA7
FB79
FB66
FB7A
FB75
FB4E
FB3C
FB4E
FB54
FB3A
FB2F
FB52
FB75
FB5D
FB24
FB1E
FB4A
FB45
FADC
FA78
FAA0
FB35
FB84
FB28
FAB2
FB50
FDAC
0133
045D
05E2
05BA
04F9
04B4
050C
055E
0530
04C1
0496
04BE
04D3
04A1
046E
0480
04AC
04A7
0482
0491
04DB
0501
04CA
047F
048C
04E3
050C
04D7
04A3
04CC
051C
0515
04BC
04A4
04FE
04EC
033C
FFD7
FC3B
FA39
FA42
FB32
FBA9
FB67
FB1F
FB44
FB7D
FB51
FAE9
FAD3
FB33
FB91
FB7A
FB10
FAD0
FAEF
FB3B
FB7A
FBA5
FBBA
FB9C
FB4D
FB12
FB24
FB53
FB3C
FADF
FAB7
FB1C
FBB6
FBCA
FB28
FAB9
FBD8
FEEB
02BF
0568
05E8
0503
0450
049C
0548
055C
04CA
045E
048B
04E4
04DE
049E
04A1
04E3
04EC
04A2
0484
04E0
053D
04FC
045A
042E
04B6
0536
050D
049B
0495
04DF
04C5
0436
041A
04FB
05E6
0527
0230
FE59
FB91
FA97
FAB1
FAD1
FA9B
FA5F
FA78
FAE1
FB4C
FB76
FB6C
FB67
FB78
FB72
FB3B
FB02
FB03
FB2D
FB37
FB13
FB14
FB6D
FBCB
FBB3
FB3F
FB0A
FB4E
FB88
FB41
FAD6
FAF0
FB6C
FB68
FAB8
FAA5
FCB3
00A6
0461
05F6
0585
04BA
04C0
053B
0542
04BE
046B
04B8
053D
055A
050F
04E0
0505
0522
04D3
044F
041E
0465
04BF
04D2
04C1
04D6
0502
04F2
04A3
047C
04B9
04FE
04D7
0480
04AF
056F
0591
03BF
0012
FC47
FA33
FA2C
FB09
FB85
FB5A
FB1A
FB32
FB70
FB66
FB0B
FABE
FACB
FB13
FB44
FB3F
FB30
FB3E
FB51
FB45
FB38
FB5F
FBA6
FBAD
FB53
FAF6
FAFB
FB3A
FB3C
FAF5
FAE6
FB53
FBAE
FB50
FAAC
FB41
FDF4
01CB
04B8
0597
0512
0493
04B9
0515
0522
04F8
04F8
0528
0533
04FA
04C9
04E3
051E
0516
04BC
046E
0480
04CE
04F3
04C3
0482
0475
0489
0480
0461
0479
04D4
050E
04E2
04AA
04FA
059D
0556
0311
FF44
FBD2
FA62
FADC
FBCA
FBEB
FB45
FAAB
FAA4
FAF5
FB28
FB1C
FB0E
FB28
FB4D
FB52
FB37
FB1A
FB07
FAFD
FB09
FB3C
FB7D
FB8D
FB5C
FB33
FB5C
FBB2
FBB8
FB49
FAE3
FB0A
FB72
FB51
FA96
FA75
FC3B
FFB9
0336
050F
0530
04C2
04BA
050A
0528
04F3
04BE
04C5
04F1
0517
0528
051C
04DD
0476
0431
045A
04DC
0546
0539
04D4
0486
0485
0496
0472
0434
0449
04CE
054B
0532
04AD
0492
0548
05E7
04D8
0192
FD7A
FAB6
FA36
FB0B
FBA9
FB7A
FB06
FAEE
FB1C
FB1E
FAE8
FADE
FB34
FB96
FB96
FB39
FAF6
FB1E
FB80
FBAB
FB7D
FB3D
FB34
FB4B
FB45
FB2F
FB46
FB80
FB78
FB06
FA9B
FABC
FB36
FB51
FB03
FB76
FDCF
0184
048C
0570
04CA
0449
04AE
053F
052B
04BB
04BC
0539
056E
04EF
0449
043B
04B4
0507
04EB
04C5
04EF
0527
04FE
0487
0447
047B
04C8
04CE
04AF
04D1
0528
052F
04AA
0426
0456
0500
04E2
02F2
FF93
FC61
FAB9
FA98
FB00
FB2B
FB1E
FB2B
FB47
FB23
FAC0
FA8A
FACD
FB4A
FB81
FB4A
FB01
FB08
FB50
FB75
FB48
FB06
FAFB
FB14
FB0C
FAE0
FAD9
FB1E
FB66
FB5F
FB39
FB70
FBF4
FBFA
FB1B
FA60
FB93
FF22
034B
05BC
05DB
0505
04B2
04F9
0510
04BA
047F
04B9
0505
04F2
04AB
049D
04CD
04F4
0501
051C
053E
0535
0508
04FF
052F
0548
0509
04B7
04AB
04BC
0484
0440
049D
056D
0535
02C4
FED6
FB8A
FA3E
FA78
FAF4
FB20
FB34
FB52
FB45
FB11
FB1A
FB76
FBA6
FB5A
FAFD
FB1A
FB80
FB91
FB35
FAEE
FAFF
FB0C
FACD
FA99
FADD
FB50
FB53
FB02
FB23
FBD9
FC1F
FB40
FA56
FB66
FEEE
0308
055D
0573
04B6
0485
04E0
0510
04E2
04BA
04D2
04E4
04BA
0485
048C
04C6
04F2
04F7
04EE
04E4
04D2
04C3
04D5
04FC
04FC
04C3
0495
04AA
04D0
04B9
0492
04DF
0577
051D
02B1
FEC9
FB83
FA79
FB32
FBF0
FBBF
FB27
FB08
FB5C
FB82
FB48
FB14
FB27
FB37
FB01
FABF
FABE
FAE8
FB04
FB1F
FB60
FB9D
FB94
FB64
FB67
FB90
FB6D
FAF4
FAD0
FB5F
FBD0
FB2F
FA42
FB3A
FEF3
0365
05AB
053D
0420
041E
04E1
0514
048E
0454
04DE
0565
0537
04B9
04A8
04F2
0511
04F4
04EF
04F8
04BE
0464
0470
04E8
051A
04A4
042A
0466
04ED
04BC
03F4
03EE
050F
058C
0369
FF30
FBA1
FAA0
FB61
FBEA
FB86
FB05
FB15
FB4F
FB1E
FAC0
FACA
FB2E
FB65
FB4A
FB38
FB60
FB84
FB73
FB5C
FB68
FB6C
FB3D
FB15
FB42
FB95
FB8D
FB2E
FB1A
FB91
FBDA
FB3D
FA77
FB58
FE9D
02BA
0542
056A
0496
0473
0521
0595
0543
04BB
04A9
04E7
04E5
0491
0460
0489
04BF
04B8
0497
0493
04A0
04A7
04CB
051D
054C
0503
0483
0463
04B3
04D6
048B
0477
0513
054F
036C
FF63
FB8C
FA22
FAD5
FB8A
FB23
FA7C
FAA9
FB55
FB76
FB05
FAED
FB7B
FBDE
FB84
FB03
FB1F
FB91
FB9A
FB3B
FB12
FB42
FB46
FAF6
FADD
FB4E
FBBA
FB87
FB1B
FB39
FB9D
FB51
FA98
FB53
FEA2
02EA
0565
0548
0452
0449
04FC
0537
04C9
0496
04FA
053B
04CC
0441
0461
04EC
0511
04B3
046E
0495
04D8
04EF
0500
0524
0514
04B1
0470
04BD
0528
04E6
042F
0436
0544
05AA
0381
FF38
FB6D
FA21
FACC
FB82
FB64
FB1E
FB62
FBC7
FB97
FB03
FAD5
FB41
FBA5
FB86
FB2E
FB23
FB61
FB7E
FB4E
FB07
FAD6
FAB2
FAA5
FAD8
FB37
FB63
FB42
FB42
FBA6
FBDC
FB37
FA58
FB1B
FE82
0304
05D0
05C9
0484
0420
04D5
054F
04D9
0433
0443
04CB
04FC
04B7
0495
04D3
04F8
04BA
0481
04B8
0514
0516
04CD
04A2
049E
047E
0451
0471
04CA
04D0
0478
0492
0580
05E4
03CC
FF58
FB3A
F9E0
FADC
FBDD
FBA9
FB14
FB2B
FB9D
FB84
FAEC
FAB7
FB27
FB84
FB46
FADB
FACE
FAEC
FACF
FAB6
FB16
FBB0
FBD9
FB86
FB5A
FB99
FBBF
FB72
FB39
FB9F
FBFB
FB43
FA0B
FA98
FE20
02D9
05B2
05AE
048F
044C
04E7
0532
04CB
0477
04BB
051E
050F
04D1
04ED
054D
056B
0532
050F
0529
0530
04EB
0494
046C
0458
042F
0425
0471
04C2
0497
0430
046F
0561
0581
0340
FF20
FB87
FA4B
FAEB
FB91
FB57
FAE4
FB03
FB77
FB84
FB13
FAAE
FA9D
FA9B
FA72
FA5F
FAA2
FB12
FB55
FB67
FB76
FB7E
FB52
FB14
FB28
FB89
FBB6
FB78
FB4F
FBA3
FBE6
FB4C
FA5F
FB02
FE48
02BF
05AA
05E4
04D7
046B
04DC
052C
04F4
04D6
053D
05A4
0576
04FF
04ED
053F
054C
04DD
048A
04C0
051B
0511
04BE
0497
04A0
0497
0497
04E8
0546
050A
0445
0409
04DD
056A
03A6
FF88
FB8C
FA0F
FAD2
FBC0
FB9F
FAFE
FAC0
FAD0
FAA7
FA5F
FA81
FB0B
FB60
FB42
FB25
FB54
FB69
FB08
FA9D
FAB9
FB2E
FB5E
FB36
FB33
FB69
FB4D
FAB3
FA60
FAF9
FBC7
FB93
FAB5
FB3D
FE72
02D3
0593
05AF
04AF
046D
0505
0565
051F
04D2
04F8
0532
050C
04C4
04D8
0524
0523
04CB
0495
04C3
0509
051F
0523
0543
0552
0516
04CF
04E4
052B
050B
048B
047B
051F
0536
0324
FF1C
FB52
F9CC
FA66
FB69
FBAA
FB6F
FB57
FB52
FB10
FAC8
FAE5
FB3F
FB41
FADD
FAB4
FB22
FBA6
FB93
FB09
FAB7
FADA
FB03
FAE9
FAD2
FAF3
FB02
FAD0
FAD1
FB60
FBDE
FB6C
FA97
FB59
FECA
0351
0608
05E6
04A2
044F
0503
0572
0516
04A8
04BC
04F0
04C7
0487
04B8
052D
0540
04E3
04BC
050D
053E
04DB
0459
0461
04D5
0514
0506
0511
052C
04D3
0414
03EB
04D4
056E
03AB
FF79
FB5A
F9B7
FA5D
FB3D
FB20
FAA2
FAB5
FB2D
FB4B
FAF7
FAC5
FAE8
FAF8
FAC3
FABF
FB3E
FBC9
FBBD
FB33
FAD0
FADE
FB1C
FB4F
FB86
FBAD
FB7A
FAFE
FADC
FB6F
FC03
FBAC
FAF0
FBA8
FEC5
02CA
0544
057C
04E7
0501
0592
0588
04C9
0459
04C8
0570
057D
0515
04DF
04F4
04E1
0490
0474
04C3
050D
04EA
0495
048F
04D2
04F3
04D8
04CB
04CD
047F
03FF
0419
0503
0558
0354
FF24
FB33
F9B9
FA77
FB60
FB31
FA8D
FA85
FB0A
FB52
FB29
FB0D
FB38
FB51
FB23
FB02
FB39
FB7D
FB63
FB0F
FB01
FB4B
FB72
FB3D
FB08
FB1D
FB43
FB47
FB77
FC00
FC3D
FB7B
FA76
FB28
FE88
02FC
05C8
05F7
0512
04E1
055B
055B
04A2
0425
047E
0512
0503
0470
0424
0473
04E6
050C
0502
0500
04EC
04AD
0484
04B2
04FC
04FA
04BC
04A4
04B1
0482
0424
0441
0504
052D
031F
FF06
FB29
F9AB
FA60
FB64
FB70
FAEC
FACD
FB2C
FB79
FB80
FB91
FBC3
FBB3
FB35
FAC5
FAE7
FB66
FBA3
FB72
FB36
FB33
FB41
FB2C
FB11
FB1D
FB3D
FB52
FB7F
FBD7
FBE7
FB39
FA6E
FB30
FE63
02BB
05BD
063B
0547
04AC
04ED
0535
04DE
0447
0422
0480
04F3
0534
0548
052C
04D5
047A
046A
049E
04BC
049B
0484
04B4
04EA
04C6
0469
0453
0493
04B2
048F
04B5
055A
0567
0364
FF6D
FB97
F9ED
FA64
FB42
FB48
FAD4
FACC
FB3B
FB7B
FB51
FB27
FB44
FB66
FB4A
FB24
FB41
FB77
FB5E
FAF9
FAC7
FB09
FB62
FB64
FB2E
FB2D
FB7B
FBCA
FBE3
FBCF
FB91
FB20
FADA
FBA5
FE1F
01A6
049B
05D0
0581
04DA
04AC
04EE
052C
0524
04E1
0493
0472
0497
04DD
04F9
04CD
049A
04AB
04EA
0504
04F2
0503
054A
055C
04E6
0442
0408
043E
045E
0445
0481
0543
0572
038A
FF9A
FBB8
FA04
FA89
FB85
FB91
FAE6
FA8B
FAE0
FB6C
FBB9
FBC6
FBA8
FB4A
FACA
FAA3
FB18
FBA8
FB97
FAEB
FA72
FAB2
FB40
FB60
FB11
FB01
FB7D
FBED
FB9F
FAE5
FAFD
FCD0
0005
034A
0563
05F8
058D
04F9
04C1
04E5
0514
050F
04DA
04A1
0481
0481
04A7
04E7
0513
04F7
04A9
047A
0493
04BA
04B8
04AD
04D9
051B
050D
04B2
04A5
0522
052E
0362
FFB0
FBF6
FA36
FA8C
FB4C
FB1F
FA5F
FA36
FAEC
FBA7
FBB3
FB50
FB1D
FB29
FB1A
FAE9
FAEA
FB29
FB41
FB08
FAEE
FB5A
FBE7
FBC5
FAE8
FA4D
FAB8
FB98
FBAB
FAC4
FA5B
FC0F
FFC8
03A7
05C9
05E8
0532
04DB
0512
0547
0515
04B5
049B
04E4
0539
053E
04F3
04A3
0489
04A0
04C3
04D6
04C7
0492
045E
0475
04E8
0551
0535
04B9
04A6
055E
05E2
0483
00D1
FC87
FA07
FA09
FB17
FB6A
FAC8
FA47
FA9A
FB40
FB70
FB26
FAEB
FAEF
FADD
FA96
FA76
FAC0
FB29
FB49
FB48
FB98
FC1A
FC14
FB43
FA77
FA9D
FB68
FB90
FA9E
F9EE
FB60
FF1E
032F
0563
0561
0499
0471
04F8
055C
0529
04B8
049A
04E0
052C
0537
0517
0505
050E
0518
0510
04F8
04D1
049C
0474
0483
04C8
04F2
04B5
044E
0466
0530
05B4
0474
0112
FD11
FA9D
FA78
FB6A
FBC2
FB24
FA81
FA9C
FB21
FB52
FB19
FAEF
FB04
FB05
FAC7
FAAE
FB0B
FB7A
FB59
FAC2
FA8B
FB1E
FBCB
FBBC
FB26
FB05
FB9F
FBFB
FB52
FA7F
FB65
FEB4
02D6
0573
05C1
04EE
047F
04C5
0512
04F6
04B9
04C9
050D
0525
04FD
04DE
04F6
051C
051B
04FD
04EF
04E9
04C0
047F
0478
04D6
0535
050A
0465
0415
04A5
0555
048A
0187
FD85
FAB5
FA28
FAE5
FB45
FACB
FA5D
FAC7
FBA0
FBEE
FB6F
FACE
FAA2
FAC2
FAC0
FAB0
FAE9
FB53
FB65
FAFB
FAB7
FB1F
FBCA
FBD4
FB21
FA8E
FAC0
FB31
FAFF
FA78
FB28
FE10
022C
0547
0623
057D
04EA
0519
0588
0588
0519
04AD
0483
0487
04AB
04FE
0563
0582
0531
04C1
04A9
04ED
051B
04E2
0483
046E
04A4
04B9
048D
04A3
0558
05F7
0502
01D0
FD99
FA94
F9E2
FAA1
FB24
FAC9
FA53
FA93
FB4A
FB9D
FB42
FACA
FAC0
FAF9
FAF8
FAB4
FA98
FAD5
FB22
FB3A
FB45
FB7A
FB9C
FB49
FAB0
FA8E
FB32
FBE0
FBAB
FAE7
FB2F
FDB5
01B4
0500
0621
0597
04ED
04FD
0556
053D
04B5
045F
0498
0518
056D
057C
0569
0543
0503
04C9
04D2
0513
0529
04DB
047D
0493
0508
0534
04C2
044D
0498
0545
04CD
0228
FE38
FB27
FA45
FADD
FB50
FAF6
FA86
FAC6
FB6E
FBA0
FB20
FA93
FA91
FAF1
FB23
FAFF
FAD6
FAE1
FAF5
FAE4
FAD8
FB08
FB4C
FB43
FAF8
FAEA
FB58
FBBD
FB70
FAC8
FB2B
FDAA
019A
04EF
061A
056A
0477
0464
04F5
0546
0506
04B2
04C0
0507
0516
04E1
04CC
050F
0563
0569
0520
04CF
04A4
0495
049D
04CD
0506
04EF
047C
043C
04BE
0583
0510
026E
FE80
FB5F
FA5C
FAD9
FB4F
FB14
FAC0
FAFB
FB82
FBA0
FB35
FAD9
FAFA
FB4F
FB55
FB07
FACA
FAD0
FAE3
FAD9
FAE7
FB3F
FBA3
FBA4
FB4E
FB32
FB9E
FC05
FBA1
FAA8
FA86
FC88
0050
03EE
05A0
0565
04B2
04C0
0565
05A8
0519
0451
041D
0491
0514
0531
04FF
04D1
04C1
04BC
04C3
04E0
04F3
04D1
0490
0481
04AE
04AC
0439
03D7
0448
0554
057A
0366
FF99
FC2C
FAC0
FB00
FB60
FB03
FA77
FA98
FB4F
FBCB
FBA2
FB40
FB24
FB36
FB16
FAD1
FADC
FB63
FBE9
FBE1
FB5B
FAEB
FAEF
FB37
FB71
FB99
FBCC
FBD5
FB59
FA92
FA9A
FC87
0023
03C4
05B1
05A2
04C6
0464
04A9
04F0
04D1
0498
04AE
04F2
04E9
0479
0416
0428
0490
04E8
0504
04FD
04E3
04A6
0462
0469
04C7
04FF
049A
03F7
03FF
04E1
0557
03C5
001C
FC3B
FA37
FA69
FB6A
FBC4
FB52
FAE8
FB0C
FB71
FB96
FB6C
FB45
FB53
FB7E
FBA1
FBAE
FB95
FB42
FAD4
FAAE
FB0C
FB9C
FBBF
FB4C
FAD8
FAFF
FB8B
FBAD
FB32
FB20
FCC7
0028
03A2
056F
0554
0498
046F
04D4
04FE
04A2
0444
0462
04C1
04CB
0473
043E
0482
04EF
0508
04CF
04B1
04DC
050A
04FE
04DF
04DF
04CA
0453
03C3
03E0
04D3
0570
041E
00A2
FCA8
FA4E
FA2B
FB0F
FB86
FB44
FAF4
FB16
FB69
FB7D
FB56
FB45
FB5C
FB59
FB26
FB02
FB1C
FB3B
FB15
FAD1
FAE4
FB65
FBCA
FBA0
FB3D
FB53
FBDC
FBF7
FB31
FA92
FBD4
FF5F
0376
05C7
05AF
0497
042D
04AC
0520
04EC
0480
048A
04FD
053C
04FD
049E
048C
04B6
04CD
04C1
04C7
04E7
04E4
04A8
047B
049C
04CF
04A9
0447
0453
0509
0572
0415
00A5
FCB4
FA5D
FA4D
FB4A
FBB9
FB3C
FAAE
FAC8
FB46
FB75
FB33
FAFB
FB1B
FB51
FB4C
FB25
FB26
FB43
FB30
FAF5
FB00
FB76
FBD2
FB8B
FAF4
FAE8
FB88
FBDF
FB36
FA75
FB80
FEFB
0334
05B1
05A4
0479
03FC
0483
051E
051C
04C9
04B8
04EC
0500
04DB
04C9
04F2
0518
04FD
04C6
04BB
04CA
04A6
0455
0448
04BA
0535
0512
0474
0447
050A
05C2
04AE
0136
FCEC
FA39
FA0E
FB31
FBCB
FB5E
FAD5
FAF9
FB6B
FB58
FAC5
FA87
FB08
FBA4
FB8F
FAEF
FAA4
FB13
FBB3
FBDF
FBA3
FB71
FB50
FAF3
FA80
FAA0
FB71
FC00
FB6A
FA69
FAFE
FE38
02B1
05C4
0633
0519
045C
049F
051C
0510
04A9
0482
04BD
04FD
0505
04F3
04E7
04CA
048D
046A
049B
04EF
04FB
04B4
048C
04D5
052B
04E5
0418
03B9
0478
0586
0503
01F1
FD8D
FA5F
F9D4
FB08
FBF5
FBA1
FACE
FAA4
FB3B
FBB4
FB83
FB0D
FAF9
FB4C
FB89
FB6C
FB2E
FB14
FB16
FB15
FB1D
FB3F
FB4F
FB25
FB09
FB6C
FC1D
FC36
FB3D
FA34
FAEA
FE0A
0225
04F5
0589
04DD
0471
04B4
050E
0504
04D2
04DF
0510
0501
04A8
046A
0488
04C8
04CF
04AA
04AA
04DE
04F3
04B8
0482
04B2
0511
04FF
0463
0405
0496
0574
04F1
0223
FE25
FB31
FA6C
FB09
FB88
FB67
FB39
FB6F
FBA3
FB57
FAD0
FAC3
FB49
FBB2
FB7B
FAFD
FADF
FB30
FB69
FB46
FB1E
FB48
FB83
FB5C
FAEE
FACE
FB2D
FB76
FB26
FAC7
FBA3
FE54
01DE
0477
0523
0480
03F1
043B
04F6
0550
050A
0499
047B
04A7
04C7
04C1
04CD
0505
0523
04E5
0481
0467
04A0
04C7
04A9
049F
04F3
054C
0523
04A9
04A8
0534
04FC
02A0
FEA3
FB4E
FA60
FB44
FC09
FBB1
FAF3
FAD6
FB47
FB7C
FB31
FAE5
FAF8
FB25
FB17
FAFF
FB37
FB9D
FBBF
FB7D
FB32
FB2F
FB64
FB93
FB94
FB4D
FAB7
FA42
FAF0
FD7A
013D
046E
05B6
055B
04A3
0460
0470
0476
0474
049B
04D6
04ED
04E3
04E2
04E6
04C6
0495
049F
04DF
04E6
0483
041F
042D
047E
04AA
04C9
0542
05B6
04CF
01C9
FDC7
FB04
FA82
FB2E
FB7E
FB32
FB12
FB6C
FBAF
FB70
FB0E
FB08
FB3B
FB39
FB0D
FB1C
FB66
FB74
FB34
FB30
FBA9
FC09
FBB9
FB1B
FAF6
FB3A
FB1D
FAAB
FB4E
FE29
023E
0525
05A5
04DD
048B
04F7
052B
04B3
042E
043B
04A3
04DB
04DA
04F0
0520
0519
04CD
0493
048D
047E
0455
045E
04A4
04B0
0453
0443
051D
05F5
04D6
0121
FCC7
FA72
FAAA
FB8F
FB6B
FA94
FA63
FB23
FBE7
FBFE
FBAE
FB6E
FB37
FAE8
FAC9
FB1C
FB82
FB60
FADD
FAC5
FB56
FBD5
FBAE
FB54
FB68
FB9C
FB3A
FAB4
FBA5
FECB
02B5
051F
055C
04C3
04B2
0513
0519
04B3
0473
048A
0497
0472
0473
04C5
0507
04E4
04A9
04C9
0511
04F3
0482
0469
04CC
04ED
0468
040D
04AA
055C
0432
00A9
FCB5
FAB3
FAD8
FB61
FB1C
FAAC
FB14
FC00
FC4C
FBB4
FB10
FB05
FB3D
FB32
FB06
FB28
FB85
FBA3
FB64
FB2A
FB26
FB1B
FAFC
FB27
FBA6
FBBF
FB06
FA84
FBF2
FF98
038D
0596
0569
0494
046E
04CB
04DA
0477
0426
042F
0463
0499
04D9
0507
04E5
0489
0461
049D
04D5
04AF
0480
04CE
054C
051B
043A
03DF
04BC
0589
042B
005D
FC50
FA5B
FA93
FB46
FB4D
FB19
FB64
FBE7
FBEA
FB7F
FB54
FB96
FBB3
FB55
FAE8
FAF0
FB41
FB56
FB21
FB0B
FB35
FB4F
FB3E
FB5A
FBAB
FB91
FACA
FA73
FC2B
0002
03EF
05CA
0574
049C
0492
0509
0507
0469
03E9
0408
048B
04F8
051B
04FE
04BB
0482
0487
04C6
04EE
04D1
04B1
04D5
04FD
04B8
0442
046B
053E
0552
032C
FF39
FBB3
FA5D
FAD2
FB60
FB28
FAC7
FB00
FB99
FBD5
FB89
FB27
FAFE
FAF9
FB05
FB33
FB6C
FB66
FB25
FB1A
FB80
FBD3
FB74
FAB8
FA9E
FB53
FBC6
FB3D
FAD3
FC78
006B
0480
064F
05AD
0479
0439
04B2
04E6
04A0
0479
04C1
0516
0513
04D3
04A8
04A3
04A4
04A2
04AC
04B7
04B5
04B7
04CD
04C4
046B
041C
0479
0551
0542
0305
FF1B
FB94
FA13
FA5E
FB0C
FB3C
FB2E
FB52
FB86
FB6C
FB14
FAD9
FADB
FAFA
FB30
FB87
FBC3
FB8C
FAFC
FAA9
FAE4
FB44
FB3D
FB05
FB3B
FBC5
FBC1
FB03
FAF2
FD24
013B
04E3
0633
0585
04AE
04B8
051B
04FC
0478
0448
04AA
0521
0537
04F0
0491
0457
0465
04BA
0514
0514
04BA
047C
04AF
0503
04F1
049E
04AF
0516
049A
0228
FE61
FB3C
FA10
FA67
FAE4
FADD
FAB4
FAD7
FB22
FB43
FB44
FB56
FB66
FB47
FB14
FB13
FB41
FB5B
FB50
FB54
FB71
FB69
FB26
FB08
FB54
FB8F
FB12
FA4F
FAE0
FDCA
0200
0544
0657
05E7
054F
0515
04E8
04A2
0495
04E4
0527
0504
04B2
0499
04B6
04C0
04B4
04CE
0507
050A
04BD
047A
0482
0498
047B
0482
0524
05D5
0517
021D
FE04
FAE1
F9C0
F9F9
FA64
FA9B
FAD7
FB26
FB47
FB33
FB2F
FB53
FB5F
FB41
FB4A
FB92
FB9F
FB14
FA69
FA78
FB40
FBD8
FBA9
FB41
FB61
FBBA
FB67
FAA8
FB2B
FE0E
0228
0514
05C0
053E
0514
0573
0588
0501
0479
047C
04C6
04D2
049F
0485
0494
0496
0488
04A2
04EA
051D
0517
04F7
04CA
0469
03F4
0413
0515
05EF
04D4
0145
FD08
FA86
FA62
FB26
FB39
FA8C
FA20
FA76
FB16
FB63
FB5D
FB55
FB63
FB71
FB88
FBB0
FBBF
FB8C
FB46
FB32
FB42
FB32
FB11
FB3C
FBA8
FBA6
FADB
FA4B
FB99
FF15
0301
054F
05A1
0536
051E
0544
052B
04EF
04FC
0541
053C
04D5
0488
049E
04B8
047E
043B
045E
04B0
04A4
0442
042D
049A
04E4
049A
0459
04EA
059A
0484
00E9
FC95
FA25
FA43
FB46
FB76
FADD
FA91
FAEF
FB44
FB0A
FAA8
FABC
FB2F
FB72
FB53
FB23
FB2A
FB67
FBB5
FBEC
FBDB
FB7C
FB2F
FB62
FBDE
FBCA
FAE0
FA53
FBD2
FF7F
036F
0591
05AA
050D
04C8
04D2
04D0
04DC
0523
054F
04F8
046C
0466
04F5
054A
04E6
0458
045A
04B8
04BD
0464
0457
04BB
04D3
043D
03D7
0485
0561
0449
0092
FC4F
FA1E
FA55
FB21
FB1B
FAB6
FAEF
FB9D
FBC6
FB30
FAB0
FAD8
FB3C
FB49
FB25
FB3C
FB69
FB44
FAF9
FB1D
FBAD
FBF1
FB8F
FB1F
FB3A
FB7D
FB3C
FB02
FC5F
FFD1
03A5
05A7
0581
04B8
0495
04F1
0516
04FB
0508
052D
04F2
0462
0428
0489
04F0
04D7
0495
04B4
04FC
04D3
0453
0437
04AB
04F8
04B0
0482
0513
0564
0399
FF8F
FBA9
FA48
FB21
FBF4
FB77
FA87
FA6A
FB02
FB56
FB2F
FB35
FB9E
FBC4
FB49
FACF
FAFC
FB71
FB6E
FB0B
FB04
FB74
FBAD
FB5E
FB26
FB72
FB9C
FAFC
FA91
FC47
0054
0450
05C2
04ED
041B
0496
056D
0554
0490
044E
04CA
051B
04C3
0464
049A
04FD
04E7
048E
049F
050A
0520
04B4
0468
049D
04D4
049C
046E
04DD
051D
0384
FFCB
FBF0
FA25
FA77
FB31
FB38
FAF9
FB25
FB79
FB5A
FAFE
FB19
FBA8
FBDB
FB5C
FADA
FAFC
FB69
FB73
FB27
FB0B
FB24
FB06
FAC2
FAEE
FB80
FB80
FA92
FA42
FC90
0124
051B
0628
0515
045F
04FA
05A9
0542
045D
0437
04D1
051C
04AE
044C
048F
0502
04FD
04B4
04BE
0509
050E
04CE
04C9
0511
0520
04D9
04EE
0594
0575
02EE
FE75
FAB7
F9C5
FADE
FBB6
FB51
FAA2
FAAF
FB2B
FB4B
FB0B
FAFF
FB35
FB26
FABF
FAA0
FB17
FB93
FB81
FB31
FB39
FB74
FB53
FAF2
FAF6
FB5C
FB46
FA84
FA98
FD2C
019A
0523
05E4
04D7
043D
04D1
0575
053C
04A2
048B
04EB
051A
04FA
0500
0547
0554
04F2
04A3
04C8
0501
04D7
048A
049B
04D6
04A8
0449
0499
0583
0553
0290
FE32
FAFF
FA78
FB54
FB85
FACA
FA77
FB26
FBDE
FBA4
FAE0
FA9B
FAF6
FB2E
FAEA
FAB5
FAFB
FB4B
FB1F
FAB8
FAB6
FB1A
FB67
FB79
FB97
FBB1
FB4E
FAA4
FB12
FDB8
01BC
04C6
0576
04C0
046D
04F6
056F
0535
04BF
04B6
04F7
04F7
04AB
0485
04AF
04DA
04D6
04E2
0524
054C
0517
04D1
04DD
050C
04EF
04B3
04ED
055F
049F
01A6
FD7A
FA88
FA24
FB3D
FBDE
FB72
FAE8
FAFF
FB51
FB36
FAE0
FAFB
FB92
FBE3
FB75
FACB
FAAB
FB14
FB4D
FAFB
FA9E
FAD7
FB76
FBA5
FAFA
FA44
FB05
FDF7
0212
0542
0629
0545
0444
0441
04E3
052A
04D6
048D
04C8
0526
0519
04BE
04A4
04DE
04E6
0481
0440
04B1
0565
0570
04C5
047B
053E
05F6
04BC
0122
FD00
FAA8
FAA7
FB92
FBDD
FB58
FADE
FAFD
FB63
FB87
FB51
FB0C
FAE4
FAC8
FAAE
FABB
FB0D
FB73
FB91
FB4D
FAFB
FAF8
FB21
FAF0
FA4B
FA16
FB99
FF17
0319
058B
05A1
047D
03D9
0444
04EE
04FF
04A5
0494
04EE
0528
04EA
04A1
04D1
054B
0568
04FC
04A1
04CF
0528
0500
0473
046A
0549
05F3
04B5
012F
FD09
FA7B
FA42
FB35
FBC8
FB88
FB1A
FB0D
FB35
FB23
FAE7
FAED
FB4E
FB8E
FB47
FABC
FA8D
FAE3
FB3C
FB26
FAE1
FB00
FB7E
FBA3
FB07
FA81
FB8F
FEB1
0295
0530
05A0
04D3
044A
0491
0511
0525
04EB
04E1
0511
0512
04BD
047C
04B4
051F
0525
04BB
0488
04F3
0571
052F
0451
03F8
04BF
058F
0485
011E
FD10
FAA9
FA92
FB73
FBB3
FB20
FAA3
FAD2
FB41
FB48
FAEB
FAB1
FAD8
FB0C
FAFD
FAD9
FB01
FB68
FB98
FB5B
FB18
FB43
FBA2
FB7E
FAB2
FA4B
FBB8
FF32
0326
0584
059B
0498
041B
049D
0553
0574
0525
0501
0523
051B
04C6
04A5
0520
05C1
05A7
04B7
03DD
03E5
0482
04CE
049A
04AC
0565
05BE
042D
008C
FCA0
FA76
FA77
FB50
FB99
FB29
FABA
FABC
FAE7
FAE1
FACB
FAF8
FB57
FB76
FB20
FAB9
FAC9
FB4C
FBB2
FB95
FB3B
FB32
FB7C
FB7A
FADB
FA74
FBBB
FF23
033E
05D3
05FC
04E1
0451
04D8
0586
0570
04D4
049A
04FB
0551
0511
0491
046E
04A8
04BC
0489
048E
0510
0577
0511
0432
0406
04EF
0594
0427
007C
FC7D
FA4B
FA3E
FAFA
FB32
FAD8
FA9C
FAC8
FB01
FB03
FB00
FB34
FB70
FB58
FB04
FAED
FB47
FB9F
FB6E
FADF
FAAE
FB30
FBC3
FB8C
FAB0
FA8C
FC6A
000C
03AF
0599
0594
04D3
0494
0504
057C
057C
0527
04DA
04AD
0488
047E
04C6
0546
057C
0515
0474
044E
04C7
0533
04F8
046D
0477
0531
055C
038B
FFD5
FC07
FA09
FA26
FB10
FB70
FB19
FABC
FACB
FB09
FB17
FB05
FB1B
FB49
FB32
FACA
FA8E
FAE6
FB81
FB9C
FB07
FA76
FAA7
FB53
FB81
FAE9
FAB2
FC60
0005
03E9
061D
063B
056E
04EE
04E4
04CE
0489
0480
04E9
0556
0540
04C3
047A
04A8
04E8
04D2
0499
04BC
0532
055C
04EA
0479
04DE
05D2
05CB
037E
FF69
FB9D
F9D5
FA01
FAB9
FAE5
FAA8
FAB8
FB39
FB9A
FB6B
FAF8
FAE0
FB41
FB9D
FB8E
FB42
FB23
FB3C
FB3C
FB09
FAF9
FB40
FB6B
FAE2
F9FE
FA2C
FC98
00B4
0473
0622
05E9
0543
0540
059F
059A
0517
04B0
04C6
04FE
04D9
046C
0440
048E
04F1
04F7
04B8
049D
04C9
04F1
04E2
04E0
053D
05A8
0525
02F1
FF6D
FC08
FA22
F9EF
FA81
FAD1
FAA4
FA7B
FAB3
FB0D
FB19
FAE2
FAE3
FB4D
FBB5
FBA1
FB38
FB08
FB3E
FB64
FB20
FAC5
FADA
FB36
FB26
FAA1
FADB
FD13
00F4
048D
0627
05D7
0510
04EB
0544
056E
0541
051A
0529
0532
0501
04C8
04C7
04DE
04BD
0466
0447
04A5
0525
0530
04B7
0464
04C8
0575
0519
02C3
FEF9
FB7F
F9DB
FA15
FAEB
FB37
FAEE
FABE
FAFC
FB42
FB1E
FABD
FAA5
FAF3
FB36
FB26
FB0E
FB53
FBBD
FBB3
FB27
FACF
FB2D
FBB3
FB70
FA8F
FAA4
FCFD
00F5
0461
05BA
0577
0517
054E
058E
053B
04A8
0490
0501
0555
0528
04D9
04E6
0524
0502
0471
0410
0453
04D2
04D5
045B
0434
04E5
05BB
0542
02BF
FF0E
FBF4
FA99
FAB0
FB0F
FAED
FA7D
FA66
FAD1
FB3B
FB2C
FAD7
FACA
FB21
FB60
FB2F
FAEA
FB1D
FBAD
FBE7
FB7E
FB09
FB2A
FB8B
FB48
FA75
FA91
FCF9
0111
048E
05BD
051B
0476
04CB
0583
05A4
052B
04DC
0513
0557
0529
04BB
0499
04CF
04E3
0499
0460
04AF
053C
053F
0493
041F
04B7
05BC
0565
02A8
FE99
FB7B
FA8B
FAFD
FB42
FADE
FA8F
FAE7
FB6E
FB62
FADA
FAA0
FB04
FB6D
FB47
FAE5
FB02
FB98
FBC4
FB09
FA29
FA42
FB4B
FBF9
FB64
FA60
FAC9
FD7F
0165
046D
0585
0541
04DC
04E6
050D
04E9
04A3
04A8
0507
0548
050B
048E
0468
04C3
0529
0524
04DD
04DD
0540
057E
052F
04BB
04D8
0550
04CD
0240
FE57
FB28
FA2F
FAEF
FBB5
FB8B
FAF1
FACD
FB2B
FB57
FB0A
FACB
FB1C
FBB1
FBD2
FB5C
FAE7
FAE6
FB09
FAD2
FA75
FA9A
FB4C
FBA5
FAF8
FA17
FAD5
FE06
0251
054D
05D3
04E0
043A
048C
051F
0520
04B3
048C
04E0
0527
04EB
0479
046A
04CE
0519
04F4
04BA
04EB
0559
055B
04CE
0477
04FD
05B8
0501
0205
FDEE
FAEA
FA20
FACB
FB65
FB48
FAF7
FB08
FB59
FB66
FB1F
FAF3
FB21
FB58
FB2F
FACC
FABB
FB28
FB96
FB79
FAFC
FAD2
FB3A
FB87
FB10
FA61
FB0D
FDF0
01F2
04E0
0598
0501
04B7
0528
0577
0504
0465
0481
0537
058E
0515
047F
049B
0528
053A
049D
042A
048E
0543
053E
047A
041F
04F0
05F6
0548
0225
FDF3
FAFB
FA41
FADC
FB4D
FB10
FABE
FAE2
FB34
FB1A
FA99
FA5F
FADA
FB94
FBCD
FB6F
FB1A
FB32
FB5A
FB1F
FAC9
FAFD
FBA9
FBD9
FAFF
FA19
FAF4
FE2D
0240
04F2
056E
04C6
047C
04FA
0591
0597
052E
04E5
04F5
0514
04EE
049B
046D
047F
049A
049B
04AD
0501
055F
0545
04AB
0450
04D3
058F
04D4
01C0
FD8F
FAA3
FA2D
FB1E
FB9D
FB19
FA84
FAB8
FB52
FB6D
FAF3
FAA5
FAF5
FB77
FB90
FB51
FB3B
FB6E
FB7B
FB20
FAC9
FAF7
FB72
FB6E
FAB3
FA3D
FB77
FEBC
02B8
0577
060C
053D
0484
049B
050B
051B
04C3
0493
04CD
0508
04D4
046A
045B
04B9
04FB
04D1
04A8
04FF
0583
0569
04A9
044B
04FD
05BD
049A
00FF
FCB7
FA32
FA1E
FB0A
FB60
FB0B
FAF2
FB5E
FBA2
FB3E
FAB2
FAC6
FB65
FBB6
FB52
FAD4
FAEF
FB72
FB89
FAF5
FA70
FAB1
FB5C
FB74
FAC5
FA76
FBEF
FF40
02E8
0532
05A5
051D
04AC
04A7
04C1
04C3
04D3
0511
0546
0522
04BF
0495
04DA
0528
04FC
047F
045F
04E4
0571
0548
0499
0458
04EB
0554
0414
00E9
FD40
FAE6
FA60
FACA
FB13
FAFB
FAED
FB2F
FB84
FB89
FB3B
FAF2
FAF6
FB2A
FB43
FB2E
FB22
FB43
FB64
FB42
FAF4
FAE3
FB29
FB42
FAD3
FA98
FC00
FF76
0377
05D1
05D8
04E2
048A
04F1
051F
04A5
042B
0456
04D6
0501
04D1
04BF
04E0
04D1
048B
0491
0514
0563
04E0
0426
0462
0565
0541
027C
FE20
FADF
FA2B
FAF2
FB4F
FAD1
FA77
FAE5
FB8A
FB9E
FB40
FB17
FB43
FB52
FB1C
FB06
FB48
FB7D
FB43
FAF3
FB24
FBA4
FB96
FAD2
FAA7
FC96
0066
0408
059F
054B
04A4
04C2
054B
056B
0506
04B1
04B5
04C5
04A4
049B
04F2
055A
0547
04C2
0473
04AE
04FE
04E7
04B6
04FD
054D
043E
0113
FD0A
FA5E
FA0B
FAF9
FB85
FB41
FAE9
FB08
FB55
FB5D
FB36
FB2F
FB38
FB0C
FAC6
FACA
FB17
FB31
FAF1
FAE8
FB83
FC1F
FBB8
FA92
FA8D
FD2A
018B
050D
05FA
0519
0463
04A9
0521
04F6
047A
047E
0504
054B
04FD
04A1
04C1
0521
0534
04FC
04EC
050F
04EB
0472
0456
04F5
0538
0379
FFAD
FBEF
FA65
FAF9
FBC6
FB89
FAD7
FAD1
FB63
FB8F
FB07
FA9D
FAF1
FB85
FB90
FB2F
FB0B
FB3B
FB2C
FABF
FAA1
FB2F
FBA3
FB2A
FA88
FBA7
FF2E
034B
057D
0544
044E
0435
04E1
054B
051E
04E2
04F2
0504
04D9
04B8
04E1
0503
04BB
045A
0483
051F
0553
04C7
0459
04F3
05EB
054F
0220
FDCD
FADE
FA6F
FB55
FBD0
FB68
FAE4
FAE4
FB26
FB27
FAF5
FAF6
FB35
FB50
FB15
FAD6
FAE6
FB20
FB31
FB28
FB52
FB92
FB5A
FAA1
FA84
FC60
0025
03F8
05E1
05A2
04AE
0463
04C5
0507
04D3
0494
04A8
04DF
04E1
04C6
04DF
0525
0540
0516
04F2
0503
0506
04C2
0494
04E8
053D
0431
0115
FD25
FA9A
FA69
FB5E
FBB1
FB09
FA84
FAF5
FBC8
FBF4
FB66
FAF8
FB2B
FB86
FB73
FB12
FADD
FAE3
FAD7
FAC1
FAFB
FB6A
FB65
FADC
FB1D
FD8D
01A4
04FB
05CC
04D7
0434
04C1
0576
053D
0479
0441
04B7
0501
04B7
046F
04AF
050E
04F6
04A7
04C6
052E
051B
0485
046D
053E
059C
03AA
FF8D
FBB2
FA3E
FADD
FB99
FB60
FAD1
FACD
FB2B
FB43
FB10
FB19
FB6F
FB80
FB09
FA9A
FACC
FB57
FB85
FB4A
FB47
FBAA
FBB0
FAD4
FA10
FB33
FEC6
0312
05A6
05BF
04BD
0457
04CF
0539
0501
0499
049F
04F3
050C
04D0
04B1
04E8
0520
0504
04CB
04CE
04DF
049E
0453
04B7
0597
055C
02AC
FE58
FAED
FA11
FAED
FB85
FB25
FABB
FB0B
FB8A
FB64
FAD2
FAAF
FB1E
FB69
FB32
FAFE
FB3B
FB78
FB1F
FA98
FACA
FB93
FBB4
FAB4
FA28
FC17
005A
046C
0610
0582
04AD
04C1
0541
0549
04E2
04AF
04D8
04F1
04CB
04B6
04E7
050E
04DC
0496
04BA
052E
054F
04E2
0493
0505
0589
0475
010C
FCC1
FA07
F9E3
FB0C
FB94
FAFF
FA5F
FAA5
FB6F
FBC4
FB6F
FB11
FB16
FB32
FB10
FAE2
FAF5
FB18
FAF6
FAC2
FAF2
FB5C
FB3B
FA95
FAEF
FDBA
022F
059B
063D
051F
0487
0529
05C1
0540
0453
0434
04D2
050C
0485
0429
04AA
0566
0569
04E4
04CB
053C
0551
04B3
0457
04F6
055F
0387
FF49
FB28
F9A9
FA94
FB94
FB3C
FA62
FA6B
FB3F
FBAF
FB52
FB00
FB5D
FBDD
FBB0
FB08
FAC9
FB24
FB5D
FB0D
FACD
FB32
FBB5
FB76
FAF5
FBF8
FF58
037F
05E3
05C4
04BE
0498
054B
05A2
0527
0498
0497
04CE
04AF
046C
048D
04EE
04E7
046A
043A
04B9
052D
04CB
0410
0428
04FA
04B5
01EC
FDAD
FA9D
FA18
FAFB
FB61
FADE
FA74
FACA
FB57
FB68
FB27
FB28
FB64
FB5C
FB0B
FB03
FB7C
FBE0
FBA8
FB3D
FB67
FBFD
FBFC
FB24
FADE
FCD6
00CC
0481
0602
0588
04CA
04DB
054C
0551
04F0
04BE
04DF
04E9
04AD
0486
04B4
04DF
04A2
043D
0441
04A3
04B6
0444
0411
04B7
0554
0422
009B
FC7D
FA2D
FA42
FB39
FB76
FAEF
FA9E
FAEA
FB44
FB30
FAF5
FB07
FB41
FB3B
FB0E
FB34
FBAF
FBDC
FB6D
FB02
FB4F
FBEF
FBD7
FB0C
FB33
FDC8
01FF
0543
05E4
04C6
0410
04A9
0593
05A2
04F9
048F
04C4
0515
050D
04D9
04C6
04BB
0493
048C
04EB
054E
0511
045A
0427
04D5
0519
0336
FF45
FB88
FA1D
FACE
FBB2
FB8C
FADB
FAA3
FAF1
FB1F
FAF9
FAF6
FB48
FB7A
FB39
FAE9
FB06
FB52
FB37
FAD2
FADE
FB7F
FBD2
FB3A
FAB1
FC07
FF9F
039E
05C0
05A0
04BB
0479
04D4
050B
04E9
04DD
0518
0536
04ED
048F
0496
04EE
051A
04F5
04D7
04F2
04F8
04A9
0468
04BD
0539
047D
01B1
FDCB
FAE6
FA30
FAE6
FB73
FB3B
FAE1
FB03
FB5C
FB53
FAED
FAB8
FAF4
FB46
FB51
FB33
FB2A
FB1E
FAEB
FADD
FB55
FBF2
FBD1
FAF7
FAE8
FD23
0122
0493
05BD
052F
04AA
04EB
0534
04DF
0469
0498
0533
0560
04F8
04B0
04F4
0544
0511
04AA
04BB
051B
04F6
042F
03D2
0491
0551
0418
0079
FC61
FA2A
FA45
FB38
FB92
FB40
FAFA
FB0A
FB1B
FAFF
FAF2
FB16
FB26
FAEA
FAAB
FAD4
FB47
FB7B
FB46
FB29
FB84
FBE0
FB85
FACB
FB3E
FDF9
0214
0541
060F
0539
0483
04BE
0548
054D
04E0
04A2
04C6
04F5
04FA
0502
051B
04FC
0497
0461
04B3
0518
04E3
044A
0450
052C
0569
0357
FF51
FBB3
FA5A
FAC4
FB22
FAB4
FA51
FAC2
FB86
FBA8
FB2B
FAE1
FB1F
FB5E
FB39
FB15
FB56
FB93
FB33
FA90
FAA7
FB87
FBFC
FB3F
FA78
FBB5
FF56
0357
056D
0568
04E1
0502
0571
055F
04DD
049F
04D5
04FF
04CB
048D
049F
04CA
04AD
047B
04B6
0541
0559
04B4
042B
04A8
059F
0534
0247
FDFE
FACD
FA09
FAD6
FB78
FB39
FABA
FAB4
FB11
FB49
FB38
FB2D
FB53
FB75
FB69
FB56
FB68
FB74
FB48
FB13
FB34
FB84
FB5F
FAB1
FAA1
FC9E
0095
0481
0644
05AB
046C
041E
04C1
0548
0522
04B5
0492
04BE
04E7
04EC
04E2
04C2
047F
044D
0471
04C1
04BD
045D
0453
0502
057B
0420
0096
FC96
FA57
FA62
FB4D
FB94
FB1E
FAC5
FAF5
FB54
FB79
FB6B
FB4F
FB1B
FADC
FAEB
FB73
FBF7
FBD3
FB32
FB00
FB97
FC12
FB80
FA82
FB01
FDF7
0211
04EF
0595
0510
04DC
0536
0560
0503
04A4
04BE
0505
04F3
049C
0480
04B1
04B6
0459
0418
0472
0503
04F5
044B
0412
04D2
0550
03A7
FFAB
FB8C
F9A6
FA22
FB34
FB66
FAFD
FAEB
FB45
FB5E
FB09
FADE
FB34
FB8F
FB76
FB38
FB5B
FBA9
FB87
FB12
FB13
FBAE
FBE5
FB0D
FA55
FBC5
FFA1
03B0
059A
054C
0486
0485
04FE
0533
0515
0504
0508
04E8
04AE
049F
04B0
0497
0474
04B3
0533
0530
047D
040A
048E
0507
03A0
0013
FC5E
FAA4
FAEC
FB8F
FB70
FAFA
FAE9
FB1C
FB22
FB0E
FB33
FB61
FB3E
FAFB
FB12
FB67
FB66
FAFE
FAE0
FB5A
FBAF
FB3F
FB04
FCC6
009F
0457
05C9
0531
0468
047B
04EA
0509
04F6
0509
051A
04DE
0490
049C
04D5
04BB
0469
0486
0514
0545
04D9
04B7
0554
055A
0309
FEC7
FB23
FA0E
FAD1
FB63
FAFF
FA95
FADE
FB53
FB46
FAFD
FB07
FB3B
FB2E
FB13
FB50
FBA2
FB77
FB07
FB15
FB95
FB82
FA9D
FA8E
FD29
01B7
0544
05F2
04EF
047C
0517
0595
054F
04DF
04D7
04EC
04B9
048A
04C5
0520
050A
04B1
04B8
050E
04F9
047B
048B
053D
04E0
0201
FDBA
FAC4
FA5E
FB2F
FB63
FAD7
FA93
FAE9
FB1D
FADB
FABC
FB24
FB82
FB55
FB0D
FB30
FB63
FB1D
FAC4
FB10
FB9F
FB64
FA9A
FB31
FE78
02F6
05B8
05AC
0497
0476
052B
0574
0512
04D8
051B
0552
0520
04DA
04D4
04DD
04C4
04C8
0511
0531
04CC
047A
0502
05A5
046B
00B7
FC92
FA7B
FAA4
FB45
FB31
FAD8
FAF1
FB36
FB18
FACE
FAF3
FB5A
FB4B
FAC7
FAA5
FB1F
FB64
FB06
FAC9
FB3C
FB85
FABE
FA06
FB9B
FFCE
040E
05BD
051A
0475
04FB
05A3
055F
04CB
04E6
055C
0537
048E
0454
04C6
0524
0503
04DD
0505
0503
0487
0453
051C
05C6
0428
FFFD
FBD8
FA54
FB25
FBF2
FB77
FA8B
FA54
FAB7
FAED
FAD3
FAD9
FB1C
FB45
FB35
FB34
FB4B
FB2B
FAEC
FB15
FB91
FB74
FA8F
FA72
FCCA
00FE
047E
0580
04C4
0435
0498
0535
0561
0555
0560
0546
04DE
04A2
04E6
0536
0508
04AD
04BB
04FE
04D1
0464
04A3
058D
0572
02CB
FE76
FB1D
FA49
FAF6
FB5B
FB13
FADB
FAFA
FB0A
FAEA
FAF0
FB28
FB2D
FAE9
FAD8
FB36
FB77
FB21
FAC2
FB1E
FBBB
FB5C
FA41
FA9D
FDDC
026D
055B
05AD
0503
0508
0581
0565
04C1
048B
04FB
0537
04D3
0480
04CF
053A
0518
04B9
04BA
04E0
049C
0456
04EA
05D9
051A
018A
FCDB
FA0D
FA1A
FB33
FB5F
FABC
FA81
FAEE
FB44
FB2C
FB0F
FB27
FB2C
FB0E
FB22
FB73
FB75
FAF5
FAB2
FB48
FBEE
FB6E
FA67
FB44
FF1D
03D1
063B
05C5
0495
0480
052B
0554
04DB
0499
04D7
04FE
04C9
04B4
04F8
050F
04A9
0463
04BA
051B
04DA
0472
04C3
053B
03F9
004D
FC17
F9F3
FA53
FB5A
FB72
FAEC
FACA
FB10
FB27
FB0B
FB29
FB65
FB4A
FAF2
FAF8
FB6E
FBAC
FB61
FB20
FB66
FB9E
FB16
FAB0
FC53
0047
043F
05D9
0546
048C
04C6
0543
0531
04DA
04E5
052E
051D
04BC
04A4
04EC
04FD
049D
0459
047D
0491
045C
0486
0555
0579
0348
FF22
FB7E
FA49
FAEB
FB70
FB0C
FA90
FAB1
FAFC
FAE3
FAB7
FAF2
FB4A
FB3D
FB08
FB2E
FB83
FB7C
FB3B
FB60
FBCD
FB90
FA8F
FA7E
FD14
0184
04EB
0598
04C2
0481
0523
058D
054E
0513
053E
054F
04E8
0483
04A9
0505
04F3
049E
04A9
04F7
04CD
044B
0484
057C
0544
024A
FDC9
FAB7
FA64
FB56
FB93
FAF4
FA95
FAD6
FB04
FACA
FABC
FB2D
FB83
FB49
FB01
FB37
FB7B
FB37
FADD
FB2E
FBC2
FB78
FA8A
FAF9
FE26
02A2
0584
05B2
04CC
04A4
051A
0526
04C5
04C0
052E
0560
051C
04E7
0503
0506
04B4
0485
04D6
0521
04C6
0457
04D5
05AD
04BD
0118
FCB7
FA59
FA69
FB19
FB13
FAC9
FB0A
FB8C
FB85
FB09
FAD6
FB09
FB02
FA9F
FA8E
FB12
FB73
FB32
FAF9
FB5F
FBB2
FB0E
FA56
FBA2
FF7B
03B4
05BB
056C
04BF
04F9
0570
0532
049F
0490
04EC
04FF
04C6
04D2
052E
054F
0514
04F5
051D
0505
0479
0446
0505
0591
03E9
FFDF
FBDB
FA39
FAB8
FB56
FB09
FA7F
FA86
FAE7
FB0D
FB03
FB24
FB60
FB5A
FB20
FB19
FB3D
FB23
FADF
FB0D
FB9E
FB96
FAAF
FA76
FCA9
00D0
0468
05A5
052B
04C2
0510
0562
0539
0506
052C
0549
0500
04AE
04C1
04F0
04CA
0494
04C9
051B
04DB
0444
046F
0572
0587
02ED
FE71
FAF2
FA2E
FB0B
FB7A
FB07
FAAE
FAE8
FB26
FAFD
FACE
FAFD
FB3D
FB29
FAFD
FB2A
FB7E
FB70
FB24
FB40
FBA7
FB6D
FA8E
FAC4
FD96
0204
0547
05D8
04DC
0452
04C0
0537
051B
04DD
04F9
052E
0517
04EA
04FB
0516
04EA
04A9
04A8
04B2
0470
043C
04BA
0578
04C7
01A0
FD58
FA86
FA44
FB3A
FB9C
FB2D
FAD6
FAFB
FB2C
FB21
FB12
FB23
FB1E
FAEB
FAD2
FAFF
FB28
FB14
FB1C
FB90
FBE1
FB4F
FA82
FB6D
FEEF
0347
05C9
05C1
04CB
048C
04FC
0536
0503
04E8
0515
051B
04CC
049D
04D2
0509
04ED
04C1
04C8
04AD
043B
0416
04DA
059C
046B
00B0
FC62
FA24
FA6B
FB61
FB64
FAC0
FA8B
FAE7
FB20
FAF9
FAE1
FB11
FB42
FB48
FB4B
FB5F
FB53
FB2B
FB4D
FBC6
FBDC
FB17
FA8C
FC1E
000A
0419
05E9
057A
04AA
04BE
0546
0563
050E
04D9
04F1
0506
04F2
04DC
04CA
0493
0465
049C
0500
04DF
0440
0430
0511
0569
0359
FF2B
FB62
FA0B
FAAC
FB59
FB2B
FAD3
FB00
FB53
FB42
FB07
FB14
FB3F
FB2E
FB13
FB49
FB8C
FB63
FB0C
FB36
FBBC
FB99
FA9F
FA7C
FD03
018A
0532
0615
0534
04B0
0516
0564
0506
0492
0497
04CF
04C9
04A8
04C2
04EE
04CD
048D
04A7
04ED
04C4
045B
04A5
0594
055B
027E
FE16
FAE1
FA3B
FAF4
FB3C
FACF
FA9B
FB02
FB62
FB45
FB10
FB26
FB49
FB35
FB34
FB79
FB96
FB39
FAEB
FB40
FBA9
FB30
FA50
FB00
FE51
02A8
0547
0567
04BA
04DE
057A
0570
04CF
0483
04C2
04EA
04B8
04A0
04E0
0502
04B8
0471
04A1
04E3
04A4
045A
04EB
05C3
04CA
0115
FCA4
FA51
FA9D
FB86
FB66
FAB4
FAB1
FB61
FBB8
FB54
FAF1
FB20
FB73
FB60
FB21
FB2C
FB5D
FB5A
FB4C
FB76
FB7E
FAF4
FA8F
FBE4
FF6F
0381
05C0
05A1
04B3
0481
04F4
051A
04B6
0460
0478
04BE
04E3
04E0
04CB
04AE
049C
04A5
04A4
0467
042D
048E
057B
05AB
03B2
FFD7
FC28
FA72
FA8A
FB0D
FB2E
FB2C
FB54
FB70
FB49
FB20
FB46
FB86
FB7B
FB39
FB31
FB6C
FB85
FB6C
FB95
FBFF
FBE3
FAED
FA68
FC26
0025
041E
05CE
054A
047C
04A8
053F
0534
0493
0438
0471
04BA
04B0
0495
04B4
04DC
04BC
047B
0478
04A3
0498
045D
0488
053F
0575
03D3
0060
FCD4
FAF8
FAF5
FB86
FB8F
FB26
FAF9
FB3C
FB82
FB7D
FB5E
FB67
FB72
FB3E
FAF8
FB0D
FB7D
FBC2
FB86
FB2B
FB30
FB67
FB35
FAC4
FB59
FDF0
01BD
04A5
0561
04AD
0429
0474
04E5
04D4
047B
0468
049C
04B4
04A5
04BE
04F7
04DD
0456
0404
046A
050A
0507
047E
047C
054D
0584
0369
FF4D
FB99
FA4F
FB04
FBCA
FB96
FB12
FB26
FB99
FBA4
FB36
FB06
FB65
FBCA
FBAF
FB57
FB48
FB6B
FB4A
FAFA
FB11
FB97
FBA9
FACA
FA1E
FB84
FF4A
036D
059A
057A
049F
0468
04BB
04D9
04A4
048F
04AB
048D
041B
03E8
0458
04F5
050B
04AC
0488
04D6
04FF
049E
044D
04C9
058D
04EF
0203
FDF5
FB0B
FA6A
FB36
FBD9
FBA9
FB1D
FAD1
FAE3
FB28
FB87
FBE3
FBEF
FB86
FB02
FAEF
FB4D
FB85
FB3F
FAF4
FB3E
FBD5
FBC7
FAF6
FAC3
FCB7
0089
040C
0561
04C9
0408
043F
04F6
0534
04DB
0488
0487
048E
0469
045B
049D
04E8
04E7
04C6
04E5
0518
04D0
0422
03FD
04D5
0580
042F
00A2
FCC8
FAD7
FB10
FBDA
FBD7
FB36
FAE9
FB34
FB85
FB74
FB45
FB4F
FB71
FB5E
FB24
FB11
FB31
FB3F
FB28
FB3F
FBA5
FBD9
FB56
FAA1
FB2F
FDDD
01B6
04A1
0565
04AF
0415
0456
04E7
0509
04C7
04A5
04C8
04DD
04C2
04BF
04F8
0517
04C8
0452
043D
0483
0498
045C
046C
050D
0533
035C
FF97
FBF4
FA78
FB07
FBDA
FBBC
FB1F
FAFC
FB59
FB82
FB3E
FB09
FB1E
FB1D
FACE
FAB7
FB4F
FC10
FC11
FB60
FB02
FB70
FBC6
FB24
FA65
FB82
FF18
0346
058D
056F
048C
0467
04E7
051C
04C8
0483
04A7
04DE
04CD
04AA
04C7
04F2
04C4
0465
0465
04D7
0510
04A6
043D
04AB
057E
04FB
0211
FDE1
FAD7
FA3B
FB1C
FBB2
FB5A
FACE
FAC9
FB22
FB4B
FB35
FB34
FB5B
FB60
FB29
FB00
FB1C
FB3F
FB29
FB19
FB6B
FBD1
FB8B
FAA7
FA90
FCB9
00BB
045E
05BF
0519
0434
0445
04F2
054A
0519
04DD
04E0
04E5
04C4
04C0
050F
0562
054F
04F6
04D3
04F3
04D6
0455
041A
04AE
053F
0418
00A9
FC98
FA50
FA85
FBB0
FC01
FB45
FA9A
FAB7
FB2E
FB4E
FB16
FAF0
FAEF
FACC
FA90
FA9D
FB06
FB50
FB2B
FB00
FB46
FBA2
FB54
FAA4
FB2C
FE13
024B
054E
05B7
04A0
0410
04A8
055F
0547
04B9
0496
04F3
0532
050C
04E9
0513
0537
0500
04B5
04C6
0501
04D6
0468
048F
056C
0590
035B
FF31
FB86
FA5A
FB28
FBD9
FB5B
FA8B
FA90
FB33
FB6A
FAF4
FAA0
FAF7
FB76
FB6C
FB0B
FAFE
FB49
FB52
FAFB
FAE9
FB67
FBAB
FAFF
FA4F
FB88
FF2F
034A
0560
0519
0443
0461
0522
056A
0511
04DD
051E
0541
04DE
0472
0492
04F4
04EB
048A
0489
050A
0542
04B6
0433
04B8
05AD
051F
020D
FDEA
FB2E
FABB
FB54
FB79
FB08
FAC5
FAF1
FB15
FAEE
FADF
FB38
FB9F
FB91
FB38
FB29
FB6F
FB72
FAF8
FAA6
FB15
FBBE
FB86
FA7E
FA5F
FCBB
00EE
0481
05AF
0507
0465
04AC
0537
0534
04D2
04BC
04FB
0501
04A0
045E
049D
04FD
04F1
04A0
049B
04E2
04DC
0471
0475
055D
05FE
0478
008A
FC54
FA44
FA97
FB85
FB91
FB00
FAD3
FB26
FB46
FAF7
FAC9
FB1A
FB73
FB44
FAD2
FAD1
FB4E
FB99
FB5F
FB25
FB5C
FB83
FAE8
FA24
FAEC
FE16
0241
0510
0589
04CF
0476
04CD
051F
0508
04EB
0512
0528
04D5
0473
0498
0527
0560
04F4
047C
0496
04F4
04DD
046F
0491
056B
058D
0362
FF4D
FBA3
FA4B
FADD
FB87
FB4C
FAC4
FAC5
FB23
FB32
FAEB
FAE5
FB44
FB7A
FB32
FAE9
FB22
FB7F
FB4C
FAB5
FAB5
FB8D
FC1B
FB66
FA6A
FB61
FF06
035A
05B0
0581
0494
048F
0534
0561
04DF
0486
04CE
0528
04FE
04A0
04B2
0519
0526
04BA
047D
04C7
0500
0491
0403
0459
054D
0509
023D
FDFE
FADF
FA3A
FB0C
FB8D
FB40
FAEE
FB1A
FB4C
FB0D
FAB6
FAE2
FB64
FB88
FB20
FACB
FAFD
FB59
FB59
FB30
FB6D
FBE1
FBB6
FAD7
FAB3
FCCF
00C3
0453
05B1
0538
0499
04C4
0531
051F
04B9
04A6
04FD
0532
04FF
04C3
04CF
04E5
04B2
0473
04A1
050C
04FD
045F
0421
04E4
0598
044B
0088
FC5A
FA4B
FABB
FBC2
FBA2
FAA0
FA1F
FA9E
FB4A
FB5F
FB1D
FB1E
FB55
FB4C
FB09
FB0D
FB68
FB8B
FB31
FAF3
FB5C
FBDC
FB7B
FA8E
FAE9
FDCA
0211
0531
05DF
0524
04B4
04FA
052E
04E9
04A8
04D8
0521
04FF
04A1
0496
04DC
04E1
0478
043B
04A6
053B
0529
048D
045E
04E8
04FA
0321
FF84
FC01
FA53
FA7C
FB2D
FB69
FB3F
FB25
FB2B
FB19
FAFD
FB16
FB51
FB51
FB08
FAEC
FB52
FBD3
FBC3
FB2D
FAD6
FB21
FB61
FAE8
FA71
FBB6
FF4B
0379
05CA
0595
046D
0418
04B7
053F
052A
04F2
0506
051A
04D2
0476
0479
04AE
0498
0456
048A
0537
0578
04CA
041B
04A3
05D5
057A
0251
FDE2
FAF5
FA8D
FB3C
FB55
FAD7
FAC4
FB4C
FB97
FB2E
FAB2
FAD4
FB4F
FB74
FB48
FB63
FBCA
FBC4
FB09
FA66
FAB3
FB7B
FB82
FAA6
FA85
FCAC
0093
03F8
0545
04FD
04A9
04EC
0539
0509
04B4
04C5
0516
0511
04A3
0460
04A0
04F5
04D9
0485
0498
050C
0529
04AC
0463
0500
05B0
0494
0109
FCCE
FA5D
FA62
FB5A
FBA6
FB37
FAF0
FB15
FB21
FADE
FACE
FB46
FBC0
FB9D
FB1C
FAFE
FB4F
FB54
FAD6
FAA2
FB4C
FC01
FB8B
FA5D
FAA0
FDAB
0218
051D
0588
04AE
045C
04C3
04F1
049B
0478
04F0
0563
0526
0492
047B
04EC
0521
04CB
048F
04EF
0557
04EF
0418
0419
0526
0586
036D
FF56
FBC4
FA90
FB1B
FB89
FB20
FABA
FB17
FBB4
FBA8
FB0C
FAC4
FB22
FB7C
FB4B
FAF4
FB19
FB7E
FB65
FAD2
FAAE
FB5D
FBF0
FB6F
FAA8
FBA6
FF28
034E
057F
0536
043D
0440
04FE
0535
04A2
0430
0477
04E7
04CB
0469
0483
0514
0553
04E9
0478
049E
04FB
04D8
0465
047B
0513
04B2
0215
FE07
FAE5
FA2F
FB22
FBF9
FBEB
FB8F
FB84
FB9C
FB71
FB2C
FB3B
FB8B
FB93
FB2C
FACC
FAD5
FB0D
FB16
FB16
FB5F
FBAE
FB5F
FAA3
FADC
FD32
00F5
0410
0523
04C1
045B
0481
04B1
048B
0476
04CA
051B
04D3
043A
042B
04D0
0552
0505
046A
0470
0508
0539
049F
0427
04AB
0562
0471
0136
FD45
FAD5
FA88
FB2E
FB81
FB66
FB63
FB83
FB5E
FAF3
FACE
FB38
FBB0
FB95
FB0F
FADC
FB45
FBB3
FB82
FAF0
FACF
FB5F
FBD5
FB5D
FA57
FA3C
FC30
FFC4
033B
0515
0537
04AF
047F
04C7
0507
04E8
049C
0483
04A7
04C5
04AF
048B
0493
04C6
04F9
0518
052E
052C
04E2
045F
0424
04B0
05A8
05C0
03D3
0032
FC9F
FAD0
FAEA
FB96
FB88
FAC2
FA47
FABB
FBA1
FC09
FBAC
FB20
FB01
FB43
FB6D
FB50
FB26
FB22
FB25
FB12
FB1F
FB7D
FBCD
FB6C
FA77
FA31
FBEB
FF7E
0326
0528
0560
0508
051B
0564
0531
0485
0421
0479
0517
0539
04C9
0467
0489
04E8
04F9
04B5
0495
04CA
04EA
048F
0417
0455
0553
05CA
0436
008F
FC9F
FA6E
FA5F
FB24
FB62
FB0C
FAF3
FB63
FBBE
FB6F
FACE
FAAF
FB3A
FBB9
FB97
FB24
FB0D
FB5D
FB7C
FB2E
FAFD
FB66
FBED
FBA3
FA9B
FA58
FC4E
001D
03B8
0560
0531
0499
04A0
0509
051B
04BD
047C
04B1
0504
04EE
0470
040E
042A
049A
04F6
0515
051A
0513
04D9
0469
0435
04B3
058A
057B
0373
FFD4
FC5E
FAAF
FAD0
FB6D
FB65
FADC
FAA8
FB0D
FB74
FB56
FB03
FB23
FBB5
FC03
FB97
FAEB
FAC5
FB30
FB78
FB33
FAD3
FAF3
FB5B
FB45
FAA5
FAAA
FC8F
0011
0376
0538
0558
04FB
04F6
0527
0519
04D2
04B7
04DB
04E7
04A2
0459
0475
04E0
051A
04E4
049A
04B2
0516
0538
04D9
0476
04B5
056B
056C
039B
0024
FC92
FA87
FA54
FAF0
FB27
FAC4
FA73
FAB1
FB37
FB75
FB58
FB4C
FB7F
FB9B
FB50
FAE5
FAE0
FB3E
FB6E
FB28
FAE8
FB3A
FBC0
FB8D
FA9D
FA64
FC64
004B
03F6
058F
0544
04B3
04E9
0579
0582
04FA
0498
04B7
04F1
04CF
047D
0475
04C1
04EF
04C7
049B
04C1
04FC
04D0
0450
0438
04F6
05CF
0558
02DB
FF2C
FC01
FA7D
FA76
FAF9
FB49
FB4C
FB37
FB24
FB0C
FAFE
FB19
FB54
FB70
FB47
FB0E
FB1B
FB6D
FB9F
FB68
FB12
FB24
FB9F
FBD4
FB3E
FA6E
FAD1
FD46
010D
0447
05A2
055A
04B2
0497
04F4
0535
051A
04E4
04DA
04EF
04F0
04D7
04C4
04BF
04A5
0471
045E
049C
04EE
04E1
0469
0422
0496
0551
04FB
02A5
FEF1
FBB7
FA5D
FAA7
FB3F
FB33
FABC
FA96
FAF3
FB5A
FB5F
FB28
FB1E
FB53
FB79
FB63
FB3F
FB4A
FB75
FB89
FB82
FB97
FBC8
FBB6
FB28
FAA6
FB48
FDAA
0119
0405
0552
053D
04DE
04F2
054D
0562
0510
04B7
049A
048E
045B
042F
0464
04E4
0529
04E5
047B
0479
04C5
04BA
0424
03C3
045E
0570
0548
02C7
FEC9
FB74
FA35
FAA1
FB4B
FB61
FB1F
FB04
FB10
FAFC
FAD6
FAFD
FB8A
FC09
FBFC
FB6F
FAEB
FAD2
FB0A
FB44
FB73
FBBA
FBFA
FBC0
FADF
FA19
FAC9
FDA0
01AC
04E7
05F5
0548
0478
0489
0517
0538
04CA
0481
04CC
0535
050F
0475
042B
048D
0514
0518
04B8
048E
04B9
04B9
0452
0427
04DA
05C8
0547
026D
FE54
FB30
FA36
FAB4
FB36
FB23
FAF3
FB1F
FB70
FB67
FB05
FAC5
FAE5
FB1D
FB15
FAF0
FB11
FB79
FBAD
FB60
FAF3
FB0D
FBAC
FBFA
FB58
FA71
FAE9
FDAC
01BC
04E7
05CE
050C
044B
0472
0503
0523
04CC
04AC
0515
058D
0586
0521
04E9
0500
04FB
049B
043F
045D
04BA
04B3
0436
0413
04DC
05C4
0515
020E
FDF2
FB04
FA61
FB2F
FBCE
FB89
FAEE
FABE
FAF7
FB12
FAD4
FA96
FAB0
FB01
FB21
FAFD
FAE2
FB0D
FB4D
FB58
FB4B
FB82
FBF9
FC11
FB5D
FA89
FB1B
FDE9
01F2
050E
05E6
051A
0457
0481
0514
0530
04D3
04AF
0511
0575
054E
04D1
04A5
04F3
0537
0510
04C8
04D3
0501
04BD
040C
03CC
0492
057C
04C4
01B0
FD98
FABB
FA20
FADD
FB6B
FB47
FB09
FB3D
FB9B
FB87
FAFF
FAA0
FAD1
FB43
FB65
FB26
FAFF
FB3B
FB8F
FB85
FB33
FB22
FB81
FBC0
FB55
FACC
FB93
FE71
0260
0542
05E9
0516
0471
04B1
052D
051D
04A9
0489
04E5
0527
04E6
0486
049B
0506
0518
0499
0427
045A
04E1
04F5
047D
0447
04D6
0553
043D
0127
FD6E
FAFF
FA85
FB0E
FB56
FB11
FAD8
FB19
FB83
FB86
FB17
FAB8
FACD
FB2B
FB6A
FB6D
FB68
FB70
FB59
FB11
FAF6
FB61
FBFC
FBEB
FAF2
FA36
FB61
FED3
02EA
0579
05C9
04FE
0492
04D3
0510
04DA
0492
04B5
0510
051A
04C7
0496
04D5
0522
04F8
0475
043B
0492
04F9
04CE
0435
0407
04AE
055C
049D
01CD
FDEE
FAE7
F9E3
FA6E
FB27
FB34
FADB
FAD3
FB3C
FB8E
FB61
FAFB
FAE4
FB2E
FB6B
FB56
FB2A
FB2F
FB48
FB35
FB20
FB6F
FC07
FC24
FB5A
FA8E
FB64
FE77
026F
052C
05BF
0515
04A6
04F4
0565
0559
04EC
04A5
04B5
04DB
04DA
04CD
04E6
050E
0506
04C8
049B
04AC
04C2
0484
0419
0423
04DC
055F
043E
010D
FD2F
FAB2
FA60
FB1D
FB5D
FAD8
FA7D
FAED
FB8F
FB7C
FACE
FA79
FAF0
FB86
FB6C
FADD
FAC5
FB66
FBED
FB9D
FAEB
FAE4
FBA3
FC14
FB76
FAB1
FB9A
FED9
02F0
0599
05EF
0506
0474
04B4
0517
04F5
0488
0480
050A
0590
057F
04F2
0487
048E
04C0
04BD
0495
048E
04A7
0497
0465
048F
053D
0582
03F9
0063
FC64
FA1F
FA2B
FB32
FB99
FB2E
FAE4
FB47
FBC9
FBA7
FB00
FA9D
FAD4
FB2A
FB1F
FAE6
FB03
FB73
FBA6
FB5A
FB0D
FB4C
FBC7
FBA1
FABD
FA5A
FBFC
FFA5
038D
05B6
05BE
04F6
04C0
052E
0562
04EA
0458
046A
0500
0550
04FB
0488
04A1
0521
0554
04F8
049A
04BA
0501
04C1
0417
03F5
04BF
0555
03FD
006B
FC6B
FA35
FA50
FB59
FBBD
FB44
FAC6
FADA
FB2F
FB30
FAD8
FAA3
FAD5
FB2E
FB55
FB49
FB42
FB4E
FB42
FB15
FB07
FB4E
FBA9
FBA0
FB38
FB55
FCFC
002F
0397
0591
05A5
04D3
0467
04AD
04F3
04B4
044D
0473
0526
05A5
056F
04EA
04D1
052F
0556
04E3
0451
0452
04D0
0510
04C5
0480
04B8
04BF
0340
FFF3
FC4C
FA2D
FA12
FAD7
FB2F
FAF3
FAD4
FB2C
FB97
FB9D
FB52
FB16
FB09
FAFF
FAED
FAFC
FB30
FB41
FB02
FABB
FAE7
FB7D
FBDA
FB7D
FAD1
FB07
FCFB
0055
03A9
0594
05CD
0536
04E4
051D
054F
04F9
0463
043C
04B1
052D
0525
04CD
04BC
0505
0524
04DF
04AB
04EE
0532
04BC
03CD
039A
049C
056E
0410
0052
FC4F
FA3E
FA49
FAE2
FAE4
FA9B
FAC4
FB51
FB99
FB64
FB26
FB32
FB43
FB06
FAB3
FAB9
FB1C
FB73
FB73
FB3A
FB0B
FB16
FB70
FBFE
FC48
FBCC
FAD6
FAC3
FCD2
009B
041E
05A6
055A
04A5
047C
04B4
04D1
04D1
04ED
050D
04F4
04C6
04E0
0533
0544
04EE
04AA
04CF
04FF
04C0
044A
0439
0486
0483
0408
03E4
04A1
052A
03AC
FFEC
FBF8
FA0E
FA56
FB35
FB6F
FB30
FB1C
FB35
FB25
FB00
FB23
FB73
FB71
FB0D
FAD9
FB20
FB6E
FB4B
FB06
FB2D
FBA2
FBCF
FBA9
FBB4
FBF9
FBB0
FAA6
FA57
FC94
00FD
04D3
05E4
04E4
042F
04CB
059B
0567
0495
0455
04DB
0541
0500
049D
04B8
0519
0527
04CE
0463
0415
03F0
0429
04CF
054C
04F8
0432
0435
0548
05B4
037C
FF05
FB1A
F9E8
FAC8
FB8F
FB4E
FADF
FB09
FB63
FB41
FAE8
FB04
FB6F
FB62
FACC
FA93
FB3C
FC1E
FC56
FBF6
FB97
FB46
FABA
FA4A
FAB5
FBC0
FC11
FB1B
FA86
FC8F
0102
0501
0633
0540
047B
04D7
054D
04F2
0457
046F
0510
0549
04DF
0481
049B
04B9
0476
0428
0442
048F
04AE
04CC
0537
0588
051D
0457
046B
0579
059A
02ED
FE46
FABA
FA27
FB48
FBB9
FAFF
FA7F
FB05
FBAD
FB78
FAD3
FAD7
FB8F
FC00
FBAD
FB36
FB39
FB6E
FB55
FB1C
FB29
FB4E
FB20
FAE2
FB29
FBAA
FB67
FA65
FA79
FD52
0203
058B
0619
04E2
0440
04D6
057A
054C
04C8
04A5
04B9
0484
042D
0445
04BF
04EC
0496
0454
0496
04FD
0511
0508
0537
0541
04B7
042B
04A8
05D7
059D
0271
FDA5
FA52
F9F0
FAFA
FB3C
FA85
FA35
FAE5
FBAD
FBAE
FB48
FB4B
FBB2
FBD9
FB97
FB69
FB85
FB81
FB20
FACB
FADB
FAFB
FACB
FAA9
FB15
FB9C
FB4F
FA75
FAE0
FDE4
025E
05A3
0652
0582
04F8
051A
052C
04E5
04BA
04E3
04EC
0486
041E
0434
049A
04C5
04B2
04D1
0526
0537
04EA
04D5
053D
0572
04E5
0445
04A4
058A
04E7
0189
FCF5
FA0A
F9EA
FB15
FB98
FB30
FACF
FAE5
FB04
FAF0
FB07
FB7B
FBD6
FB9F
FB18
FAD4
FAEA
FAFD
FAF7
FB24
FB77
FB77
FB19
FB09
FB97
FBE8
FB27
FA38
FB3D
FEFC
0382
0601
05C1
048A
0435
04CB
053E
052A
0503
050F
0509
04D5
04C6
0502
0525
04E4
0497
04BC
051E
0516
049E
0467
04BC
04F9
04A3
0457
04D7
0573
0469
0112
FD0E
FAA5
FA66
FAFB
FB19
FAD0
FAC2
FAF4
FAFF
FAE5
FAFB
FB35
FB2E
FAEB
FAE9
FB50
FB97
FB50
FAE8
FB09
FB7C
FB70
FAD6
FAA6
FB50
FBD7
FB44
FA82
FBAE
FF5B
037C
0592
055C
04AF
04EC
0598
05A2
050A
04A5
04C6
04FC
04F6
04E9
04FE
04FA
04B3
0473
0488
04C3
04CE
04D1
0525
057C
051C
042A
03E8
04F0
05CF
0456
0055
FC20
FA1D
FA59
FB15
FB21
FADB
FAEA
FB1D
FB05
FAD9
FB11
FB71
FB59
FAD1
FA9E
FB15
FB8D
FB5A
FACD
FAB3
FB1D
FB5B
FB35
FB3C
FBA7
FBB4
FAED
FA81
FC3F
0033
042B
05F2
0589
04A6
047B
04BD
04C4
04A8
04CD
0515
051F
0500
0510
0538
050E
04A1
0487
04F1
053F
04EA
046B
048F
0526
0534
0496
0467
0535
0592
038D
FF60
FB9B
FA57
FB01
FB86
FB02
FA6C
FABB
FB7F
FBC1
FB73
FB39
FB47
FB31
FAD2
FA9A
FACE
FB19
FB1C
FB01
FB1C
FB3B
FAFC
FAA4
FAE3
FB99
FBBB
FAF1
FAA7
FCA3
00AA
046F
0600
059B
04E0
04B7
04CD
04B3
04A6
04DD
04F6
049A
042F
0452
04D8
050D
04D1
04C1
0532
0599
0565
04EB
04E4
0535
0518
0484
0470
0530
054B
0300
FEB5
FAF3
F9BF
FA9A
FB8B
FB83
FB12
FAFF
FB32
FB3D
FB34
FB64
FBA0
FB80
FB1A
FAEC
FB19
FB45
FB40
FB4F
FB8F
FB8D
FAFD
FA73
FABA
FB76
FB6D
FA7F
FA79
FD16
018F
051A
05E9
04EA
0439
0497
051A
04F4
048B
048D
04E0
04FD
04EB
0515
0575
0586
051A
04A2
0484
0496
0485
0470
0498
04C6
0499
045E
04D1
05B5
0569
02A7
FE61
FB17
FA4E
FB33
FBF3
FBC4
FB3C
FB09
FB22
FB40
FB5B
FB6B
FB2C
FA97
FA3C
FA9B
FB55
FB9B
FB46
FAFB
FB2C
FB74
FB5F
FB3E
FB8D
FBDF
FB4E
FA38
FA92
FDA3
0213
0515
056C
047F
043F
04DC
0525
0498
040C
0452
0508
0553
051D
04F1
0500
04F5
04AA
046D
0475
048D
048E
04B5
052A
057C
052B
049C
04AF
0543
04CE
0223
FE2C
FB28
FA4F
FAD2
FB3C
FB21
FB13
FB62
FBAF
FB9E
FB5D
FB30
FB07
FAD6
FAE2
FB4C
FBAA
FB8D
FB39
FB4E
FBC3
FBD7
FB3A
FAA6
FACD
FB2B
FAC8
FA1F
FB16
FE97
02F2
057B
0578
0496
0486
0521
054A
04CB
0476
04B4
04F2
04BC
0482
04C8
0530
04FE
044E
03F7
0455
04DA
04FB
04E7
04FC
050B
04C2
048F
0519
05CD
04E1
0172
FD10
FA4B
FA06
FAE0
FB3C
FAFF
FB01
FB78
FBBC
FB71
FB08
FAFD
FB2A
FB3D
FB4C
FB7D
FB88
FB2B
FAC5
FAE7
FB5E
FB60
FACE
FA8E
FB35
FBE9
FB83
FAA2
FB6F
FEE5
0335
05AE
05B4
04F7
04F9
0570
0562
04D0
0487
04BC
04CF
047E
0461
04DC
055B
0533
04B3
04A1
04F9
050A
04AE
0492
0502
0548
04C4
0423
0471
051E
0424
00A8
FC83
FA51
FA80
FB42
FB23
FA98
FAB5
FB65
FBAC
FB42
FAE7
FB19
FB64
FB45
FB02
FB09
FB1D
FAD0
FA75
FABB
FB86
FBEA
FB8A
FB27
FB64
FBA8
FB1C
FA89
FBEA
FFC5
03F5
05E7
0574
049F
04CB
0565
0554
04B5
0470
04B6
04DC
049A
047B
04D8
0531
050B
04C5
04F0
0546
051E
049A
0486
0505
0539
04A9
043A
04CD
055E
03C7
FFAB
FB81
F9EA
FAC1
FBBA
FB6F
FAA6
FA9C
FB2C
FB60
FB0C
FAE2
FB24
FB3F
FAE2
FAA3
FB07
FB97
FB9D
FB43
FB3C
FB8A
FB83
FB0C
FAE6
FB62
FB9C
FADB
FA41
FBF2
003C
04A3
067A
05C3
04A9
04A5
052F
053B
04DB
04D2
053F
057E
0544
0502
0510
0529
0503
04DC
04F1
04EC
0475
03FE
0435
04E6
0522
04AE
0479
0511
0542
033E
FF21
FB53
F9EF
FA93
FB57
FB52
FB1D
FB4B
FB6B
FB00
FA86
FAC3
FB74
FB8B
FABA
FA00
FA4A
FB34
FBB1
FB79
FB21
FB14
FB28
FB2F
FB4A
FB71
FB44
FAD0
FB27
FD68
0126
0468
05A9
0553
04E7
0515
0553
0512
0495
046F
04B0
04F8
051A
0532
053F
0513
04B8
0486
049D
04B5
04A4
04A8
04E8
0501
049E
0444
04CE
05EB
05D8
0335
FEE4
FB61
FA35
FA99
FAE3
FA8F
FA5C
FAC5
FB50
FB6B
FB42
FB53
FB91
FB7D
FB08
FAC1
FB09
FB82
FB99
FB5A
FB45
FB7A
FB92
FB48
FAEA
FAE9
FB29
FB1F
FA9A
FA3D
FB0C
FD79
00E6
0405
05B8
05D5
0527
04B2
04D2
051D
0511
04BA
047F
048F
04B5
04BB
04B2
04BF
04D2
04C3
04A6
04BA
04FF
052D
0523
051C
053D
053B
04CE
044D
0468
050A
04FD
030C
FF85
FC2D
FA90
FAA4
FB32
FB4E
FB0D
FAF1
FB1C
FB51
FB64
FB68
FB69
FB52
FB1C
FAFE
FB29
FB75
FB87
FB40
FAEB
FADE
FB0E
FB2D
FB1C
FB1B
FB5F
FB9C
FB4C
FA9B
FAB5
FCD0
00AB
0461
0603
0568
042C
03E2
0499
0536
050C
048B
0468
04AC
04DC
04C9
04C0
04F3
052A
0525
0505
0502
04F9
04A0
0426
0422
04B5
052F
04ED
0457
0468
0531
054D
0353
FF8E
FBF6
FA46
FA76
FB38
FB8B
FB80
FB8D
FBB9
FBA5
FB35
FAC8
FAC3
FB17
FB63
FB63
FB2E
FAFA
FAE0
FAE4
FB0E
FB56
FB86
FB60
FAFC
FAD5
FB40
FBDD
FBDC
FB14
FAB1
FC45
FFF9
03F3
05F7
0590
045E
0427
04FB
058F
051F
0457
0442
04E7
056C
0550
04FC
04F8
0527
051A
04D7
04CF
0517
0535
04DE
047C
0498
04F8
04EA
0460
042B
04C4
053C
03FE
00BC
FD0A
FAD9
FA8D
FAFA
FB00
FAA4
FA80
FAB6
FAD6
FAB1
FAA2
FAF4
FB5C
FB59
FAF3
FAAF
FAD6
FB19
FB17
FAF3
FB15
FB77
FB9B
FB46
FAF1
FB30
FBC4
FBCB
FAFF
FA7A
FBCF
FF43
033E
05AD
05EE
052B
04E2
0565
05E9
05C8
054C
0524
056C
0591
052A
0484
043C
0478
04CB
04DB
04BE
04B8
04C9
04CB
04C7
04E0
04FA
04CA
046D
048B
0560
05E2
046B
00A6
FC58
F9D9
F9C4
FAA9
FAEF
FA85
FA5F
FAD3
FB2D
FAE4
FA74
FAA2
FB4C
FB9E
FB53
FB16
FB76
FC01
FBDF
FB0D
FA6C
FA90
FB0D
FB3A
FB28
FB59
FBB9
FB91
FABB
FA59
FBDB
FF54
032F
05A6
063F
05D3
055E
0530
0524
051C
0524
0530
051D
04E4
04B6
04BF
04E7
04E9
04B0
047B
0492
04E4
051B
0508
04E4
04FA
0527
04F8
0469
0427
04B3
054C
044B
00FF
FCD1
FA1F
F9DD
FACB
FB20
FA90
FA2F
FAAE
FB6C
FB80
FB04
FAC1
FAF9
FB1F
FADA
FA9D
FAF7
FB98
FBBA
FB3D
FAE0
FB21
FB8B
FB77
FB1B
FB33
FBBB
FBC7
FAEC
FA50
FBA5
FF21
0303
0554
05C4
057F
0581
05AC
057A
04FB
04C1
0502
0553
054D
0512
0509
0534
0531
04D7
0482
049B
0503
0532
04ED
048B
0473
0489
045F
0400
0414
04F0
05AE
04B5
0172
FD49
FA6F
F9DA
FA91
FB06
FAC7
FA86
FAC8
FB2D
FB22
FAC9
FAB8
FB10
FB51
FB2C
FAFD
FB2F
FB7D
FB49
FA9E
FA4B
FAD3
FBA2
FBD0
FB67
FB47
FBCA
FC20
FB7B
FA8F
FB34
FE4A
0278
0564
0609
0565
0500
053C
056D
0523
04BF
04C3
050F
0522
04E6
04C5
04F7
052A
0507
04C6
04DD
053D
0555
04EC
0487
04AC
0502
04B9
03CF
035F
0432
0558
04CE
01BB
FD99
FACC
FA45
FAEC
FB3D
FAEC
FAB8
FB11
FB7C
FB5F
FADB
FA8D
FAB1
FAED
FAF2
FAEF
FB2D
FB83
FB80
FB1A
FAD0
FB00
FB58
FB4C
FAF1
FAF7
FBA7
FC46
FBF9
FB2C
FB8B
FE32
0230
0539
05EE
0508
043E
045D
04D4
04F0
04D3
0509
058B
05C4
056E
04F5
04D0
04DA
04AD
045B
0461
04D9
052C
04DE
044D
0445
04D1
051E
04A6
0410
0452
0517
04B1
01F9
FDEA
FAD9
FA22
FAF8
FBA9
FB88
FB32
FB42
FB70
FB29
FA8E
FA4F
FAB5
FB47
FB7D
FB66
FB60
FB70
FB4E
FB00
FAF9
FB6D
FBDE
FBB4
FB24
FB02
FB9C
FC26
FBB7
FAB7
FAD8
FD55
016B
04E6
062B
059C
04CA
04B0
04FB
04EA
0477
0443
049D
0517
0528
04E5
04CA
04F4
04FC
04AB
0462
0489
04EE
04FE
04A0
045B
0486
04BA
0478
0413
0458
052E
0520
02DE
FEF3
FB82
FA29
FA87
FB09
FAD9
FA7A
FAB3
FB66
FBD2
FBA2
FB3D
FB14
FB15
FAF8
FAD6
FB08
FB8E
FBE9
FBB8
FB3E
FB04
FB26
FB46
FB31
FB36
FB91
FBD5
FB62
FA8A
FAC6
FD3F
014A
04C2
060A
0582
04C8
04DE
0557
055E
04E5
0495
04CC
0532
054D
051E
04EF
04D3
049C
044F
043C
0489
04E0
04D6
0484
046B
04BD
050C
04E4
0488
04A7
0544
0535
032E
FF51
FB74
F98B
F9DD
FAFD
FB75
FB1F
FACB
FAEF
FB27
FAF8
FA9A
FAA0
FB1C
FB86
FB81
FB53
FB5F
FB8D
FB7C
FB28
FAF5
FB0C
FB1D
FAEE
FAD0
FB26
FB99
FB6A
FAB5
FAD9
FD1D
0102
0475
05D6
056C
04BE
04C4
052F
054B
050B
04EC
051C
053D
0503
04A6
048F
04BD
04D6
04AD
047F
0497
04DE
0509
0508
0517
054B
0553
04F6
048E
04B7
0557
0545
0350
FFAE
FC1B
FA4C
FA62
FB0D
FB20
FAAA
FA7D
FAE5
FB55
FB3C
FACA
FA9E
FAF5
FB68
FB88
FB5F
FB3B
FB2E
FB13
FAE9
FAE5
FB11
FB20
FAE8
FAC2
FB1E
FBB5
FBB0
FAD5
FA52
FBC3
FF57
034E
059D
05DB
054C
0525
055A
053F
04C5
048B
04E7
0566
057A
0531
04F8
04E8
04B9
046B
046B
04E7
0563
0549
04C5
048F
04E2
0529
04DD
046E
04C2
05CE
0626
0453
0082
FC99
FA79
FA5E
FB01
FB1D
FA9C
FA46
FA99
FB33
FB71
FB40
FB16
FB30
FB46
FB0F
FAC6
FAD4
FB33
FB6B
FB45
FB1C
FB49
FB8D
FB70
FB07
FAE4
FB1F
FB16
FA7B
FA4C
FBFD
FF9B
0355
0539
051D
0478
048A
0529
0579
0539
04EB
04E7
04F2
04C3
048D
04A8
0505
0531
04FC
04BA
04C7
04FC
04E3
0473
0435
048E
0525
0548
04E7
04B2
0517
054B
03E7
0091
FCC4
FA85
FA65
FB2E
FB75
FB1F
FB01
FB79
FBF3
FBCE
FB3B
FAE0
FAF7
FB27
FB2C
FB37
FB70
FB99
FB62
FB04
FAFC
FB4D
FB68
FAF8
FA82
FABC
FB83
FBD8
FB2E
FA7F
FB88
FEE3
0315
05D1
061D
0506
044B
049A
0542
0562
0500
04BE
04E1
050E
04E7
0495
046F
0478
0470
0450
0451
047F
0497
047A
047E
04EF
0576
0569
04D0
0491
0534
05C7
0499
0131
FD21
FA99
FA45
FAF8
FB3F
FADF
FA9C
FAED
FB6A
FB7F
FB29
FAD5
FAB7
FAAC
FAA7
FADF
FB6C
FBEE
FBE8
FB66
FB07
FB39
FBB2
FBD1
FB74
FB10
FB00
FB07
FAD4
FACC
FBF2
FEC8
026E
052F
05EF
051E
0429
0420
04E6
0599
0590
04F7
047B
0490
0504
054E
0522
04B2
046B
047E
04CB
0500
04EC
04A8
048B
04C3
0508
04E2
0452
0411
04B4
0593
04FB
01F5
FDB2
FAA5
FA14
FAF6
FB75
FB0B
FA99
FACC
FB31
FB0F
FA91
FA7E
FB07
FB89
FB8D
FB61
FB7B
FBB2
FB93
FB31
FB0F
FB5C
FBAB
FB8F
FB28
FAE4
FAF5
FB32
FB63
FB59
FAF3
FA6E
FAB4
FCC0
0057
03D6
05A4
05B2
0533
0510
0528
050A
04C7
04BE
04EF
04FF
04D6
04C6
04EE
04FC
04B9
0472
0483
04C4
04D7
04BE
04CB
0500
050F
04E7
04E1
0518
0512
0482
0416
04B2
05CF
0571
0265
FDFB
FADC
FA4A
FB20
FB93
FB27
FAA0
FA8F
FABB
FAD5
FB01
FB61
FBA0
FB6B
FB12
FB23
FB9E
FBEC
FBB3
FB3C
FAEA
FABA
FA80
FA60
FA9D
FB14
FB54
FB4E
FB65
FBA5
FB77
FAAA
FA5C
FC1F
FFFC
03F2
05E0
059B
04BC
0492
04EF
0507
04BE
049F
04DE
051A
050A
04DF
04D5
04CF
04A2
047E
04B3
051E
0547
0511
04DF
04EC
04FA
04D2
04B3
04DA
0500
04CD
04A5
052D
05F3
0542
020C
FDA2
FAAD
FA5B
FB4E
FB9E
FB17
FACE
FB31
FB87
FB42
FADD
FB01
FB71
FB76
FB04
FAC2
FAF3
FB1F
FAF6
FAE2
FB39
FB93
FB71
FB1E
FB3A
FB9F
FB95
FB10
FAE3
FB60
FB8E
FA9D
F9BE
FB3D
FF84
0411
0618
0583
047C
0488
0524
0538
04BB
0468
047F
049F
04A7
04E7
0561
0587
0519
04A8
04BF
050E
04FA
04A0
049D
0501
0533
04EB
04A5
04C4
04DE
047D
042A
04C3
05BF
051E
01C9
FD54
FA88
FA68
FB78
FBE4
FB83
FB4E
FBA7
FBF0
FBAF
FB3D
FB19
FB21
FAF8
FAB9
FACA
FB23
FB54
FB34
FB0E
FB16
FB13
FADF
FAC0
FAF8
FB32
FAF9
FA9A
FAE7
FBDB
FC42
FB66
FA97
FC0D
0027
0487
0670
059B
041F
03C9
046E
04E6
04D0
04AF
04CD
04DE
04B4
049F
04D5
0505
04D1
047D
0491
0504
053F
0508
04D3
04FC
0534
0517
04CC
04AA
048B
042B
03F6
04A5
05BC
054F
0215
FD66
FA3E
FA09
FB46
FBB3
FAF8
FA65
FABA
FB50
FB63
FB3A
FB79
FBF6
FBFA
FB68
FAF0
FB01
FB40
FB3B
FB11
FB03
FAE9
FA9E
FA89
FB08
FBA8
FBA9
FB29
FB1F
FBD3
FC32
FB5D
FA77
FBBE
FFAB
03F0
05F5
059E
04D4
04DE
0544
0526
04A7
047E
04C6
04F8
04DF
04D8
050B
0514
04BA
046D
04A2
0517
0541
0528
0537
0568
053D
04A1
042E
0446
046D
0413
03B4
0446
056F
053D
0259
FE00
FAEB
FA66
FB36
FB7A
FAE0
FA77
FAD9
FB68
FB60
FAEB
FABB
FAF4
FB1E
FAF4
FAC1
FADD
FB2E
FB63
FB5C
FB33
FB02
FAE5
FB07
FB6F
FBC4
FBB1
FB72
FB96
FC09
FBEE
FAEB
FA42
FBCE
FFC6
040D
0635
05E7
04D9
048E
04F1
052B
0511
0517
0553
055C
0512
04E0
0509
052C
04DB
0458
043F
049A
04DA
04C0
04A6
04C5
04C1
0461
0426
0487
0508
04D5
042D
043C
052C
0539
0296
FE07
FA7A
F9C7
FAD0
FB54
FAC3
FA54
FAD1
FB7F
FB6D
FAD3
FA98
FAF1
FB42
FB2A
FB03
FB2B
FB6C
FB72
FB55
FB51
FB50
FB30
FB2B
FB78
FBC1
FB98
FB43
FB75
FC18
FC1B
FB07
FA4B
FBF2
000C
0432
0615
05D0
0527
0524
0557
0527
04D3
04D6
0503
04E2
048E
0491
04F5
0521
04D2
048D
04C4
0510
04DE
0463
0454
04BF
04EC
0480
040B
0423
046F
0445
03E6
0440
0537
050B
0245
FDCB
FA50
F98C
FAA6
FB94
FB67
FACC
FAA2
FAE4
FB08
FAEF
FAEE
FB2A
FB6B
FB7D
FB75
FB79
FB82
FB77
FB55
FB27
FAFF
FB03
FB5E
FBEC
FC29
FBCA
FB4E
FB78
FC1F
FC2C
FB2D
FA7F
FC1C
0025
044C
0628
05A7
04BA
04C5
0554
055A
04D3
048C
04C8
0509
04F8
04DB
04ED
04E4
0485
0439
0489
052B
0542
04A3
0420
0457
04D4
04DA
047F
0455
0466
0446
0411
046C
0534
04DB
020D
FDB0
FA5F
F9AA
FA95
FB33
FAF2
FAA5
FAE6
FB58
FB7C
FB65
FB5A
FB4F
FB1B
FAEC
FB00
FB2D
FB1B
FAE9
FB12
FB86
FB99
FB1C
FAD6
FB60
FC16
FBF9
FB3B
FB09
FBB2
FC09
FB3A
FA82
FC13
0030
046C
0645
05BC
04C4
04B0
051F
0533
04DB
049D
04A9
04C2
04CD
04EF
0522
051F
04D9
04A8
04CB
0504
0501
04D9
04D2
04D9
04A9
045B
0458
04A5
04B7
0447
03F5
0478
0547
04B8
01DA
FDD5
FAE4
FA26
FACB
FB61
FB5E
FB26
FB12
FB06
FAE5
FAD6
FAF5
FB0D
FAF7
FAEE
FB2E
FB7B
FB67
FB00
FACB
FB04
FB40
FB1E
FAF6
FB50
FBE7
FBE8
FB44
FAEF
FB7B
FC10
FBA7
FAEF
FBEF
FF76
03B0
05F6
05B2
04AE
0498
053B
0573
0506
04B5
04E6
052F
0521
04E0
04BE
04B0
048F
047A
04A2
04D9
04D0
04AC
04D9
053D
0539
04A9
0444
0480
04CD
0482
041A
0490
0588
051A
0213
FDC9
FAE0
FA66
FB00
FB05
FA6E
FA32
FA92
FAF6
FB11
FB35
FB85
FB9F
FB58
FB2C
FB89
FC0B
FBFA
FB67
FB18
FB58
FB87
FB2F
FAC8
FAED
FB53
FB49
FAF2
FB22
FBE5
FC24
FB3B
FA69
FBC0
FF9B
03E1
062B
061D
053E
04EA
052D
0564
054C
0517
04F0
04CA
049C
0470
0449
0425
0422
0461
04B2
04B9
0471
0451
04A9
051A
050F
049B
046E
04C9
0510
04B9
0443
0498
0574
052A
0278
FE47
FAF3
F9E5
FA6A
FAEF
FAD5
FAA3
FACA
FB00
FAED
FAC8
FAF0
FB4C
FB81
FB8C
FBB6
FBFB
FBF9
FB8F
FB29
FB2A
FB5D
FB5A
FB33
FB4D
FB94
FB8B
FB36
FB3E
FBD0
FBF7
FAFF
FA07
FB3F
FF3C
03D2
063A
05FB
04F5
04D2
0559
058A
054B
0541
0587
058C
0516
0497
0471
0468
0433
040B
044C
04BE
04D6
0497
0490
04ED
0524
04DB
0483
0490
04A9
044F
03F4
0473
0574
0530
026F
FE47
FB2F
FA6B
FB05
FB62
FB12
FAA9
FA83
FA7B
FA7B
FAA9
FAF4
FB0D
FAF1
FB08
FB76
FBC7
FB83
FAF4
FAC9
FB1C
FB52
FB18
FAE2
FB1F
FB78
FB65
FB2F
FB89
FC4A
FC57
FB48
FA82
FBF3
FFB7
03A4
0581
0531
0463
0465
04FF
0555
0531
050A
0521
052E
04EF
04A6
04BC
052C
0580
0562
04FC
04B3
04B8
04E9
0509
04EB
0496
044E
045F
04BB
04E1
047C
0402
0440
0515
050D
02C7
FEBC
FB21
F9CC
FA80
FB86
FBB6
FB54
FB15
FB0F
FAEF
FAB4
FAA4
FAC5
FAE6
FB08
FB5E
FBCB
FBD7
FB52
FABA
FA9C
FAD6
FADF
FAB0
FAD0
FB61
FBD8
FBD3
FBAC
FBB6
FB83
FAB5
FA38
FBB7
FF7D
039C
05BC
0588
04A5
047D
04DB
04F1
04B8
04BB
0507
0526
04F3
04C9
04D4
04D5
04A9
049B
04E1
052C
0513
04C1
04B9
04F4
04E1
0462
0423
048B
04F9
04B1
041F
0456
054E
055D
0311
FF11
FBA9
FA79
FB02
FB9C
FB5C
FAB2
FA71
FAD4
FB6C
FBB4
FB87
FB2D
FB0D
FB42
FB83
FB85
FB51
FB30
FB44
FB63
FB5D
FB46
FB5B
FBA6
FBE7
FBD4
FB6E
FAFB
FACA
FAF2
FB44
FB5C
FAF7
FA6C
FAA1
FC63
FF8A
02EB
0533
05DC
056A
04CF
0494
0495
047C
0446
0438
0471
04BD
04E1
04EA
04FC
0503
04CA
0469
044E
04A5
04F4
04B9
0444
0461
0529
05B2
0551
0495
0480
050E
0544
04BD
0461
0501
05BA
04AA
014B
FD60
FB1B
FAEC
FB89
FBC2
FB88
FB5A
FB67
FB88
FBA1
FBB1
FBA5
FB5E
FAF5
FAB8
FAD1
FB1A
FB55
FB6A
FB55
FB18
FADD
FAE3
FB21
FB3A
FB03
FAC4
FAD0
FB0F
FB3F
FB71
FBCE
FC08
FB93
FAB5
FAE4
FD56
014B
0472
0540
0472
03D6
042A
04BC
04D7
04BA
04EF
055F
0576
0510
04AE
04BC
0500
04FF
04B5
048D
04C2
050E
0518
04EE
04E7
0529
0571
0563
050D
04DE
0501
0504
0475
03C6
03F2
0508
0582
03B5
FFE0
FC3F
FAC9
FB32
FBAA
FB33
FA8D
FAB9
FB6A
FB8D
FADF
FA41
FA6F
FB16
FB6E
FB4B
FB30
FB6F
FBB9
FB9B
FB28
FAD4
FAD7
FAFB
FB01
FAEF
FAE5
FADE
FAC5
FAB2
FAF4
FBA2
FC36
FBED
FACE
FA35
FBC3
FF87
038E
05AA
0584
04A3
047A
04FE
054D
052B
0528
0578
057F
04D3
0415
0426
04DF
053A
04BB
0412
0420
04C8
052F
04F3
04A0
04CC
0540
055B
0507
04D6
0520
057C
0548
0494
0435
04B4
055B
0497
0198
FD7D
FA7D
F9CA
FA8D
FB16
FAC5
FA62
FAC6
FBA4
FC07
FB9D
FB0D
FB00
FB63
FBB9
FBCC
FBAF
FB67
FAFB
FAB5
FAE1
FB57
FB92
FB58
FB10
FB30
FB91
FB97
FB0D
FA7E
FA87
FB03
FB36
FAC2
FA4F
FB1A
FDCD
01AF
04F5
0639
05B0
04CE
04A6
04FB
0501
049D
0470
04BB
04EB
0484
0407
044B
0529
0585
04DC
0411
0439
0515
0574
04E4
043B
0459
0503
0558
0513
04C6
04DF
050E
04E2
049A
04CC
0561
054F
0395
0050
FCC7
FA7A
F9FC
FAA6
FB4A
FB4E
FAFC
FADB
FB05
FB33
FB41
FB4E
FB5E
FB40
FAEA
FAC4
FB31
FBE9
FC27
FBAC
FB11
FAEE
FB14
FAFB
FAAA
FAA3
FB05
FB4D
FB20
FAED
FB4D
FBFA
FBF2
FAED
FA2F
FB71
FEF3
02FF
056E
0594
0496
040F
048A
054C
056A
04E8
047E
0498
04DF
04DD
04AA
04A3
04CC
04CC
0490
0484
04EE
055D
0534
0491
043F
0498
050E
050A
04C4
04CB
0509
04EE
046F
0450
04FF
05A8
04CD
01EB
FE2C
FB57
FA49
FA90
FB34
FB86
FB6B
FB2A
FB0E
FB24
FB41
FB53
FB66
FB6E
FB3F
FAEE
FAE4
FB59
FBDA
FBBD
FB0C
FA9B
FAF7
FB9A
FB9A
FAFA
FAA5
FB0A
FB7E
FB4D
FAD7
FAEA
FB67
FB5B
FAA6
FAAA
FCD8
00CC
046D
05FE
05A9
04DF
04AC
0507
0560
0561
050C
0498
044A
044F
0491
04D0
04E1
04C8
04AC
04AF
04D4
04F5
04E5
04A9
0481
04AC
050F
0546
0519
04C9
04B5
04C6
04A6
0474
04C3
0591
05B0
03CC
000F
FC48
FA43
FA38
FAEE
FB36
FAED
FAA4
FAB1
FAEE
FB1E
FB3C
FB5B
FB6B
FB4E
FB0D
FAEC
FB30
FBBD
FC02
FB92
FABC
FA54
FAB5
FB58
FB92
FB63
FB4E
FB73
FB68
FB02
FAC8
FB2C
FBA8
FB64
FABE
FB67
FE65
028C
0586
0639
059B
0530
0563
0594
0548
04C4
0488
04AD
04F3
052F
0559
0559
051A
04BB
0477
046B
048E
04C6
04E7
04CD
048E
0470
0495
04C8
04CD
04B2
04A6
049C
0468
043B
048E
053B
0505
02B8
FED6
FB77
FA2F
FA83
FAE1
FA9F
FA5B
FA9D
FB02
FAF2
FA9E
FAB3
FB3A
FB7E
FB16
FA8D
FA9D
FB31
FB8E
FB5B
FAFD
FAF7
FB49
FB97
FBA3
FB82
FB61
FB4A
FB29
FB0D
FB32
FBB3
FC2D
FC07
FB3E
FAE2
FC58
FFD7
03C6
060B
0608
0509
04A1
050D
057A
0569
0537
0558
059E
058D
0513
049F
0487
04A7
04B7
04B7
04D6
051B
054E
0541
04F6
0497
045A
0464
04A0
04CE
04BA
046C
0413
03EA
0424
04B6
0501
0405
014B
FDB5
FAFC
FA2A
FA9C
FAE8
FA87
FA2E
FA7C
FB09
FB13
FAB3
FAAC
FB39
FBA6
FB56
FAB2
FA9C
FB37
FBB7
FB77
FAD0
FA91
FAEC
FB52
FB53
FB23
FB29
FB5E
FB68
FB36
FB32
FBA4
FC1E
FBDE
FB03
FAF8
FD22
011E
04C4
0637
05B2
04FD
0545
05FD
0608
055B
04E0
0506
052D
04C6
043F
0459
04F4
053C
04E1
048B
04D8
0576
0598
0512
048B
0491
04E9
050F
04F4
04EB
0501
04E1
0474
0436
04A4
056B
0557
0356
FFA8
FBF8
F9FC
F9F1
FA96
FAB0
FA44
FA2C
FABC
FB4B
FB35
FACC
FAD6
FB59
FB8F
FB1D
FAA7
FADC
FB6B
FB81
FB05
FAB2
FAF8
FB5D
FB45
FADE
FAD1
FB33
FB64
FB0D
FAB8
FAFF
FB8F
FB84
FAC7
FA7A
FBF3
FF4E
032A
05BB
0637
0561
04AD
04E2
058E
05CC
0559
04C3
0494
04AB
04A1
0489
04CA
0554
0582
0514
04A6
04DC
055F
0555
049F
041B
0469
0512
053D
04E7
04D3
0547
0590
051E
0485
04B2
0551
04C0
01F0
FDDF
FAD2
FA15
FADE
FB6E
FAFC
FA48
FA59
FB29
FBCD
FBAC
FB24
FAEB
FB23
FB55
FB34
FB02
FB0E
FB2C
FAFB
FA9B
FA95
FB14
FB8D
FB7E
FB20
FB03
FB2F
FB2B
FADB
FACA
FB54
FBDA
FB69
FA40
FA14
FC61
009F
048D
064C
05F2
0507
04C5
051C
054C
04FE
0499
0489
04A8
0497
046F
04A5
053F
0599
0536
048A
0478
051F
0596
052E
0474
0478
0540
05BA
0549
04A2
04AC
051A
04F1
0436
041D
0530
0605
0494
00B1
FC88
FA5F
FA6C
FB26
FB42
FAC8
FA63
FA6B
FAB6
FB02
FB34
FB51
FB60
FB6F
FB82
FB82
FB4A
FADC
FA77
FA68
FABE
FB35
FB71
FB48
FAEB
FABE
FAEA
FB1D
FAFB
FAB6
FAE2
FB83
FBC7
FB14
FA44
FB1F
FE63
02A5
0587
060B
0543
04C4
04FE
0551
0549
0525
0530
053F
0500
0492
0468
04AE
050B
0509
04AA
045E
047E
04F4
0560
057C
0549
04F6
04B3
04A1
04C8
0510
053A
0506
0492
0467
04DF
056B
04C2
0221
FE53
FB27
F9DD
FA24
FABC
FADE
FAC4
FAF0
FB5F
FB9C
FB70
FB28
FB1F
FB49
FB57
FB20
FAD7
FABD
FAD4
FAE1
FAD3
FAE2
FB38
FB95
FB8D
FB26
FAEC
FB3D
FBBC
FBBC
FB28
FAB2
FADD
FB50
FB78
FBB5
FD33
0051
03C8
05D5
0604
055D
04F5
04E0
04AF
0468
0478
04E1
0517
04CA
0468
047F
04EC
0522
04F8
04D8
050A
0548
0531
04D3
0495
049D
04A7
0480
0466
04AF
0533
0556
04CA
041A
0424
04FE
057D
0426
00BE
FCD4
FA6D
FA25
FAD9
FB28
FAE4
FAC9
FB2B
FB7C
FB3F
FAD6
FAFF
FBB9
FC2F
FBD3
FB1A
FACB
FB00
FB2F
FB03
FAC4
FAD3
FB23
FB66
FB82
FB8E
FB88
FB50
FAF3
FAC2
FAEB
FB35
FB53
FB4F
FB64
FB88
FB70
FB37
FBAB
FD95
00B7
03B7
054A
0550
04C5
0496
04CD
04E2
04A5
0476
04B6
0537
0576
0538
04CA
0495
04B3
04ED
050A
0503
04E8
04CF
04D1
04FB
0535
054F
0538
0508
04CE
0486
044F
046D
04E4
052F
04C1
03DF
038F
045F
055E
04D1
0213
FE63
FBA4
FA9A
FAA3
FAE5
FB26
FB7F
FBBC
FB81
FADD
FA5B
FA63
FAC7
FB20
FB4E
FB77
FBA1
FB9B
FB53
FAFF
FADB
FADE
FAD6
FABB
FABC
FAFA
FB55
FB8F
FB98
FB98
FBA1
FB90
FB4F
FB1C
FB4A
FBB8
FBCE
FB46
FAE8
FC13
FF34
02EE
053A
0569
04AE
048C
052F
059D
054A
04CC
04E2
0550
0541
0485
03E3
0408
04AE
0517
0513
050B
053C
055B
0522
04CC
04BB
04E1
04DD
0496
045F
0474
0499
0488
0467
0480
04A9
046D
03E0
03C3
0477
0506
03D8
008E
FCB8
FA74
FA59
FB30
FB82
FB1A
FAC2
FAF3
FB51
FB59
FB16
FAF3
FB11
FB30
FB1D
FAF7
FAED
FAFF
FB10
FB1C
FB29
FB24
FB05
FB00
FB52
FBCC
FBE9
FB79
FAFA
FB02
FB72
FBA6
FB6F
FB58
FBC6
FC27
FBA1
FA8B
FA98
FD15
013A
04C0
060F
0598
04E7
04E1
0536
054A
0517
04FE
051E
0531
050A
04DA
04DC
0502
050E
04F0
04CD
04BD
04B5
04A9
04AE
04D0
04EA
04CE
0494
048B
04C3
04E6
04AD
045F
0477
04DB
04D6
041B
0378
03F1
051D
0506
0234
FDA3
FA14
F944
FA54
FB27
FADD
FA58
FA93
FB3E
FB6C
FB08
FADD
FB4E
FBB2
FB58
FA98
FA60
FAEC
FB7D
FB6E
FB00
FAE0
FB2B
FB6D
FB62
FB52
FB80
FBBA
FBB3
FB8C
FB94
FBBC
FBAB
FB6A
FB72
FBE5
FC20
FBA0
FB2C
FC5E
FFBC
03B3
05FD
05EF
04ED
049B
0527
0597
055D
04F4
04FE
0556
0568
0510
04BB
04B4
04CA
04B1
0484
048A
04C4
04E8
04CB
0492
046A
0452
043E
0440
0462
0478
0455
042E
0461
04DA
04FA
0464
03AC
03C7
04AD
04F6
0330
FF8D
FBEE
FA1A
FA39
FB0D
FB6F
FB38
FAE2
FAC0
FAC6
FAE0
FB18
FB5E
FB75
FB46
FB15
FB2D
FB7B
FBA4
FB8B
FB71
FB8D
FBA9
FB7A
FB1E
FB08
FB5D
FBAE
FB8D
FB31
FB25
FB7B
FBB3
FB81
FB55
FBA8
FC1F
FBE4
FB0F
FB18
FD5C
0152
04C7
0606
0571
04B7
04CE
053C
0534
04C3
0489
04B1
04C9
0487
0443
045F
04AA
04B0
0477
0482
04FE
056D
0548
04BE
0468
0472
0478
0443
042E
048E
050E
0517
04AC
0472
04B6
04F6
04B4
045C
04B0
0556
04B9
01CC
FDA5
FAA6
FA1D
FB20
FBDF
FB9A
FAFC
FAD3
FB15
FB49
FB4C
FB5B
FB83
FB82
FB3E
FAFC
FB0B
FB5A
FBA1
FBBC
FBB7
FB94
FB48
FAF5
FAEB
FB44
FBAE
FBCD
FBAF
FBA6
FBBD
FB96
FB0A
FA8E
FAB3
FB4B
FB7C
FAEF
FA9A
FBF3
FF44
030E
0565
05B6
050C
04B9
050C
0571
0570
0526
04E8
04C4
049C
0479
047E
04A0
04A3
0475
044D
0458
0479
0480
0477
0487
04A3
0491
0459
045E
04CC
0533
0503
0459
03FE
045C
04E7
04E7
0497
04E0
05D2
05F4
03B0
FF5E
FB4D
F998
FA2C
FB3E
FB6D
FAED
FAAE
FAF9
FB4D
FB4B
FB30
FB54
FB93
FB9E
FB81
FB97
FBE7
FC09
FBBC
FB49
FB21
FB41
FB4C
FB31
FB47
FBB0
FC09
FBEB
FB8A
FB5E
FB66
FB25
FA88
FA3D
FAC4
FB88
FB80
FAD3
FB24
FDC3
01E0
0524
0616
0562
04B7
04D3
0524
04FB
0480
0443
0462
0488
0486
048A
04AD
04BC
048E
0453
045C
04AA
04EE
04EF
04BF
0484
0444
0407
03FE
044F
04C6
0504
04FE
0508
054C
056D
0503
045F
0460
0541
05D2
046D
00C8
FC9C
FA23
FA0B
FB18
FBB2
FB6E
FAFA
FAF4
FB39
FB66
FB6E
FB88
FBAD
FB9D
FB51
FB1A
FB2D
FB56
FB51
FB36
FB4E
FB8E
FB98
FB50
FB18
FB4B
FBAB
FBB1
FB55
FB1C
FB4E
FB7F
FB37
FABC
FABC
FB38
FB5F
FADA
FABD
FC93
0060
042F
05F1
058C
04A3
048D
050C
0526
04AA
0450
0494
050C
0515
04BA
0486
04A7
04C5
04A1
047E
04A8
04E6
04C9
0462
043A
0485
04CD
04A8
0463
048E
0513
053C
04BB
0433
0453
04D5
04E1
0466
0447
04E7
0514
032B
FF38
FB5D
F9B3
FA3F
FB44
FB67
FADB
FA92
FAD7
FB35
FB52
FB59
FB76
FB79
FB31
FAD9
FADF
FB47
FBA2
FB9D
FB63
FB44
FB48
FB44
FB3D
FB66
FBB6
FBD7
FB9A
FB46
FB3B
FB62
FB57
FB0F
FB02
FB6E
FBC9
FB66
FAB2
FB36
FDF4
01F9
0509
05D0
050F
047B
04D2
0571
058C
0539
0507
0517
0504
04AA
0464
047F
04CB
04F6
0510
054E
0585
0548
049B
041A
0438
049D
04A8
0455
0431
0474
04A8
047A
045E
04E5
05B1
05BA
04CE
0418
0499
057A
04A8
0147
FCFE
FA5A
FA29
FB04
FB45
FAC8
FA7C
FAD4
FB47
FB4A
FB12
FB1B
FB51
FB39
FAC2
FA6F
FA9C
FB02
FB36
FB4B
FB90
FBDE
FBAD
FB00
FAA3
FB2C
FC0A
FC23
FB4D
FA96
FAD6
FB91
FBB5
FB27
FADE
FB4F
FBAD
FB37
FAC8
FC34
FFF1
041D
064E
060B
04EB
048B
04F9
0557
0541
0514
050D
04ED
0491
045E
04B6
054F
057C
0514
04A6
04B7
0513
052F
04ED
04A9
0494
047E
044A
0443
04A8
051B
0502
0467
040F
0472
0501
04E6
0446
0424
04CB
04E4
02D2
FED4
FB2B
F9D2
FA84
FB5D
FB27
FA6B
FA45
FAD9
FB5E
FB55
FB10
FB03
FB17
FB08
FAEF
FB16
FB63
FB66
FB0D
FAD2
FB11
FB7F
FB94
FB54
FB3C
FB74
FB8E
FB42
FAF7
FB37
FBC6
FBE2
FB5F
FB02
FB60
FBDF
FB83
FAA6
FB13
FE03
025B
058D
0637
055A
04D1
0532
05A2
056E
04F8
04EF
053A
0539
04D5
04A1
04F0
0548
051B
04A0
0484
04EA
053B
050C
04AD
0499
04B4
0490
043E
044B
04D9
0545
04FF
046B
045A
04D6
0510
04AA
045B
04CF
053E
03F9
008B
FC9D
FA57
FA2B
FABB
FAC4
FA69
FA76
FAFA
FB47
FB0F
FAD1
FAF9
FB32
FAF5
FA6F
FA5A
FAE6
FB6E
FB5C
FAFC
FB01
FB78
FBBD
FB71
FAFF
FAF5
FB36
FB3C
FAE9
FAAD
FAC6
FAE7
FADB
FAF7
FB89
FC0D
FBA8
FA96
FA79
FCB8
00AC
0419
0575
0541
0501
0556
05B5
0597
0542
052E
0536
04EF
0476
045F
04D3
0537
050B
04AA
04C6
0560
05BF
0574
04EE
04CB
04F5
04DB
0462
041D
047B
0524
0572
0547
050A
04F1
04CC
0485
046D
04B4
04F6
04BB
044A
0466
0509
04E5
02B2
FEDD
FB58
F9BC
F9E3
FA89
FAE3
FB12
FB51
FB5F
FAF3
FA67
FA53
FABC
FB0E
FAF4
FAC7
FAFA
FB65
FB7D
FB22
FAC7
FACB
FAF8
FAF0
FAC0
FAC7
FB18
FB5A
FB51
FB2F
FB3D
FB69
FB71
FB4D
FB34
FB37
FB2B
FB16
FB4B
FBD2
FC0B
FB6D
FA9D
FB3C
FE29
0244
054A
0608
054B
04A8
04BE
050E
051A
050E
0541
058D
0585
0528
04E3
04F4
0518
0502
04CD
04CC
0507
0533
0524
04F5
04CA
049C
046C
046F
04C8
0539
0557
0517
04D5
04C7
04B4
046B
043A
0484
0507
0505
045A
03E7
046D
0534
0474
015E
FD4B
FA7E
F9E6
FA8B
FB07
FAFF
FAEF
FB10
FB0A
FAAE
FA68
FAA3
FB2D
FB74
FB48
FAFC
FADC
FAD4
FAC2
FAC0
FAEB
FB13
FAF7
FAB7
FAB9
FB0C
FB41
FB0D
FAC7
FAEE
FB68
FB9C
FB54
FB0B
FB34
FB88
FB7E
FB36
FB52
FBD9
FBF3
FB2A
FA99
FC05
FFB1
03B5
05D8
05C4
04FB
04D2
052B
0534
04CA
0485
04B6
0502
050D
0506
053B
0580
056B
0504
04CA
04F5
0525
04FB
04B3
04C5
0520
053E
04E6
0485
0487
04C0
04C0
0489
047F
04B0
04A9
043F
03F8
044E
04DD
04DE
0463
0466
0538
0580
0381
FF62
FB78
F9EC
FA9A
FB9B
FB9B
FAFA
FAAF
FADC
FAF2
FABA
FA9B
FACC
FAF5
FAC6
FA90
FAC5
FB38
FB47
FACF
FA6D
FAA8
FB3B
FB7D
FB45
FB01
FAFD
FB09
FAF4
FAF6
FB48
FBA1
FB90
FB38
FB2A
FB8A
FBBF
FB57
FACC
FAE2
FB6B
FB6C
FABF
FAD4
FD28
0137
04AF
05D7
0543
04C2
0524
05AA
057E
04EE
04CB
0531
0582
056B
0547
0567
0582
052D
049B
0463
04A7
04E9
04CD
0498
04B4
04FE
0506
04C1
049B
04C6
04EF
04CD
04A3
04D5
0533
052B
04A9
0445
0460
0491
045B
0422
04A2
0575
04E6
01D1
FD5F
FA2F
F9A7
FAB6
FB66
FB17
FAAC
FADD
FB3E
FB1E
FA9F
FA7F
FAEF
FB5A
FB49
FB01
FB03
FB48
FB66
FB45
FB32
FB4F
FB54
FB0F
FAC8
FADD
FB30
FB53
FB35
FB36
FB7C
FBA8
FB68
FB0D
FB20
FB87
FBA3
FB3F
FAF5
FB3A
FB8B
FB28
FA90
FB70
FEAA
02E4
05AE
0602
0518
04A6
0501
0545
04F4
049C
04DA
055F
056C
04E3
0465
046B
04BE
04EE
04EB
04E9
04EE
04CE
0493
0489
04C7
0503
04FF
04E0
04E1
04DF
0494
0423
0415
0492
0512
0509
04AD
04A0
04F9
0520
04D4
04B7
055B
05F5
04D2
0157
FD0C
FA3D
F9BF
FA75
FAEC
FADF
FAE5
FB32
FB55
FB03
FA9F
FAAD
FB18
FB5C
FB3D
FAFD
FAE1
FADE
FAD1
FAD3
FB05
FB40
FB40
FB05
FAD9
FAE3
FB01
FB18
FB4C
FBAD
FBE8
FBA0
FB00
FAA7
FAD1
FB06
FAD1
FA80
FAB3
FB4B
FB67
FABC
FA81
FC4D
001E
03FC
05E0
05A0
04B5
0467
04B7
0501
0510
052A
0566
0579
053E
0501
050F
0546
054F
051D
04F5
04F8
0503
04F7
04EE
04FB
04F8
04BE
047D
0489
04D9
0510
0500
04F2
051C
0533
04D7
044F
044E
04E9
0546
04BE
03F5
0428
0548
0581
0325
FED4
FB12
F9C2
FA73
FB5D
FB77
FB20
FB08
FB25
FB0C
FAB8
FA8A
FAA8
FAD3
FAE2
FAF9
FB36
FB5C
FB32
FAE4
FAD3
FB03
FB18
FAED
FAD0
FB05
FB4E
FB47
FB01
FAEC
FB1D
FB2F
FAF3
FADC
FB58
FC00
FC02
FB5B
FB0A
FBA3
FC4A
FBC9
FA86
FA96
FD6B
01E3
0547
061A
054F
04BB
04F8
054B
0524
04D8
04E4
0521
0513
04BD
0490
04B5
04D3
04B1
0499
04E0
0550
056D
052A
04F0
04F5
04FB
04CE
04B1
04F4
0555
0545
04BB
0456
047B
04C1
0498
0432
0435
04A6
04C8
0449
03FE
04B9
05B2
04EB
0184
FD1D
FA4E
F9FE
FAD6
FB35
FAF7
FAF6
FB6B
FBA3
FB2D
FA9E
FABE
FB6A
FBCF
FB8E
FB1F
FB05
FB24
FB17
FADB
FABF
FAD6
FAE0
FAC3
FAC5
FB0D
FB52
FB40
FB08
FB19
FB72
FB98
FB57
FB1E
FB55
FBB0
FB96
FB1D
FB00
FB75
FBB5
FB25
FAA5
FBEB
FF62
034D
057E
0593
0502
0512
0579
054B
048B
0426
0499
0544
0558
04E4
049A
04BD
04E0
04AA
0463
0483
04FE
0562
0571
0552
052B
04EE
049F
047A
04A5
04DC
04CE
0495
0495
04D9
04EF
049A
0449
047A
04ED
04F4
0488
047C
0535
059D
040E
005D
FC61
FA2A
F9FF
FA86
FA9E
FA6E
FA9A
FB15
FB42
FAF7
FAC4
FB13
FB8A
FB92
FB2D
FAE7
FB01
FB2B
FB0F
FAD1
FACE
FB08
FB35
FB36
FB38
FB59
FB71
FB61
FB51
FB6D
FB8F
FB75
FB3A
FB39
FB79
FB85
FB18
FAA9
FAD2
FB55
FB50
FA9F
FA8E
FC95
0072
0419
05BE
0580
04E3
04EE
0559
0572
0536
051D
0544
0550
0517
04E5
04FD
0523
04F5
0490
046E
04BB
0511
0506
04B7
0487
048E
0495
0482
0484
04B6
04E5
04DE
04BA
04AE
04AA
047F
0454
048F
0523
0561
04DA
042A
0454
0538
053D
02F8
FF02
FB99
FA5F
FAE2
FB80
FB5F
FAF5
FAF0
FB35
FB3B
FAED
FAB5
FAD3
FB07
FB0E
FB00
FB15
FB37
FB29
FAF5
FAE6
FB0E
FB22
FAF0
FABC
FAE6
FB5A
FBA6
FB8E
FB50
FB3A
FB43
FB49
FB5E
FB9D
FBC6
FB78
FAE0
FAB7
FB4C
FBDD
FB7E
FA99
FAF5
FDC4
0200
0537
05FC
0519
0455
0476
04E6
04F4
04C2
04D1
0523
0544
0500
04AB
049E
04D2
050B
0534
0550
054A
050B
04C3
04C8
051F
055F
0538
04DD
04B2
04C0
04B7
047E
0463
049B
04E1
04DD
04B2
04C9
0512
0502
0474
042B
04D1
05A2
04CC
0178
FD16
FA27
F9CA
FADD
FB8E
FB4B
FAD0
FACA
FB09
FB11
FAE7
FAEF
FB3C
FB76
FB5F
FB28
FB1B
FB32
FB39
FB1F
FAFB
FACF
FA95
FA71
FA9F
FB0F
FB5B
FB42
FB09
FB1D
FB72
FB92
FB53
FB1F
FB52
FB9C
FB76
FB00
FAEC
FB70
FBCC
FB5C
FAE2
FC08
FF63
0368
05DB
0607
052B
04C5
0504
0525
04D4
0497
04E0
055C
0563
04DE
0451
042C
045B
049A
04CF
04FE
0513
04F9
04D2
04D4
04F9
0504
04E5
04D4
04EE
04F6
04AE
044D
0446
04A1
04E7
04CF
04AF
04EC
053F
0503
0449
03FB
048F
04EE
0366
FFBC
FBD1
F9D1
FA0D
FB01
FB43
FAE3
FABA
FB05
FB31
FAE5
FA87
FAA0
FB12
FB51
FB2C
FAFF
FB1E
FB66
FB86
FB72
FB57
FB42
FB1A
FAE8
FADE
FB09
FB35
FB39
FB3A
FB62
FB8D
FB72
FB1D
FAF2
FB1F
FB5B
FB5C
FB53
FB89
FBB7
FB48
FA7A
FAC0
FD5A
01A1
0541
0676
05B4
04DA
04F6
0577
0564
04CC
0481
04DA
0542
0524
04B7
0499
04E8
0531
0521
04ED
04E6
04FE
04F1
04BB
049D
04B8
04E3
04ED
04E1
04D9
04D2
04BD
04B5
04D8
04FF
04E5
0492
046C
04A9
04F8
04E6
0492
047D
04C3
04D6
0461
03F5
0457
051C
049E
01C4
FD90
FA5C
F98C
FA5E
FB1F
FB19
FADA
FAFB
FB40
FB24
FABB
FA91
FAD7
FB21
FB0C
FAC5
FAB0
FAD3
FADE
FAB8
FA9F
FAC5
FB04
FB18
FAFF
FAE5
FADB
FAD3
FAD0
FAF0
FB20
FB19
FACE
FA9D
FADF
FB5E
FB8F
FB49
FB00
FB1A
FB5B
FB52
FB18
FB3B
FBC1
FBE7
FB39
FAAD
FBF0
FF6F
037E
05D7
05D5
04C7
0443
0497
050D
052C
0531
055C
0574
052F
04C4
04B6
0520
0588
0584
0530
04EF
04E0
04DB
04D0
04DC
050E
053E
054D
054D
0558
0554
051D
04CD
04A5
04B1
04AE
0480
0467
04A0
04EA
04D0
045E
0426
0476
04D2
04A5
0436
046E
0563
05B1
03CB
FFE4
FC0A
FA29
FA47
FAEC
FAFA
FAA4
FA9A
FAED
FB15
FADA
FAA0
FABF
FB00
FAF4
FA9D
FA65
FA87
FAC5
FAD4
FAC2
FAC9
FAEC
FAF8
FAE3
FADD
FB07
FB41
FB5B
FB55
FB45
FB28
FAFB
FAF6
FB4E
FBCB
FBE0
FB5E
FAD2
FAD8
FB48
FB6C
FB11
FADE
FB50
FBD0
FB72
FA8A
FADB
FDA4
01E7
052D
05FE
052D
048A
04E0
0589
05B5
0571
054A
055B
0546
04DB
0474
0476
04CF
051B
0524
050E
0509
0511
0506
04DF
04B9
04AD
04BA
04CB
04C9
04A9
0478
045F
0480
04C0
04D4
049B
045B
0475
04E6
0538
0517
04C3
04B2
04D9
04AB
0406
03A9
0450
0555
04E2
01EA
FD9F
FA81
F9DB
FAB0
FB2C
FAB5
FA2B
FA56
FAE2
FB0E
FACC
FABA
FB21
FB91
FB8E
FB2C
FADD
FAD7
FAF1
FAFD
FB04
FB12
FB17
FB0A
FB0B
FB29
FB46
FB42
FB33
FB3C
FB47
FB27
FAF0
FAEF
FB34
FB66
FB40
FB01
FB20
FB96
FBC9
FB65
FAEE
FB16
FBB9
FBF0
FB5C
FB01
FC5F
FFB4
0375
05AB
05CA
04F8
04A5
051D
059D
0583
0507
04CE
0504
053D
0514
04AB
0475
04A0
04EA
0509
04F8
04D9
04BE
04A9
04AB
04D2
050A
0527
0518
04F2
04CF
04B4
04A1
049C
049C
048A
046C
047F
04E4
0548
0529
0497
043B
047C
04DD
04B0
0424
0426
04DE
04F4
02E2
FEF7
FB5D
F9EB
FA5D
FB0D
FAFA
FA90
FA98
FB13
FB6C
FB5E
FB30
FB21
FB1C
FB06
FB09
FB4B
FB97
FB97
FB4F
FB16
FB18
FB25
FB0E
FAED
FAF7
FB29
FB52
FB59
FB59
FB59
FB3A
FAF3
FAC8
FB00
FB76
FBB1
FB7F
FB40
FB61
FBC4
FBDB
FB76
FB10
FB29
FB80
FB67
FAF8
FB79
FE09
01FD
0521
05EE
0508
0453
04B8
0565
0540
0475
0412
047A
04FB
04EE
04A4
04BF
052B
0544
04E1
0494
04CF
0539
0537
04C8
0478
048C
04B8
04B2
04A3
04C5
04EB
04C7
047B
0465
0485
047C
042A
03FB
0446
04BB
04C4
045D
0414
0434
0466
045D
047B
051D
0592
0461
010A
FD05
FA8F
FA81
FB9B
FC15
FB75
FAAA
FA95
FB01
FB25
FAC4
FA62
FA83
FB00
FB51
FB3E
FB13
FB23
FB5A
FB6D
FB4D
FB37
FB56
FB90
FBB1
FBAD
FB9C
FB87
FB6C
FB54
FB4B
FB43
FB25
FAFF
FB09
FB58
FBB0
FBC6
FB9F
FB79
FB66
FB4B
FB34
FB5A
FB9E
FB75
FABC
FA7A
FC20
FFCD
03AC
059A
054E
0473
0491
0577
05EF
057A
04C6
0490
04C4
04DD
04B4
048F
0498
04AE
04B7
04C8
04E1
04C7
0466
0414
0432
04A5
04F9
0504
0508
0530
053F
04F2
0478
0444
046B
048D
046C
044A
0472
04B9
04BC
0482
047D
04CE
04FE
04AE
044F
049C
054F
04EF
0251
FE33
FAD7
F9D8
FAAD
FB7D
FB37
FA6F
FA3D
FACF
FB67
FB6F
FB1D
FAF1
FB07
FB21
FB34
FB69
FBB0
FBB3
FB53
FAF2
FAF9
FB47
FB67
FB3B
FB1B
FB4A
FB8B
FB83
FB40
FB14
FB0B
FAE5
FA9C
FA92
FAF5
FB5D
FB53
FB00
FAF3
FB4E
FB9B
FB97
FBA2
FC09
FC43
FB9C
FA9E
FB19
FE20
0270
0574
05E7
04E3
044D
04BF
055C
0558
04F0
04D0
0511
0542
0528
04F7
04DC
04BA
0476
0448
0477
04E9
053A
0535
0507
04EB
04E7
04E5
04F2
0526
0560
0564
0532
050E
051C
0525
04E6
0480
0456
0481
04A8
0485
0454
046F
04B4
04A7
0441
0428
04B7
0510
03B4
0052
FC83
FA61
FA74
FB5F
FB9D
FB09
FA8F
FABB
FB26
FB36
FAF2
FAC2
FAC3
FABC
FA9E
FAA5
FAEF
FB3A
FB42
FB1E
FB0C
FB07
FAD4
FA78
FA51
FA94
FAFC
FB2B
FB27
FB36
FB55
FB38
FAD7
FAA1
FAED
FB72
FBA1
FB6B
FB48
FB73
FB95
FB61
FB2E
FB70
FBD6
FB95
FAB7
FAA5
FCC0
009E
0427
05A4
0556
04C2
04DD
054B
055B
0506
04CA
04E3
0518
0531
0544
0564
0563
051D
04C9
04C6
0519
0569
0576
0562
0563
056A
0540
04EC
04B6
04C2
04E5
04E9
04DE
04EE
0509
04F1
049F
045C
045A
0475
0473
046F
04A4
04ED
04D2
0445
03FF
04A2
0590
0524
026A
FE67
FB4D
FA5A
FADD
FB58
FB2F
FAE2
FAF5
FB2F
FB13
FAAE
FA76
FA94
FAB3
FA9E
FA94
FADA
FB40
FB56
FB0E
FACB
FAD1
FAF6
FAF9
FAEA
FB00
FB2C
FB21
FAD9
FAAA
FAD0
FB19
FB3C
FB45
FB6A
FB9A
FB90
FB52
FB3E
FB74
FB88
FB23
FAB0
FAE6
FBA8
FBEB
FB23
FA64
FB77
FEC5
02A4
0500
055B
04E5
04D8
053D
0562
0509
04A9
04B4
0508
053D
0531
0518
051D
0531
0533
0521
051A
0529
053A
0534
051A
04FF
04F1
04EC
04E7
04DC
04CB
04BB
04B4
04B8
04C3
04D1
04E2
04F5
04FC
04E1
04A7
0484
04B3
051B
053F
04CD
0434
0446
0510
0554
0398
FFDF
FC07
FA13
FA49
FB36
FB7D
FB1B
FADD
FB13
FB48
FB17
FABA
FAA5
FAEA
FB40
FB6C
FB6B
FB41
FAED
FA94
FA79
FAAC
FAF0
FB18
FB39
FB6D
FB87
FB57
FB0F
FB09
FB43
FB54
FB07
FAB4
FAC5
FB18
FB38
FB21
FB4A
FBD4
FC23
FBAD
FAE8
FACD
FB80
FBFD
FB69
FA65
FAA7
FD2A
010E
0459
05BE
0583
04DC
04B3
0511
0572
0574
052E
04F2
04E2
04DB
04BF
04A3
04A6
04C4
04DD
04E2
04D9
04C4
04A7
0496
04A8
04D3
04E5
04C5
04A1
04AD
04D4
04DE
04D8
0502
0550
0558
04F3
0495
04B6
051D
0525
04B3
0460
048D
04C5
0483
0430
049F
0575
04F5
01FC
FDB5
FAA6
FA14
FAF6
FB81
FB22
FA96
FA96
FAF9
FB3E
FB48
FB4A
FB4D
FB2F
FAFC
FAE8
FAFE
FB16
FB14
FB04
FAF2
FADC
FACC
FADD
FB14
FB57
FB88
FBA6
FBBC
FBBE
FB95
FB47
FAFF
FADA
FAD4
FAED
FB25
FB57
FB4B
FB11
FB02
FB45
FB8D
FB8D
FB68
FB6D
FB85
FB57
FAF9
FB03
FBA2
FC04
FB64
FA86
FB50
FE8D
02A3
052E
0578
04CF
0498
04E3
04F9
04B2
0493
04DD
0530
052F
050D
0526
0568
057C
054E
0515
04F1
04D8
04CC
04DD
04EE
04D3
0497
0481
04B5
04FD
0511
04F7
04EB
04FF
0505
04ED
04DE
04EA
04E8
04C9
04C9
0503
0533
0517
04D5
04BC
04C5
04B5
049B
04C1
0512
0506
0479
042A
04BB
0559
0434
00BD
FCB2
FA5E
FA38
FADB
FB07
FAD8
FAF6
FB5E
FB83
FB3B
FAF8
FB04
FB16
FAE0
FA95
FA95
FADD
FB28
FB5D
FB81
FB77
FB28
FAD4
FACF
FB0D
FB33
FB1E
FB14
FB4C
FB8D
FB87
FB50
FB48
FB74
FB7B
FB40
FB21
FB53
FB7E
FB4F
FB03
FB02
FB35
FB3D
FB1C
FB2D
FB77
FB93
FB5B
FB44
FB9E
FBD4
FB44
FAB0
FBE2
FF71
0391
05DB
05CD
04E9
0494
04C6
04CD
0497
049E
0501
054E
0540
0528
0558
05A1
05AD
0583
055D
0539
04FD
04C3
04B5
04B9
04A3
048E
04B4
0505
052F
0513
04F9
0513
0520
04D1
045F
0453
04B1
04F1
04D4
04C2
04FB
0516
04B0
0429
0423
0484
04A8
0471
046F
04DD
051E
04BD
0463
04EE
05A4
0484
00D5
FC80
FA19
FA14
FACB
FADD
FA82
FA8A
FAF2
FB20
FAEF
FAD3
FB04
FB24
FAF5
FAC9
FAF6
FB3C
FB3C
FB14
FB1C
FB43
FB38
FAFC
FAE0
FAFC
FB13
FB04
FAF7
FB0D
FB1C
FAF7
FAD2
FAFC
FB60
FB99
FB91
FB97
FBB6
FB8B
FAFD
FA99
FAC8
FB2B
FB39
FB1A
FB4D
FBB4
FBAA
FB1F
FAE2
FB67
FBDE
FB66
FAD3
FC2F
0003
0433
0641
05FF
0538
0530
057E
0555
04D1
0495
04BF
04E0
04D4
04E6
052B
0548
0517
04FD
053C
0570
0532
04C7
04B6
04ED
04F2
04B8
04A9
04EC
0521
04F6
04AB
04A7
04D4
04C9
0487
047D
04C7
04F6
04D0
04B6
04F5
0534
050B
04B7
04AB
04C6
0495
0431
042C
0499
04CD
0475
044D
04F9
0573
03CC
FFC3
FBA3
F9D1
FA41
FB0B
FB03
FAB1
FAE1
FB5E
FB76
FB14
FABC
FAA6
FA8C
FA54
FA53
FAA8
FAEF
FAE0
FACB
FB02
FB48
FB3B
FB07
FB18
FB5D
FB67
FB2A
FB13
FB57
FB97
FB76
FB30
FB38
FB76
FB64
FAFA
FACD
FB21
FB76
FB60
FB39
FB77
FBD5
FBC7
FB64
FB3D
FB6D
FB81
FB53
FB5D
FBC9
FBE6
FB3E
FAEC
FCBD
00BA
0495
061F
059F
04F0
050A
0552
0522
04D0
04F4
0563
0584
054B
052E
054C
053C
04D8
04A0
04EC
0559
0566
053A
053B
0551
051E
04BA
0496
04C7
04E6
04BE
049F
04CE
0501
04C6
044D
0430
0486
04C0
04A2
04A0
0505
054C
04E8
0431
03E4
0413
0433
0415
041F
0479
04B1
0489
048B
051B
053C
0355
FF6B
FBAB
FA1C
FA80
FB13
FAE3
FA76
FA74
FAAF
FAB9
FAA8
FAD2
FB20
FB29
FAEE
FADD
FB17
FB31
FAF3
FAC0
FAEF
FB38
FB37
FB14
FB2E
FB66
FB5D
FB22
FB26
FB7A
FBA5
FB5B
FAFB
FB00
FB42
FB3D
FAFF
FB15
FB8F
FBC8
FB6B
FB11
FB50
FBC8
FBC9
FB71
FB6A
FBC9
FBF1
FBA5
FB76
FBBA
FBD2
FB36
FAEE
FCC5
00CC
04AB
061A
055E
0482
04AC
053C
054A
04FB
04F3
053B
0554
0515
04EA
0513
0545
0536
0515
0527
0545
052E
0501
04FB
050D
0500
04E5
04E7
04EB
04B5
045F
0447
0489
04C7
04B8
0495
04BB
0501
04F0
0491
0470
04B5
04DB
0490
044B
047C
04C7
049D
0437
043E
04A5
04AF
043C
0437
0510
0557
031B
FEA3
FAB5
F996
FA9D
FB84
FB52
FAEE
FB2F
FB9E
FB6C
FAC3
FA6E
FA9F
FAC3
FA86
FA4E
FA7C
FACA
FAC7
FA93
FA95
FAD0
FAF5
FAF5
FB05
FB34
FB58
FB64
FB74
FB80
FB57
FAF4
FAAE
FAD0
FB33
FB7B
FB9B
FBCF
FC0C
FBFA
FB91
FB4B
FB6B
FB99
FB7B
FB4A
FB57
FB6F
FB3A
FAFB
FB45
FBE5
FBE0
FB02
FADA
FD2A
0174
050F
060D
0537
049F
04FF
0569
051F
04A3
04B5
0533
0572
0552
0550
05A4
05E7
05BD
0564
0540
0543
052B
0506
050E
0530
0528
04F4
04CA
04B8
049F
0484
0497
04DC
0512
0502
04D3
04C3
04BF
0487
0439
043C
0499
04D8
04B7
0490
04AD
04CA
0496
045B
048B
04EA
04D0
044C
0442
04EA
04D9
0272
FE39
FAC4
F9EC
FAD7
FB66
FADA
FA39
FA62
FAE4
FAE6
FA71
FA3D
FA8A
FAD9
FAC0
FA82
FA8A
FAC7
FAE2
FACF
FAC4
FACF
FAD2
FAD0
FAE8
FB13
FB2B
FB25
FB11
FAF9
FAD7
FAC0
FADB
FB23
FB5F
FB61
FB48
FB49
FB56
FB44
FB2E
FB5B
FBAD
FBAF
FB4E
FB17
FB5D
FBAC
FB7F
FB2D
FB64
FBF4
FBE3
FB17
FB2F
FDD0
0240
05BD
067B
0576
04D8
054D
05C4
056F
04DC
04E1
055B
0584
052D
04F3
053D
05A9
05AA
0553
051D
0531
054D
054D
054D
0562
0571
0561
053E
051C
050E
051D
0540
0555
0537
04EB
04A1
0480
047C
0479
0480
04A1
04BF
04A8
047D
048E
04CD
04D1
0486
046A
04C7
0519
04C3
0421
042B
04D3
0483
01DF
FDC4
FAB5
FA22
FB01
FB6E
FAF0
FA79
FAA4
FAF2
FAC8
FA62
FA5A
FAB2
FADC
FAA2
FA6D
FA96
FAE1
FAE6
FAB7
FAAB
FAD0
FADF
FAB9
FA95
FAAC
FAF6
FB45
FB75
FB7E
FB6E
FB5F
FB67
FB7D
FB7D
FB55
FB25
FB1C
FB38
FB53
FB63
FB79
FB80
FB4D
FAF7
FADB
FB16
FB4C
FB3A
FB21
FB54
FB87
FB2F
FAA8
FB65
FE62
029C
05B9
0662
057C
04CC
04FA
055E
0552
0507
04F6
0523
0541
0534
0529
0535
053A
052B
052B
0549
054F
0514
04C3
04A5
04C1
04E0
04E0
04C6
049D
0472
045D
0472
04A0
04C5
04DC
04FF
052D
0534
04F8
04AC
0493
04A0
048E
045E
0459
0494
04BF
04AA
0496
04BF
04DF
049C
0441
0470
04E3
042C
0143
FD2F
FA5B
FA16
FB45
FBEB
FB6A
FABD
FACA
FB44
FB65
FB0F
FACF
FAF5
FB37
FB34
FAFE
FAE5
FAF8
FB07
FB00
FB09
FB38
FB6C
FB7D
FB6D
FB60
FB6D
FB83
FB82
FB5F
FB3B
FB3F
FB65
FB7E
FB73
FB61
FB6D
FB88
FB82
FB54
FB31
FB3D
FB59
FB5A
FB5B
FB87
FBB3
FB8E
FB40
FB59
FBDD
FBF5
FB0D
FA23
FB22
FEA7
02EC
0577
05A2
04EB
04D9
0552
0563
04ED
04B4
051B
0591
0579
0505
04D4
0504
0521
04EF
04BE
04DD
051B
051E
04EB
04D0
04DA
04D1
04A2
0479
0478
0482
0475
0466
0477
0499
04A3
04A0
04C0
0505
051E
04DC
0481
0472
04A5
04AE
0469
044D
04DD
05C3
05BC
03AD
FFE3
FC1E
FA21
FA37
FB21
FB82
FB18
FA9E
FAA5
FAF8
FB1B
FB01
FB04
FB3E
FB5E
FB2F
FAED
FAE7
FB0D
FB1B
FB04
FAF8
FB09
FB11
FB04
FB06
FB2D
FB4D
FB3D
FB23
FB42
FB83
FB8D
FB51
FB2C
FB46
FB4A
FAF3
FA9C
FAC7
FB45
FB6A
FB11
FAF4
FB8F
FC2C
FBBE
FA9A
FA98
FD09
0101
0443
0588
056E
0535
0549
054E
0510
04DA
04E5
0501
04F0
04CF
04D7
04F0
04D8
049A
048D
04D1
051C
051E
04F0
04E1
0509
052C
0521
050B
0520
0549
053B
04EA
04A9
04C2
0515
054B
054B
0549
055B
0543
04CE
0442
0422
0477
04B6
048E
0483
052B
05F1
0538
022C
FE10
FB2B
FA81
FB0F
FB53
FB0A
FAFB
FB76
FBD9
FB9C
FB23
FB0E
FB49
FB4D
FB14
FB26
FBAD
FC10
FBC5
FB24
FAE7
FB24
FB41
FAEC
FA9C
FAC5
FB1B
FB0D
FAAE
FA92
FAE6
FB26
FAF5
FAAA
FACD
FB3A
FB5E
FB1B
FAF6
FB3A
FB80
FB5B
FB22
FB72
FC09
FBEB
FADD
FA42
FBCE
FF82
0363
056B
056F
04D0
04B0
04F0
04EE
049B
0475
04AD
04DE
04B3
046B
0471
04B4
04BC
0463
0419
0449
04C1
04F8
04D6
04C6
0503
0541
052A
04ED
04FC
0552
0576
052E
04DA
04E0
0519
0517
04E2
04E6
0530
0544
04E3
0482
0496
04C9
047E
03F9
0436
0547
058B
034C
FF00
FB33
F9DD
FA7F
FB38
FB24
FAEE
FB42
FBBA
FB99
FB09
FADA
FB4C
FBB6
FB8C
FB22
FB1F
FB7D
FBA8
FB65
FB1C
FB2A
FB56
FB3D
FAF4
FAE3
FB20
FB4B
FB23
FAE7
FAF4
FB32
FB3D
FB02
FAD7
FAF0
FB12
FAFE
FAE9
FB33
FBC0
FBFF
FBB7
FB66
FB84
FBB3
FB42
FA80
FAFA
FDD3
021A
0565
063A
0569
04CE
0521
0599
0566
04E0
04D4
0547
057B
051A
04B2
04D5
0544
055A
0500
04BA
04D0
04F4
04CD
048C
0492
04D9
0502
04F2
04EF
051D
0534
04F7
04AB
04B9
0505
0511
04BA
046D
0482
04BD
04B8
0492
04B7
0517
0516
048F
0448
04EC
05AF
04CB
0182
FD45
FA67
F9DA
FA8F
FB05
FAE1
FAC6
FB10
FB55
FB22
FAA4
FA60
FA78
FAA1
FAAC
FAC2
FB05
FB41
FB33
FAF1
FAD4
FAFF
FB3D
FB5B
FB67
FB78
FB6D
FB22
FACB
FAC8
FB1D
FB59
FB29
FAD2
FACB
FB17
FB4A
FB38
FB2F
FB6E
FBA9
FB7B
FB26
FB4D
FBE8
FC12
FB52
FAB7
FBF9
FF6A
0347
056E
0578
04C6
04A7
0516
0554
0530
051C
0554
057D
0544
04E5
04CD
04F9
050D
04F1
04EE
052F
0566
053D
04DC
04B7
04F2
0538
0548
0545
0565
0581
0549
04D0
0486
04A1
04D0
04B6
0474
0471
04B2
04C8
047F
0438
045A
04A6
0499
044D
0478
052B
0528
030D
FF24
FB7C
F9EE
FA57
FB1F
FB32
FAE1
FAEB
FB4A
FB68
FB1D
FADC
FAF2
FB1E
FB0B
FAE3
FAFC
FB43
FB4E
FB03
FACC
FAFA
FB45
FB3C
FAE7
FAB2
FACA
FAE4
FAC2
FA94
FAA7
FAE9
FB0D
FB0A
FB28
FB88
FBD9
FBCB
FB88
FB74
FB97
FBA1
FB7A
FB7B
FBD1
FC04
FB89
FAD5
FB56
FDF9
01DC
04EA
05D3
0531
0498
04D1
0561
0586
0540
050E
051F
0527
04F2
04C0
04D5
050B
050E
04E7
04EB
052E
0558
0530
04F8
0508
053E
0529
04B5
0456
0469
04BB
04DB
04BF
04B6
04DA
04EA
04C4
04AB
04CF
04F1
04C8
0488
049B
04EB
04E7
046F
043C
04DB
0578
0464
010F
FD05
FA7E
FA33
FAFC
FB69
FB33
FAF5
FB08
FB26
FB05
FACC
FAC1
FAD7
FAD7
FAC8
FAE2
FB22
FB40
FB1B
FAF0
FB07
FB47
FB5D
FB2D
FAFB
FB0A
FB45
FB60
FB43
FB1C
FB1A
FB31
FB46
FB57
FB6C
FB74
FB5C
FB42
FB5B
FBA0
FBBA
FB75
FB1A
FB19
FB59
FB40
FAB2
FAB5
FC98
004A
03FE
05CC
0587
04AC
0494
052C
058A
054B
04EA
04DB
04F8
04ED
04D1
04E6
0515
0502
04A6
046D
0498
04DF
04DE
04A6
049E
04D9
04FB
04CD
0493
049F
04D4
04DA
04B1
04A8
04D5
04F6
04E0
04C8
04E5
0504
04D2
046E
0454
049A
04BC
0474
0453
0506
0600
0598
02C5
FE88
FB25
F9FF
FA85
FB2A
FB1B
FAB2
FA88
FAAD
FACD
FACA
FAD2
FB05
FB44
FB68
FB73
FB7D
FB7B
FB53
FB17
FAFD
FB1F
FB54
FB69
FB67
FB78
FB98
FB95
FB55
FB0F
FB09
FB42
FB72
FB6A
FB43
FB25
FB11
FB01
FB13
FB5B
FB99
FB7C
FB2D
FB3D
FBC9
FC11
FB63
FA6A
FAF3
FDF7
0235
053D
05E2
052D
04CD
052C
057D
0536
04C8
04CC
0521
053B
04FE
04D1
04E7
04FB
04D8
04BE
04F9
0555
055D
050C
04D2
04EC
0512
04EF
04A8
04A1
04D9
04ED
04AA
0457
044A
0471
0488
048E
04B3
04E2
04C2
044A
03F4
0429
04A9
04DE
04C1
04EE
059D
05D2
0425
007D
FC90
FA64
FA65
FB41
FB85
FB0F
FAB3
FAEB
FB46
FB2D
FABA
FA81
FAB8
FAF9
FAE7
FAAB
FAA5
FAE1
FB18
FB2A
FB3D
FB5F
FB5E
FB12
FAB7
FAA9
FAE3
FB07
FAEA
FAD5
FB0A
FB5D
FB71
FB45
FB29
FB49
FB76
FB82
FB7D
FB82
FB71
FB34
FB12
FB5A
FBB6
FB6A
FA86
FA6F
FC8D
0086
0436
05C2
0552
048C
049D
053D
058D
055C
0522
0529
053A
0512
04CF
04B5
04C8
04E2
04F1
0504
0517
050A
04DE
04C6
04E2
050C
050C
04E5
04D4
04F1
0516
051C
050A
04FF
04FD
04FB
0502
0521
053C
0517
04AE
0461
0486
04ED
050A
04BA
0496
0523
05CA
0514
0231
FE23
FB0A
FA28
FAD8
FB86
FB65
FAE9
FAC6
FAF9
FB10
FAEE
FADA
FAF8
FB07
FADD
FAB9
FAEB
FB4E
FB6F
FB34
FAFC
FB0E
FB33
FB1E
FAE7
FAE2
FB18
FB3D
FB2D
FB1C
FB36
FB4F
FB34
FB14
FB3D
FB86
FB6C
FADB
FA71
FAAD
FB2F
FB49
FB01
FB07
FB88
FBC1
FB25
FAA4
FBEE
FF5C
032A
0531
051B
0468
0475
051A
0567
0510
04B1
04CC
0527
0549
052A
0520
053D
0535
04DC
047A
046C
04B2
04FD
0515
0502
04DC
04AF
0493
04B3
0514
056A
0560
0502
04B0
04A6
04B9
04B0
04AD
04E3
051F
04E1
0427
03A3
03F4
04C3
0520
04D5
04B8
055E
05CE
044C
0086
FC6A
FA4B
FA85
FB70
FB83
FAE1
FA9B
FB08
FB7A
FB5A
FAF3
FAD5
FB03
FB14
FAEF
FADD
FB01
FB22
FB0E
FAF1
FB04
FB2D
FB37
FB34
FB63
FBB2
FBBB
FB5F
FB04
FB04
FB23
FAF8
FAA5
FAB2
FB38
FBA5
FB90
FB5C
FB9A
FBFD
FB9F
FA88
FA47
FC6A
007C
0427
0587
04EC
041D
043D
04DE
050E
04AE
0467
04A7
051C
0544
0510
04D8
04D4
04EE
04FE
04F6
04DE
04B4
0488
047E
04A5
04D7
04E0
04C4
04B6
04CF
04E6
04D9
04C3
04C9
04D0
04A2
0458
0453
04A1
04C7
046E
040F
0472
0556
0523
028A
FE50
FAE6
FA02
FAFD
FBE1
FBAD
FB0B
FAF2
FB52
FB72
FB25
FAF4
FB38
FB93
FB87
FB33
FB10
FB3C
FB6B
FB75
FB80
FB9E
FB95
FB3F
FAE3
FADF
FB24
FB4D
FB3F
FB45
FB87
FBB4
FB82
FB36
FB3C
FB7E
FB7F
FB36
FB34
FBB7
FC05
FB5D
FA64
FAF2
FE08
0254
0554
05D9
04F8
0476
04DC
0561
0552
04ED
04C9
04F3
0504
04CC
0492
0491
04A2
048B
045D
0456
047A
0491
0482
047A
049B
04BF
04AC
0471
0452
0466
0481
0481
0483
04A3
04BB
04A1
047C
049F
04F5
0506
04B2
0492
051D
0598
046F
010B
FCE7
FA52
FA1D
FAFA
FB3B
FAA5
FA35
FA84
FB16
FB42
FB18
FB15
FB4A
FB53
FB17
FAFD
FB3D
FB7C
FB52
FAF6
FAF4
FB5A
FBA4
FB77
FB1D
FB09
FB3D
FB63
FB61
FB68
FB82
FB72
FB2B
FB08
FB3C
FB6F
FB39
FADC
FAF9
FB83
FB9E
FAEA
FA89
FC29
FFE9
03D8
05D1
05A2
04D3
04AE
050D
0520
04C6
0493
04D2
051B
0504
04C3
04D2
052C
0558
051A
04C1
04A6
04B3
049A
045E
044F
0487
04BD
04AB
0472
0465
0495
04CF
04EC
04F4
04E6
04AA
045C
045A
04C7
0524
04DC
042D
040C
04BD
0504
0345
FF8B
FBDD
FA37
FA90
FB39
FB0C
FA7E
FA85
FB10
FB45
FAD0
FA59
FA82
FB0F
FB54
FB36
FB27
FB5D
FB82
FB51
FB18
FB3A
FB8D
FB8D
FB24
FAC4
FACD
FB1B
FB5E
FB8C
FBB6
FBBB
FB73
FB1B
FB26
FB8C
FBAB
FB30
FAA7
FAC1
FB3C
FB37
FAAE
FB05
FD84
0184
04CF
05E2
055D
04F0
054F
05C1
0587
04E7
04A5
04E8
052E
0521
0505
0526
0551
0527
04B7
0473
048F
04C4
04BF
0494
0486
04A5
04C2
04C9
04D0
04D8
04BD
0483
046F
04A7
04E5
04CD
0478
0464
04B1
04E1
049F
046A
04EE
05AC
04FE
01E0
FD81
FA5A
F9C0
FABA
FB6F
FB3D
FAEA
FB1E
FB74
FB44
FAB0
FA67
FA9E
FAD9
FAC5
FAB5
FB0E
FB91
FBA7
FB3D
FAE1
FAF6
FB3B
FB43
FB12
FAF8
FB08
FB12
FB13
FB3B
FB80
FB8B
FB3F
FB0A
FB4D
FBAB
FB7C
FADA
FAAC
FB57
FBF8
FB92
FAC0
FB6B
FE87
02A4
054C
059C
04DE
04AB
0525
0563
0504
04A3
04CA
0527
0527
04DA
04CE
0529
056C
0530
04B3
0473
0484
0497
0486
0482
04AD
04DC
04E3
04DF
04FC
0518
04F5
04AC
049A
04CF
04E0
048C
043C
0478
0509
0527
04A6
0460
04F8
0583
042D
007B
FC42
F9EF
FA12
FB18
FB64
FAED
FAAD
FAF8
FB2F
FAE2
FA83
FAAB
FB30
FB6D
FB37
FB05
FB2A
FB63
FB51
FB0F
FAF7
FB0D
FB0B
FAEE
FB0D
FB7C
FBCA
FB91
FB15
FAE1
FB04
FB16
FAF1
FAF0
FB48
FB89
FB43
FAD9
FB11
FBD1
FC09
FB4B
FAE3
FC9F
007F
0451
05FA
058F
04D4
04F4
0571
055A
04C1
0476
04C6
0525
0518
04DA
04D7
04F8
04D7
0475
044B
0493
04F3
050A
04F6
0505
052B
0516
04CA
04B1
04F5
052E
04EF
0475
045A
04B9
050E
0500
04D7
04EC
04F4
047F
03EA
041B
050B
051E
02C0
FE7C
FAD2
F9AD
FA7D
FB49
FB18
FAB1
FB08
FBCC
FBF6
FB4E
FAA9
FAB3
FB23
FB5B
FB4E
FB5A
FB86
FB6E
FAFB
FA9B
FAA5
FAD9
FAD2
FAB4
FAF7
FB92
FBE9
FB9D
FB1A
FAFA
FB37
FB55
FB38
FB3E
FB8E
FBBE
FB83
FB3E
FB6D
FBB6
FB53
FA88
FAFF
FDF5
025C
058E
05FF
04BD
03F9
0486
0560
0564
04C0
045F
0491
04DB
04DF
04D7
0505
0532
050C
04BC
04B8
0509
0532
04DC
045B
0432
046B
049D
0492
047D
0495
04BF
04CB
04C6
04D3
04D5
049A
0446
043B
047C
048A
042A
03F4
0491
056E
04D8
01D2
FD89
FA71
F9DD
FAE0
FBAD
FB93
FB36
FB3D
FB6E
FB4A
FAE8
FAC6
FAFC
FB15
FACF
FA8C
FAC5
FB54
FBA1
FB6B
FB0E
FAFB
FB36
FB6D
FB72
FB59
FB44
FB41
FB51
FB6B
FB67
FB2B
FAEE
FB16
FBAA
FC1B
FBF2
FB7E
FB79
FBF0
FC09
FB43
FA9C
FBD4
FF55
035E
05AC
05B3
04DC
04A7
051D
0554
04E7
0468
046F
04D0
04FA
04CB
049D
04AC
04C3
049F
0459
0442
0477
04CD
0509
0512
04F1
04C6
04B9
04D5
04E4
04A6
0439
0419
047F
04F0
04C7
041F
03CC
0447
04EA
04C6
0408
03DF
04C5
0568
03EB
0030
FC4B
FA61
FA8F
FB2F
FB00
FA62
FA5F
FB29
FBF1
FC0D
FBA9
FB55
FB43
FB3F
FB24
FB0A
FB05
FB07
FB06
FB15
FB36
FB45
FB35
FB2E
FB52
FB7C
FB76
FB61
FB92
FBFC
FC1B
FBA8
FB28
FB53
FC08
FC56
FBC3
FB08
FB17
FBB3
FBBC
FAF7
FADF
FD0A
0107
047E
059E
04E6
0431
0479
051B
052B
04BB
0487
04D2
0527
0525
04FE
0502
051E
050B
04D5
04C6
04E6
04E6
04A2
0460
0466
0491
048E
045F
044E
046B
0472
044B
0444
0494
04E1
04AF
042B
0408
0475
04BE
0451
03C7
0433
0558
0559
02BA
FE68
FB07
FA38
FB1A
FBB2
FB3F
FAA2
FABE
FB43
FB60
FAFC
FABE
FAF6
FB34
FB03
FA9E
FA95
FAFE
FB68
FB81
FB76
FB8B
FBAC
FB99
FB58
FB34
FB50
FB8E
FBC7
FBEE
FBED
FB9E
FB20
FAE4
FB34
FBAE
FBAF
FB3B
FB0A
FB7B
FBDC
FB58
FA7E
FB21
FE4A
02A7
059D
05EC
04CB
0436
04BF
0561
0538
049C
046D
04D9
0547
0545
050A
04F7
0504
04F5
04C8
04B0
04B6
04AB
0480
0469
048A
04BB
04C8
04B9
04B8
04BD
04A1
0476
0485
04CD
04E1
0481
0416
0437
04C2
04F6
048C
0445
04D4
0579
0471
010C
FCDE
FA4F
FA2A
FB1C
FB7F
FB1F
FADE
FB2B
FB7C
FB46
FACA
FAA5
FAEB
FB2D
FB36
FB4E
FBA7
FBFB
FBE7
FB79
FB16
FAEC
FAD7
FAC4
FAE1
FB42
FB96
FB86
FB35
FB16
FB49
FB7A
FB6B
FB4B
FB60
FB86
FB76
FB50
FB7A
FBE0
FBD1
FB10
FAB2
FC3C
FFCA
0387
056B
053B
047E
0487
0523
0553
04CD
0442
0447
049B
04AA
0465
043A
0463
04A4
04BD
04C5
04F0
0526
0527
04F1
04C2
04C3
04DB
04F0
0510
053F
0545
04F2
0482
0464
049F
04BD
0470
040A
0400
0430
040F
03A5
03B7
04A1
0541
03D4
0015
FC01
FA04
FA95
FBF6
FC57
FB9B
FAEA
FAFC
FB6F
FBA0
FB86
FB76
FB75
FB45
FAEF
FAD1
FB10
FB54
FB43
FAFE
FAE6
FB02
FB06
FADE
FAD6
FB17
FB53
FB3B
FB0B
FB3A
FBB5
FBE3
FB8B
FB46
FBA0
FC1B
FBC7
FAD7
FAFB
FD8E
01C2
052C
062F
0566
0488
046E
04A2
0493
046C
0492
04DB
04D0
0473
0447
0488
04D6
04CB
048E
0487
04B7
04C1
0490
047C
04B1
04D6
0495
043F
046C
050C
0561
04FD
0468
045E
04BD
04BC
043A
041F
0504
05E1
04D1
014D
FD12
FA7F
FA3F
FB00
FB39
FABD
FA5F
FA9F
FB1F
FB58
FB46
FB38
FB4A
FB5E
FB6B
FB88
FBA7
FB98
FB5A
FB3A
FB6A
FBAA
FB97
FB44
FB2F
FB89
FBDF
FBB2
FB2B
FAEF
FB2F
FB6C
FB46
FB27
FBA5
FC67
FC4C
FB09
FA1B
FB7D
FF57
0381
059E
0561
047C
0475
052E
0597
0542
04BC
0496
04AD
049B
0465
0462
04A0
04D0
04C4
04B0
04C4
04DB
04B7
0473
0460
048C
04B0
04AC
04B8
04F0
04FC
0491
040B
041A
04B9
0505
0470
03BC
041A
0551
0572
02E5
FE80
FAE6
F9DB
FAAB
FB64
FB1D
FA8E
FA9F
FB2F
FB7A
FB42
FAFD
FB0A
FB37
FB2F
FB06
FB07
FB32
FB3E
FB12
FAE9
FAF1
FB01
FAF1
FAEE
FB39
FBAA
FBCA
FB7A
FB2D
FB46
FB80
FB59
FAEF
FAF8
FBAA
FC29
FB93
FA83
FADE
FDC5
0206
0525
05D8
0517
04A7
0511
057D
052E
0485
044F
04A0
04DB
04AE
0479
049E
04EA
04F9
04DC
04FD
0560
0581
0513
0483
0476
04E9
0540
0523
04DE
04CC
04C3
047B
0425
042E
047E
0479
0408
0402
04FA
05E3
04C3
0101
FC8D
FA11
FA3D
FB62
FBA8
FAFA
FA83
FAD3
FB4C
FB46
FB01
FB16
FB7A
FB9D
FB4F
FAFF
FB01
FB1E
FB06
FAE2
FB0A
FB5D
FB5B
FAF1
FAA8
FAE2
FB40
FB37
FAF2
FB17
FBB9
FC19
FBB5
FB22
FB42
FBE0
FBE0
FAF5
FA9A
FC8C
008D
044E
05C7
0530
0453
0459
04D9
04EF
048F
0463
04B2
0518
052E
0515
0514
0519
04EA
04A6
04B4
0524
0583
0570
051E
04FB
050C
04F7
04AC
048E
04D0
0509
04BB
0426
0404
047C
04C5
044C
03B5
0427
0576
05BE
035C
FF05
FB4E
FA0D
FAAE
FB4A
FAF3
FA56
FA5B
FAE2
FB31
FB17
FB09
FB47
FB74
FB33
FAC3
FA9D
FAC0
FAC6
FA9B
FA9F
FB06
FB70
FB71
FB33
FB35
FB7B
FB84
FB1F
FAD1
FB10
FB81
FB71
FAF7
FAE9
FB90
FBFC
FB4C
FA49
FAF9
FE3E
0288
0553
05C4
0522
04FA
0562
0577
04E9
0463
047D
04EC
0512
04E1
04C5
04E4
04F2
04C9
04B5
04FA
0555
0553
04F5
04A8
04A4
04B0
049F
04AE
050C
0553
04F3
041C
03C0
0465
055B
058E
04FA
04B4
0540
057A
03AE
FFCE
FBE5
FA1D
FA95
FB8D
FB83
FA9E
FA06
FA47
FAE0
FB26
FB18
FB1D
FB4F
FB6D
FB5B
FB51
FB74
FB8F
FB5E
FB05
FAEC
FB34
FB8B
FB9B
FB6B
FB34
FB04
FAC9
FA9E
FABF
FB1A
FB46
FB14
FAF1
FB54
FBE9
FBD0
FAF4
FAB0
FC97
007C
044C
060D
05C4
0512
0527
05AA
05A4
04F5
045F
0464
04B5
04CB
04AD
04BC
04FD
0512
04D1
0487
0486
04AF
04B0
047F
0463
0486
04CB
0511
0561
05AE
05AD
0536
049F
0462
0473
0452
03E5
03DE
04CB
05DF
0551
023B
FDE1
FAA1
F9B6
FA45
FAB7
FA75
FA26
FA78
FB3A
FBBD
FBB5
FB69
FB2E
FB09
FAE3
FAC8
FAD6
FB02
FB21
FB28
FB2B
FB3A
FB43
FB3B
FB33
FB37
FB32
FB0E
FAF6
FB2B
FB9C
FBD9
FB9D
FB40
FB4E
FBBD
FBCB
FB0F
FA6F
FB8D
FEF9
033A
05FB
063F
052A
0486
04E2
055C
0515
044C
03EC
044E
04ED
0532
0525
0526
054D
0557
052B
0501
050B
0527
0518
04E3
04C0
04BC
04B5
049A
048E
04A2
04B3
04A9
04A5
04B9
049F
0418
038F
03DB
0505
059D
03E8
FFEE
FBDF
FA05
FA8F
FBB1
FBCE
FB04
FA7C
FABD
FB38
FB4A
FB11
FB0A
FB44
FB57
FB12
FABD
FAAB
FAD1
FAEC
FAE6
FAE2
FAFB
FB30
FB75
FBB6
FBC4
FB78
FB0D
FB01
FB79
FBEA
FBC1
FB38
FB2C
FBE0
FC65
FBB8
FA5D
FA4C
FCE2
0129
04A4
05C0
052C
04A6
04F9
0577
0545
048B
0425
0478
0510
054D
0520
04E4
04CE
04C4
04B4
04C1
0503
0547
0545
04FF
04C0
04B9
04CE
04C8
049D
046B
0449
0446
047A
04E0
0520
04D4
042A
03FB
04CC
05C0
050E
01DF
FD8E
FA8F
FA0B
FAF1
FB72
FB07
FA96
FADE
FB76
FB89
FB06
FAA4
FAC9
FB13
FB0E
FAE2
FAFA
FB4A
FB59
FB07
FAC6
FAFD
FB69
FB83
FB35
FAE5
FADA
FAF0
FB01
FB2A
FB77
FB98
FB52
FB04
FB44
FBDE
FBDD
FAE8
FA47
FBC9
FF97
039F
0597
0547
0464
046A
0528
058B
0537
04CD
04E1
053C
0555
0519
04DD
04C9
04B7
0499
04A0
04D9
04FD
04CE
047E
0478
04C8
0508
04F4
04CC
04E4
051A
0500
048E
0440
0464
049B
0463
03F4
0416
04E2
051F
0357
FF9E
FBDF
FA15
FA6B
FB53
FB68
FAC6
FA70
FADF
FB81
FBA6
FB5C
FB29
FB33
FB27
FAE0
FAC1
FB25
FBC4
FBF9
FB96
FB1F
FB1A
FB66
FB7B
FB27
FACA
FAD0
FB34
FBA9
FBF4
FC02
FBCD
FB71
FB3C
FB61
FB97
FB68
FB0C
FBAD
FE44
022A
054B
060F
04EF
03D3
03FA
04ED
057C
053D
04CB
04B9
04DD
04BF
0459
0415
043C
04A9
050E
0542
053B
04FB
049C
0458
045A
048E
04B8
04BF
04B9
04AF
0496
0480
04A3
04FA
0514
0491
03CE
03B0
0481
0530
042C
0110
FD47
FAC9
FA4E
FAF2
FB63
FB2B
FAC3
FABB
FB20
FB96
FBCF
FBBD
FB7C
FB35
FB06
FAF9
FAFA
FAF9
FB0E
FB54
FBAB
FBC3
FB74
FB0C
FAFF
FB5B
FBAA
FB82
FB12
FAE4
FB2E
FB8D
FB99
FB78
FB94
FBD5
FBA3
FADE
FA91
FC2A
FFCC
03C4
05FB
05E6
04CF
0442
048F
04F7
04EA
04A4
049E
04DB
0502
04F3
04DF
04E5
04DC
04B1
0495
04B7
04EE
04EF
04BF
04AA
04C9
04D8
04AB
0482
04AE
04FC
04E2
044F
03DF
0411
0494
04CB
04B8
04E8
0550
04CB
025B
FEA1
FB92
FA82
FAE1
FB38
FAF5
FAC2
FB30
FBCD
FBCB
FB28
FAA6
FABD
FB0A
FB07
FACF
FAE5
FB5F
FBC8
FBCB
FB98
FB86
FB8A
FB62
FB14
FAF4
FB1E
FB49
FB36
FB1A
FB47
FBA3
FBBB
FB7A
FB53
FB89
FBA8
FB1F
FA6A
FB05
FDDF
01F4
0502
05B4
04D5
0439
04B2
057B
058D
04F5
0494
04DE
054E
053C
04C2
0482
04BA
0504
04F6
04BC
04C1
0502
0511
04B4
043C
0417
0442
0464
045C
0462
0495
04BC
04A9
04A2
0504
057B
04FB
02C9
FF6F
FC6C
FAD3
FA7B
FA90
FAA9
FAF7
FB95
FC0D
FBDF
FB37
FAD0
FB0A
FB7C
FB7B
FAF8
FA81
FA85
FAD7
FB0E
FB17
FB32
FB75
FB9E
FB79
FB42
FB53
FB9E
FBB4
FB68
FB22
FB55
FBC7
FBC0
FB1E
FAEC
FC7A
FFDC
0382
0598
05BC
0514
04E0
0539
0563
04FB
0473
045C
04A3
04C1
0481
043D
0446
047D
04A0
04C0
0517
058A
05A8
0542
04BA
0487
0499
048B
044C
044C
04C1
052F
04FC
045F
0445
0505
0596
046A
0126
FD40
FAB3
FA37
FADB
FB44
FB02
FAA4
FABF
FB37
FB8D
FB86
FB62
FB6C
FB94
FB9D
FB7B
FB5A
FB55
FB51
FB36
FB1B
FB21
FB34
FB2F
FB20
FB3C
FB7B
FB79
FB04
FA96
FAE8
FBED
FC95
FC00
FAD4
FAEF
FD7B
0186
04C3
05C4
0524
048A
04C8
0549
053A
04AF
0475
04E5
056F
055B
04AC
040E
03F5
042D
0452
045E
0490
04E6
050D
04DA
0494
0497
04D8
0505
0503
0509
052A
0519
04A5
043A
047C
053C
0530
0329
FF82
FC18
FA94
FAEE
FBB9
FBC3
FB1E
FA9C
FAA2
FAD1
FAC3
FA9C
FABC
FB1F
FB63
FB5C
FB4E
FB76
FBA7
FB98
FB6B
FB83
FBE5
FC07
FB90
FAF0
FAD5
FB33
FB4F
FADE
FA9D
FB43
FC42
FC31
FABE
F996
FAD5
FEAD
02F9
055E
0570
0497
043F
049A
0506
051A
0505
0515
054B
056E
0553
0504
04A9
0474
0484
04D2
0528
054E
0534
04F9
04B7
0478
0443
0431
0457
04AC
04F0
04DC
0470
041C
0472
056E
0618
0518
01FD
FDF0
FAF1
FA1D
FAD1
FB81
FB52
FABA
FA9A
FB1A
FB99
FB8D
FB25
FAF3
FB2D
FB7A
FB76
FB2A
FAED
FAF3
FB1D
FB30
FB1E
FB06
FB09
FB32
FB75
FBAB
FB9E
FB39
FAC3
FAB6
FB31
FBAD
FB84
FAEA
FB1A
FD31
00CF
0421
058D
052A
0478
04A5
056E
05CF
0566
04D5
04C9
0522
0545
0502
04C3
04DB
0506
04D4
0463
0445
04B4
0536
0537
04C6
0473
048C
04CA
04DA
04D3
04E9
04EE
048B
03FE
0417
0510
05B2
0447
0095
FC7F
FA4A
FA6B
FB5D
FB87
FAD3
FA4D
FA92
FB2A
FB4D
FAE4
FA72
FA63
FAA8
FB02
FB49
FB6B
FB5C
FB2F
FB19
FB3B
FB71
FB75
FB3D
FB11
FB2A
FB56
FB33
FAC0
FA7F
FADC
FB88
FBAB
FAF5
FA58
FB60
FE92
0298
0552
05D2
0513
04A5
0502
0573
0553
04EE
04E8
0540
0562
0511
04C8
04FF
0576
0593
0534
04C9
04AD
04C5
04CE
04C4
04CB
04D6
04B9
048B
04A2
0512
0563
051E
047D
044B
04F2
05BD
0549
02CF
FF04
FBB5
FA4D
FAAD
FB76
FB7A
FAC1
FA31
FA5B
FAEC
FB3E
FB2C
FB0C
FB10
FB0B
FAD8
FAAB
FAB3
FAC5
FAA1
FA6B
FA84
FAF3
FB4B
FB42
FB1A
FB36
FB78
FB6F
FB15
FAF8
FB5F
FBB0
FB2C
FA2D
FA30
FC5D
0036
03E2
05D2
05E9
0538
04CC
04E7
052F
054B
0539
0529
052F
052D
0507
04D9
04E6
053E
0593
058B
0524
04BF
04B7
050A
056B
0597
057D
0531
04DA
04AF
04D1
0513
051C
04E0
04D2
0542
058E
0462
0126
FD0E
FA46
F9D9
FAC7
FB4E
FAD7
FA3C
FA58
FAF1
FB43
FB27
FB1D
FB57
FB5E
FAE2
FA5F
FA7F
FB1E
FB72
FB20
FAAA
FAAB
FAFC
FB10
FAD6
FAC8
FB18
FB4E
FB12
FACE
FB1A
FBBD
FBCE
FAFB
FA43
FB22
FE0C
01E0
04E2
061D
05E0
0527
04B6
04A9
04B3
04AC
04C5
0531
05AF
05B9
053A
04B7
04A7
04E2
04F6
04D5
04D4
050B
052A
0501
04E7
0530
057D
052E
0468
0418
049A
051C
04CB
042A
046F
0589
05AB
034B
FF23
FB97
FA3C
FA8B
FB0C
FB1C
FB09
FB15
FB10
FAE2
FAD2
FB0E
FB51
FB43
FAFD
FADA
FAF0
FAFD
FADB
FABF
FADC
FB09
FB0B
FAF3
FB07
FB4E
FB87
FB82
FB56
FB3E
FB54
FB80
FB84
FB2F
FAA9
FAB5
FC4A
FF91
034D
05AE
05F7
0523
04AD
04FC
0553
0518
04A3
0496
04F0
0524
04FD
04E6
0531
058A
056F
04F3
049F
04A2
04A1
0465
0450
04CB
0576
0577
04A8
03E8
0408
04B2
04E6
046D
043A
0500
05E4
051D
01F7
FDD2
FADA
FA08
FA90
FB19
FB15
FADE
FAE8
FB29
FB48
FB17
FAC9
FAB0
FAE2
FB2F
FB5A
FB57
FB51
FB6B
FB90
FB94
FB71
FB4A
FB2E
FB12
FB03
FB2E
FB8E
FBD3
FBC7
FB9F
FBA6
FBA7
FB24
FA55
FA8C
FCEC
00D2
0416
0531
04B2
0443
04A1
0523
0511
04AC
04A4
04FA
0515
04CB
049C
04E0
052E
0503
0499
048F
04EF
0513
04A3
0424
044F
0507
0572
050C
0451
0411
046C
04BC
0488
0432
0473
0545
0581
03DD
0059
FC9B
FA96
FAC0
FBC7
FC1B
FB7D
FAE4
FB12
FBB0
FBEA
FB8F
FB2B
FB32
FB78
FB94
FB78
FB5E
FB53
FB2F
FAF6
FAE3
FB11
FB40
FB31
FB07
FB0C
FB3D
FB40
FAF7
FAD1
FB38
FBD8
FBCF
FAE3
FA2E
FB48
FE96
02A2
0556
05D5
0506
045B
0461
04A2
04A2
0482
0492
04BF
04B4
046C
0443
0476
04D0
04FF
04FC
04F8
04ED
04AB
0446
0432
04AF
055C
0594
0535
04BC
049D
04BE
04BA
048D
04AF
0560
05F3
051A
0226
FE03
FABC
F9C3
FAAF
FBC1
FBBC
FB01
FAC0
FB53
FBE2
FBAE
FB15
FAF6
FB72
FBD4
FBA1
FB39
FB35
FB81
FB92
FB41
FAFC
FB08
FB19
FADE
FA9D
FACA
FB3D
FB60
FB0F
FAE0
FB40
FBB5
FB71
FA9D
FAA0
FCBE
0092
0437
05FB
05CD
04FB
04C0
0534
0595
055C
04D4
0498
04C1
04DB
04A3
045F
0474
04C7
04E9
04BA
0495
04C5
0511
0516
04E1
04CD
04EB
04E4
049A
0473
04B5
04F6
04A1
0404
0425
0547
060E
04A6
00E2
FCB1
FA46
FA0C
FAAF
FAE3
FAA5
FAA7
FB1A
FB6C
FB28
FA9B
FA71
FAE0
FB75
FBA9
FB75
FB2E
FB10
FB14
FB2A
FB53
FB81
FB7F
FB35
FAE1
FADF
FB32
FB74
FB59
FB27
FB5A
FBE1
FC03
FB54
FA95
FB45
FE1A
020B
0516
060C
0582
04F7
0536
05BE
05B1
04FE
0460
045C
04A6
04AF
0476
0473
04D8
0537
051B
04AA
046D
048E
04B9
04BC
04D2
052D
057F
0562
04F2
04A5
049C
0481
0437
0435
04D0
0561
049E
020B
FEA0
FBDE
FA79
FA27
FA5E
FAC6
FB24
FB46
FB33
FB25
FB3A
FB4A
FB34
FB1E
FB3E
FB6E
FB55
FAF7
FABF
FAEA
FB2E
FB32
FB06
FAE9
FADF
FADD
FB0A
FB83
FBEB
FBB8
FB0C
FABB
FB2D
FBA5
FB59
FB03
FC6E
001C
0425
061E
05B7
04B2
048A
0504
0532
04FC
0500
0559
0562
04D1
044C
047D
0524
0581
0564
0536
0536
0533
0511
0500
0515
050C
04B4
0455
0454
0491
04A4
0497
04DD
054B
04C0
025D
FECF
FBD7
FA88
FA78
FAAD
FAC2
FAE0
FAFF
FAD0
FA59
FA1A
FA64
FAE3
FB1A
FB0C
FB0E
FB2A
FB21
FAF5
FAF5
FB36
FB5A
FB1F
FAE0
FB17
FB96
FBB0
FB3D
FAE1
FB0E
FB50
FB20
FB1C
FCA1
FFFB
0393
0576
055B
04AA
0499
04FA
0513
04E6
050B
0597
05EE
05AE
053E
052C
0566
0575
053A
0507
0502
04ED
04A5
0468
0462
0462
0451
0480
0516
0580
0521
0463
0465
0539
0529
0292
FE37
FAD3
FA24
FB23
FBB4
FB2F
FA95
FAAF
FB13
FB1B
FAE4
FAE8
FB12
FAEE
FA87
FA68
FAA8
FABF
FA73
FA5D
FAF3
FBB6
FBE1
FB8C
FB62
FB87
FB79
FB18
FB04
FB7D
FBAE
FAE0
FA14
FB58
FF27
0361
0592
0583
04E2
04D8
050D
04E5
04A7
04E8
0572
0587
0509
04A6
04CD
0525
0542
054E
0582
0593
052C
04AA
04AB
050E
0515
0493
044A
04BE
054E
0514
0467
047D
0562
054B
02AF
FE7E
FB56
FAB0
FB83
FBEA
FB58
FAB1
FABA
FB30
FB71
FB59
FB2D
FB03
FACA
FA9D
FAA6
FAC7
FAB4
FA73
FA61
FAA5
FAF0
FB01
FB08
FB4B
FB8D
FB5B
FAD9
FABD
FB30
FB5E
FAB0
FA2B
FBAA
FF8C
03C3
05C4
0530
03F0
03D6
04CA
0592
0590
0534
04FA
04D0
0493
047B
04BF
0523
0540
0529
053E
0580
0585
0530
04F6
051E
054B
0516
04C6
04DD
0533
052C
04C9
04D1
0570
054C
02E1
FEAB
FB16
F9EF
FA9C
FB4F
FB4B
FB2F
FB78
FBAE
FB4C
FAAA
FA79
FAC5
FB05
FB08
FB22
FB6A
FB72
FB09
FAAC
FAC7
FB05
FAE7
FAA3
FAD2
FB54
FB69
FAE4
FA97
FB11
FB94
FB23
FA6B
FB7C
FF2C
0390
05E5
058E
0458
0413
04BE
0543
0526
04DA
04CD
04E6
04F9
0522
056A
0579
051A
04A8
04A3
04F7
052F
0527
0527
0548
0542
04F2
04B6
04E0
0520
04FB
04AE
04F5
05A7
0546
0290
FE52
FAEF
F9FC
FAD3
FBA9
FB9A
FB1E
FAE9
FAFA
FB06
FB1B
FB65
FBAA
FB7F
FAF2
FA8D
FA9E
FAD5
FAD2
FAB5
FAD2
FB15
FB21
FAF9
FB0B
FB6E
FBA0
FB4C
FAE6
FAFC
FB41
FB08
FAA9
FBAC
FEF3
0329
05D5
05F9
04EE
047B
04DC
051E
04D2
0482
049A
04C3
0491
044B
0479
0505
0557
0539
050F
0519
0516
04DF
04CA
050C
0539
04EB
047D
0493
0502
0504
048B
0488
0558
0589
033A
FEBB
FAC2
F989
FA87
FB92
FB99
FB44
FB55
FB94
FB7F
FB3A
FB37
FB56
FB29
FAD1
FAEA
FB70
FB95
FAFA
FA67
FAB7
FB8F
FBE9
FB85
FB15
FB0C
FB11
FAD8
FAC9
FB41
FBA4
FB2A
FA7D
FB88
FF17
0370
0602
0615
050D
0468
044C
0437
042A
0479
04F6
0506
0496
044D
049E
0526
0555
053E
0539
0530
04D0
044E
0445
04C6
0519
04C9
0461
04A2
054D
056E
04E0
049A
0505
04DA
0281
FE61
FAE4
F9E8
FADF
FBCF
FBB5
FB37
FB33
FB91
FBBF
FBA9
FB98
FB89
FB43
FAED
FAFC
FB67
FB8C
FB15
FA92
FAB5
FB4B
FB82
FB2A
FAF8
FB60
FBDB
FBC2
FB4C
FB17
FB17
FACD
FA94
FBC6
FF08
02F6
0560
05A3
0517
050C
0549
0502
045E
0439
04B7
050D
04C3
045B
0470
04C1
04B6
0468
0479
04F9
053B
04F8
04CA
0526
0585
053A
0493
0456
047D
0458
03EF
0441
0583
05F6
039D
FF02
FB1C
FA0D
FAF6
FB92
FB1C
FA9D
FADF
FB63
FB76
FB50
FB7D
FBC7
FB90
FAF0
FAAC
FAFF
FB39
FAE9
FAAC
FB22
FBCD
FBB6
FAF1
FA8D
FB10
FBC4
FBDD
FB8F
FB78
FB72
FAF2
FA7F
FBAE
FF19
0319
0555
0550
048F
047A
04EC
050C
04C0
04A9
0504
0550
052C
04E5
04E5
050E
0508
04DF
04D5
04DD
04B4
046B
0462
04A0
04B6
0472
044A
04A7
0519
04E6
0451
046E
055A
056B
02FE
FEC1
FB55
FA70
FB27
FB6F
FABB
FA3A
FACB
FBB5
FBD1
FB21
FA97
FAA4
FADE
FAE7
FAFD
FB5A
FBAC
FB91
FB51
FB75
FBDD
FBDA
FB4B
FAEA
FB33
FB9E
FB74
FAEB
FAC2
FAFE
FAF8
FACC
FBD5
FF04
0326
05CE
05F7
04FA
049B
0504
0536
04DA
0498
04E3
0546
0532
04D9
04C1
04EE
04EE
04A2
0465
0464
045D
0436
0446
04AB
04EF
04CA
04B1
051D
0594
053A
0451
0428
051A
0569
030F
FE89
FAC3
F9E0
FB01
FBD0
FB6A
FACE
FAE5
FB45
FB2D
FAC1
FAB2
FB18
FB5B
FB38
FB12
FB35
FB57
FB3A
FB2D
FB7C
FBC7
FB85
FAF2
FAD1
FB4F
FBBD
FBA3
FB65
FB85
FBA7
FB27
FA92
FB8A
FEC3
02B8
0524
056A
04E8
04F7
056E
0566
04BD
0437
0450
04A6
04B5
0494
04A7
04F0
0522
052A
052E
052E
04F9
049D
0472
0495
04B3
0490
0479
04C2
050D
04B4
03F0
03D4
04B3
0517
0332
FF38
FB83
FA22
FAC2
FB7F
FB52
FAE1
FB0F
FBA1
FBCF
FB7D
FB3E
FB58
FB77
FB56
FB1D
FAFE
FAE1
FAB6
FAC5
FB3C
FBB2
FB92
FB03
FAC9
FB26
FB85
FB7D
FB81
FBF8
FC3E
FB81
FA80
FB4E
FEDC
035B
05F6
05E2
04DD
04A5
0509
04F3
045D
0437
04C1
0527
04D8
045B
0470
04F0
0521
04E1
04B8
04D8
04D1
046D
0432
0487
04FB
04F7
04B5
04D2
0529
04FC
0449
0409
04A2
04BE
02A8
FEB1
FB42
FA34
FAE5
FB68
FB01
FA83
FAB8
FB50
FB9C
FB7F
FB41
FAFC
FAAC
FA9D
FB1D
FBCD
FBDE
FB41
FAE2
FB66
FC2F
FC3F
FB9A
FB16
FB0E
FB06
FAC7
FAF1
FBDC
FCA0
FC22
FB0D
FB97
FECB
02ED
0552
055C
04B5
04DD
0580
058F
050E
04E8
0562
05AE
0533
047A
0451
04A8
04D7
04B6
04AD
04D6
04C2
0443
03DF
0419
04A9
04DF
049E
0464
0464
044A
0417
0461
0535
0543
0319
FF20
FB97
FA46
FABE
FB42
FAF9
FA7B
FA79
FAC0
FAE5
FB09
FB6C
FBAE
FB4C
FA96
FA6F
FB0B
FB9B
FB7E
FB29
FB65
FC0B
FC41
FBD7
FB8E
FBCD
FBF3
FB6B
FAC8
FAEB
FB92
FBB9
FB74
FC48
FF1D
029A
0483
046F
0425
0507
064E
0668
054F
046F
0498
051F
0526
04D5
04D0
050C
04F1
0467
040D
0443
049E
04A8
0498
04C6
04F1
04A6
0414
03E1
042F
0479
0476
048A
04E6
04BA
02EF
FFB6
FC9F
FAF6
FA8E
FA78
FA5E
FA7F
FAD3
FAE7
FAB1
FABF
FB5A
FBF9
FBF1
FB79
FB5A
FBC5
FC08
FB9E
FAFB
FAD7
FB31
FB7B
FB86
FB9D
FBC8
FB9F
FB13
FACD
FB3A
FBBA
FB67
FAC7
FBB8
FF30
039F
064E
0637
04DF
0443
04AF
050B
04AF
042C
0439
04A8
04CE
048C
0460
0491
04D5
04D3
04A0
047E
0473
0464
0465
049C
04DF
04C1
0437
03E4
0461
0558
0593
0419
0111
FDA6
FB26
FA2F
FA73
FB1D
FB74
FB5B
FB32
FB4C
FB7F
FB6B
FB0A
FAC7
FAEE
FB44
FB63
FB47
FB3E
FB75
FBC9
FC0C
FC2F
FC24
FBD3
FB61
FB44
FBA9
FBFF
FB95
FAE3
FB82
FE69
0272
0540
05A9
04C6
0460
04EA
0561
04FF
043D
0405
0473
04E1
04F0
04EB
0522
0566
055A
0503
04AA
0461
03FD
0392
0394
0439
04F8
0509
0472
041E
04B2
056B
04A3
0199
FD82
FA8D
F9E1
FAAE
FB57
FB2B
FAC8
FAF2
FB8B
FBE5
FBBD
FB72
FB60
FB5E
FB21
FACD
FACD
FB35
FBA3
FBC9
FBC7
FBCB
FBB4
FB58
FB02
FB2B
FBAD
FBAE
FAC9
F9FE
FB02
FE5B
028E
0566
0601
0552
04D0
04FE
055E
0565
0516
04BC
0474
043B
042E
0479
04F2
051F
04C1
043A
041F
047A
04B9
0479
041C
044E
0509
0584
053C
04C2
04FB
059D
0513
0238
FDF5
FAA9
F9D3
FAB3
FB6A
FB1A
FA79
FA73
FAF5
FB45
FB28
FB1C
FB72
FBCF
FBAF
FB2B
FAD1
FAEA
FB3B
FB80
FBBC
FBE9
FBBE
FB1B
FA86
FAB3
FB7D
FBD0
FAFD
F9ED
FA7D
FD81
01B9
04FB
0638
060C
0597
054B
04FE
04AA
04A2
04FC
054A
051E
04A3
0467
0497
04D5
04CA
04A9
04D9
0544
0562
04F5
047B
048C
0504
0521
0498
042A
04B3
05BC
058A
02D7
FE73
FABE
F975
FA37
FB4A
FB80
FB1D
FAFA
FB50
FBA2
FB89
FB25
FAD1
FAB2
FABF
FAFE
FB66
FBAB
FB79
FAEF
FA9E
FAD3
FB2F
FB2A
FADD
FAE5
FB6A
FBB8
FB28
FA57
FAE5
FDBE
01DF
0520
0630
058D
04A8
045C
047E
0493
0487
0493
04C0
04D9
04CC
04CC
0507
0553
0565
052F
04EC
04C3
04A0
0477
047B
04DE
055C
055C
04BF
043F
04A1
057D
0540
02BB
FEA5
FB21
F9CD
FA62
FB60
FBBA
FB92
FB75
FB7F
FB71
FB46
FB3C
FB59
FB4E
FAF5
FAA2
FAB2
FAFD
FB07
FABC
FAA6
FB29
FBD8
FBEE
FB51
FAC7
FAF7
FB87
FB93
FAFF
FAF3
FCBF
0050
03FF
0603
05FD
050B
047B
049C
04D4
049D
0428
0402
0458
04D0
0507
04FD
04F2
0505
0520
052D
052E
0526
050B
04DF
04C2
04B6
048F
0440
042E
04C5
059D
0565
0319
FF51
FBF3
FA74
FA87
FAD6
FAB0
FA9B
FB38
FC2A
FC83
FC03
FB62
FB4E
FB8D
FB7F
FB14
FADF
FB26
FB6C
FB23
FA8D
FA6A
FAF0
FB77
FB62
FAF4
FAE4
FB46
FB6B
FAFB
FADA
FC6C
FFEB
03D7
0638
066C
0575
04B9
04A7
04B8
0472
0409
03F9
0455
04B3
04B9
0485
046D
0494
04D1
04F6
04FE
04F5
04E3
04DF
050A
0559
0572
051A
04AC
04CE
0575
056C
035C
FF6E
FB8D
F9B0
FA03
FB01
FB51
FB16
FB35
FBD3
FC25
FBA5
FAEB
FAE2
FB8E
FC0A
FBBF
FB20
FAF4
FB4C
FB8C
FB5D
FB0F
FAF9
FAE9
FA8E
FA2B
FA5A
FB11
FB76
FB0B
FAC1
FC3C
FFE0
03FD
064F
062E
04FA
045C
04A8
0504
04DB
0488
0499
04F8
051A
04D9
0499
04A3
04BC
048E
0447
045F
04E1
0550
0553
052A
0537
0557
0514
0480
0453
04DD
0527
03BA
0058
FC97
FA73
FA66
FB2E
FB67
FAF0
FA9F
FAEE
FB6E
FB80
FB25
FAE2
FAFC
FB3B
FB5A
FB69
FB8E
FBA5
FB64
FADD
FA8D
FABB
FB15
FB21
FAFD
FB32
FBCA
FC00
FB4F
FA9E
FBB4
FF33
0376
0600
05F8
04D4
0475
051F
05A7
054D
04A1
0488
04F3
051F
04CC
048E
04D8
053D
0516
0484
044B
04BB
053E
052E
04B1
0467
0481
049A
0483
04A6
0542
058A
042C
00D6
FCE3
FA3A
F99D
FA3C
FAD5
FAEC
FAD8
FAF1
FB1F
FB22
FB01
FAF2
FB00
FB03
FAEF
FAFC
FB52
FBB3
FBB6
FB53
FB02
FB2A
FB95
FBB6
FB6E
FB2F
FB45
FB4F
FAE0
FA7F
FB91
FEC2
02E0
05C0
065F
05C0
0578
05DC
0605
0566
04AB
04BB
056B
05B8
0532
0485
047D
04EC
050A
049B
042F
0442
0492
049B
0464
045C
049E
04C5
04A0
049E
051C
057A
046E
0171
FD93
FAA2
F993
F9E0
FA5F
FA73
FA50
FA58
FA91
FAC0
FAD2
FAEE
FB26
FB51
FB44
FB1B
FB20
FB6A
FBB0
FBAF
FB7E
FB6D
FB85
FB8A
FB68
FB6D
FBC0
FBED
FB6B
FAB6
FB4E
FE31
0262
0594
066E
05C1
0545
058D
05CC
055D
04C7
04DE
0578
05A1
04FD
0455
0476
0513
053E
04B7
0436
0462
04FB
054E
0526
04D5
0490
0431
03C1
03C1
047A
0529
0462
017F
FD8B
FA7B
F981
FA2F
FB1F
FB5C
FB0C
FADA
FB0D
FB49
FB2D
FADC
FACD
FB25
FB7C
FB67
FB00
FAC7
FAF0
FB34
FB3F
FB1C
FB04
FB00
FB0B
FB4D
FBE3
FC67
FC38
FB84
FBB9
FE26
023A
05A1
068D
0583
047B
048B
0509
04FC
0489
0484
04FD
0523
0492
040C
046A
0559
05BF
0538
0486
0476
04D6
04F2
04A9
047E
04AA
04B9
0457
0401
0456
04EF
0469
01E8
FE3B
FB3E
FA25
FA94
FB42
FB54
FAF7
FAD1
FB2B
FBAD
FBD6
FB91
FB3E
FB34
FB57
FB49
FAFB
FAC9
FAFE
FB64
FB8D
FB5C
FB1C
FB13
FB3C
FB72
FB9D
FB98
FB2D
FA9B
FAEC
FD31
0116
04AF
0629
0595
0496
0470
04DE
04F5
049C
0481
04DE
0517
04B3
0432
0453
04F2
0531
04B9
0431
044A
04CB
0507
04E4
04E5
0534
0540
04B3
043A
04BE
05D6
05C1
033A
FF10
FB8A
FA38
FAAD
FB63
FB6F
FB1E
FB10
FB4C
FB60
FB20
FAE4
FAF9
FB39
FB4A
FB2A
FB32
FB8F
FBF5
FBF8
FB98
FB32
FB00
FAE5
FAC8
FAD5
FB1B
FB34
FAB5
FA08
FA79
FCF9
00E0
0442
05A7
054A
048C
046A
04C3
04FA
04DD
04C3
04F0
053E
055C
0531
04E0
048E
044B
0431
0462
04C4
04FF
04DC
049E
04BA
0532
0577
0524
04B3
04FC
05DC
05CF
0361
FF11
FB43
F9F8
FAE1
FBF8
FBD2
FAE9
FA80
FAF1
FB79
FB72
FB25
FB24
FB60
FB58
FAF5
FAB3
FAF0
FB6D
FBAC
FB94
FB6B
FB51
FB25
FAEC
FAF8
FB6D
FBC3
FB46
FA36
FA04
FC08
FFF8
03DD
05D2
05AF
04E6
04C0
052A
0545
04D5
048A
04EC
0587
058D
04F2
0479
04A1
04FF
04EA
046F
0431
046D
04B2
049E
0477
04A1
04E9
04DB
049B
04DB
05A6
05CE
03F9
004D
FC8C
FA6E
FA18
FA6D
FA90
FA94
FADE
FB52
FB79
FB37
FAF3
FB0A
FB49
FB39
FAD5
FAA6
FB0B
FBAC
FBE3
FB96
FB4F
FB6D
FB99
FB55
FAD8
FAD5
FB60
FB98
FAF8
FA92
FC37
0021
0436
061A
0598
0486
0470
0524
058B
0543
04D9
04BE
04CC
04D2
04F2
0534
053D
04E1
048B
04AD
0507
0505
04AA
0480
04B1
04B4
0444
0407
0495
0515
03CD
0053
FC72
FA55
FA49
FAEF
FB25
FB02
FAFE
FB0F
FAED
FABD
FACF
FAFE
FAE6
FAAE
FAE9
FB92
FBDB
FB5A
FAC6
FAEB
FB74
FB78
FAFE
FAFD
FBC0
FC35
FB94
FB06
FC96
006D
0433
05AA
051A
0476
04BF
0541
052E
04DA
04FA
056C
057F
0513
04BC
04D2
04F8
04E2
04D5
0507
0519
04AD
042C
0446
04D0
04F9
049A
048D
0534
054E
0332
FF26
FB84
FA38
FAC5
FB51
FB07
FA96
FAB0
FB06
FB0B
FAE1
FAFC
FB40
FB2D
FAD1
FAD1
FB53
FBA2
FB3E
FAB8
FADE
FB83
FBCD
FB8D
FB69
FBA5
FB8E
FACB
FA99
FCAC
00C9
0484
05D4
0535
049C
04F5
057E
056D
0515
051E
0566
054E
04D6
0499
04C5
04D6
0483
0448
0492
04F0
04C9
0457
044F
04B3
04D4
048B
0497
053C
0530
02DE
FEB3
FB21
FA02
FAB7
FB62
FB44
FB0F
FB44
FB68
FAFF
FA7A
FA8F
FB1E
FB61
FB1D
FAE6
FB1E
FB6C
FB6B
FB54
FB73
FB87
FB43
FB0B
FB6E
FC08
FBD2
FADC
FAEA
FD89
01D9
052E
05F0
051A
048F
04CB
0502
04CE
04B1
04F4
0516
04A8
0427
0450
04F8
0548
04FB
04B6
04EB
052B
04F8
04A7
04C0
04FD
04B8
0423
0434
04EF
04B3
0202
FDB0
FA62
F9B9
FABE
FB76
FB3F
FAF2
FB30
FB90
FB88
FB46
FB43
FB76
FB7A
FB4A
FB41
FB6A
FB67
FB18
FAE8
FB1A
FB53
FB36
FB0F
FB52
FBAC
FB68
FAD1
FB71
FE52
0268
0568
0626
0590
051F
0526
0513
04BB
0493
04C6
04E7
04AD
0471
0494
04E0
04DE
04A2
04AA
04FE
0515
04BD
047C
04AD
04D9
047D
041C
0494
0574
04E0
01B6
FD4B
FA4A
F9E4
FAD6
FB49
FAE5
FA93
FAD9
FB50
FB7D
FB73
FB70
FB62
FB28
FAF3
FB02
FB31
FB2E
FB0A
FB1F
FB61
FB59
FAFB
FAF3
FB99
FC25
FBB0
FAD8
FB8B
FEBF
02EF
058A
05A2
04A0
044A
04D7
0552
0535
04E8
04E2
0501
04F2
04BF
04AA
04C2
04E5
0508
0530
0537
04FB
04B6
04C8
050E
04EB
0447
03FC
04A7
0559
0436
00B4
FC9F
FA67
FA97
FB94
FBB5
FAFE
FA80
FABA
FB2F
FB50
FB27
FB05
FB03
FB09
FB0E
FB0C
FAE7
FAA9
FAA8
FB1C
FBA0
FB98
FB24
FB12
FBA3
FBF1
FB3E
FA77
FB94
FF2F
036B
05C3
05A3
04A2
045A
04CB
0514
04F0
04D1
04F1
050B
04F5
04EC
0518
053A
0518
04EB
04FE
0520
04F0
0496
049A
04F7
04FD
047D
0454
051F
05C7
0457
006F
FC2C
FA0F
FA6F
FB82
FBB7
FB2F
FAD7
FAEE
FB06
FAFC
FB11
FB49
FB49
FAFA
FAC1
FAE5
FB25
FB26
FB06
FB18
FB38
FB08
FAB5
FADF
FB78
FB87
FA9E
FA1A
FBE6
0009
042E
0603
058A
04A2
04A5
0538
056F
052F
04FC
0500
04F0
04BB
04AA
04D3
04E9
04C4
04AD
04E3
0529
0520
04E5
04E2
050D
04F0
0496
04B6
057D
05AA
03AB
FFAA
FBCC
FA1A
FA8A
FB6B
FB75
FADD
FA7B
FA93
FAD9
FB12
FB3F
FB51
FB2E
FB03
FB19
FB5A
FB5F
FB0E
FAD9
FB12
FB5E
FB36
FAD4
FAEE
FB84
FBA6
FAEE
FAA3
FC7E
006A
0434
05CD
055A
049F
04C2
0554
0573
051D
04E5
04F9
0504
04D8
04AB
04A4
04AD
04B3
04CD
04F3
04E3
0498
0480
04E6
054F
0504
0448
0436
050B
0543
032D
FF2C
FB9B
FA4E
FAD0
FB5E
FB1C
FAA4
FAAA
FAFC
FB15
FB03
FB1E
FB5B
FB60
FB30
FB24
FB4B
FB53
FB1D
FB00
FB33
FB5F
FB27
FAE0
FB25
FBB9
FBAE
FAEE
FAF4
FD35
0128
048E
05CF
0569
04E9
0504
0543
0529
04EB
04E3
04F5
04DA
04A9
04A1
04A9
048A
046C
04AB
052D
0562
0511
04BA
04D4
050C
04C6
0442
0466
052C
0508
028E
FE70
FB12
FA12
FAC7
FB6C
FB3A
FACA
FACB
FB0C
FB0D
FAD9
FAD8
FB1D
FB57
FB5E
FB52
FB49
FB2A
FB02
FB0B
FB42
FB47
FAF1
FABF
FB32
FBD1
FB9B
FAB2
FAD5
FD7E
01CF
052A
05EE
0501
0465
04D6
0575
056D
0508
04E8
0507
04FE
04D5
04E5
0521
051B
04BF
047F
04A7
04E8
04EE
04EA
0523
0546
04D4
0434
0465
054C
0520
0263
FE09
FABB
F9FD
FAC3
FB29
FABC
FA73
FADD
FB5E
FB54
FB0E
FB1D
FB58
FB38
FAD1
FAB2
FAFA
FB30
FB17
FB02
FB2B
FB41
FB00
FAD2
FB37
FBBB
FB71
FAAB
FB34
FE30
0259
0530
05B3
0514
04D8
0527
0546
0509
04EE
0515
0508
049F
046F
04D7
0554
0540
04D4
04BE
0502
0510
04C9
04C1
052C
0557
04C0
0425
0495
057F
04C8
0162
FD05
FA72
FA74
FB6F
FBA6
FB13
FAAF
FAD4
FB07
FAFF
FB07
FB45
FB5A
FB14
FADD
FB14
FB62
FB46
FAF6
FB0A
FB73
FB7D
FAFD
FABF
FB4B
FBDB
FB62
FA81
FB4F
FEC5
0323
05AE
05A5
04A7
0461
04D5
0511
04D9
04BF
04FD
051F
04E2
04B7
04F8
0540
050A
0491
0473
04BB
04E0
04B5
04AB
04F4
050C
049C
0448
04D1
0578
045A
00D6
FCC3
FA93
FAAD
FB6D
FB72
FB04
FAFD
FB52
FB54
FAF7
FAE1
FB42
FB78
FB1E
FABE
FAF9
FB81
FBA1
FB57
FB33
FB52
FB41
FAF1
FB06
FBB3
FC07
FB39
FA61
FBAE
FF95
03C3
0599
050E
043E
0487
053D
0539
049D
0465
04CE
051F
04E8
049A
04AE
04E1
04CE
04A3
04BC
04E9
04C5
0481
04A4
0507
04E2
041D
03CC
04B3
05A1
0461
007A
FC2E
FA1E
FA8D
FB9F
FBCD
FB4C
FB05
FB2A
FB4E
FB47
FB56
FB85
FB84
FB40
FB18
FB42
FB65
FB2D
FAE2
FAF5
FB47
FB60
FB48
FB7C
FBF6
FBE8
FAFF
FA72
FC01
FFC1
03A0
057F
054F
04A4
049F
04F8
04FE
04B7
049E
04C6
04D2
04A6
0494
04BE
04D9
04B4
0494
04B9
04E5
04C8
049A
04C3
050D
04D3
041F
03EF
04C2
055A
03CF
0004
FC34
FA97
FB0F
FBC6
FB98
FB0B
FAF9
FB3F
FB36
FAE3
FAE5
FB52
FB83
FB1F
FAB3
FAE2
FB75
FBBC
FB8C
FB45
FB1D
FAFE
FAFD
FB5E
FBE4
FBC7
FAE3
FA94
FC7E
006B
0419
0595
0529
0480
0482
04C5
04C6
04B8
04E6
050F
04D6
047F
0498
050A
0528
04C9
0489
04CE
0518
04E0
047F
0495
04EE
04CC
0449
0466
055E
059A
0357
FF0F
FB64
FA4B
FB1C
FBD5
FB9F
FB31
FB39
FB63
FB2A
FAC4
FAC6
FB36
FB8B
FB7B
FB4D
FB44
FB43
FB27
FB20
FB51
FB77
FB50
FB1D
FB3F
FB78
FB2C
FA8E
FAEE
FD60
0138
0460
0566
04C7
0418
0433
04A8
04CB
04A2
04A9
0503
0543
0508
047F
0437
046E
04D2
04F5
04DE
04E3
0518
0516
049A
0415
0444
050A
0509
02F6
FF3E
FBF1
FAB4
FB2E
FBB5
FB5E
FAC5
FAE0
FB98
FC06
FBBD
FB42
FB2C
FB56
FB44
FB01
FB07
FB6C
FB9F
FB3A
FAB1
FACD
FB8B
FBF9
FB6B
FA94
FB0A
FD9F
015E
045C
056C
04F8
0448
0436
049E
04E8
04D6
04A2
0493
04A4
04B1
04BE
04E0
0501
04E2
0482
0447
0490
051E
0544
04C3
0444
0494
055E
051B
029A
FE8C
FB2C
FA25
FB02
FBE5
FBA5
FAD2
FAA4
FB50
FBE1
FB9D
FAEE
FABB
FB2E
FB93
FB6D
FB1C
FB34
FB94
FB99
FB2A
FAF9
FB78
FBFF
FB93
FA83
FA99
FD36
0182
0500
05FD
0521
045B
04A3
0548
0541
04A1
044F
04AC
0521
0504
0485
0451
049C
04F0
04EF
04D7
0500
052E
04D3
040D
03C9
049A
05A1
051C
0238
FE25
FB10
FA29
FAC5
FB67
FB52
FAEC
FAD9
FB21
FB58
FB45
FB2A
FB4B
FB82
FB7E
FB3E
FB1D
FB48
FB72
FB39
FACB
FAC1
FB45
FBAC
FB49
FA99
FB26
FDEE
01FF
0520
05F2
0529
0487
04E2
058E
0595
0502
04A0
04C5
04EE
049D
0425
0435
04D7
0550
051E
04AA
04AF
052A
055F
04EB
046F
04B1
054A
04B1
01ED
FDEE
FAE4
FA20
FAEE
FB9A
FB52
FAB5
FAA6
FB18
FB53
FB11
FADB
FB26
FB9F
FBA3
FB2C
FAD6
FAF8
FB28
FAEC
FA88
FAAC
FB5A
FBB3
FB28
FA8F
FB77
FE6F
023C
04F8
05C7
0554
04D3
04D5
0516
0522
04DD
0488
046B
0496
04DC
0509
050F
0500
04E3
04BB
04AD
04E9
055A
058D
053D
04CB
04DF
0545
04A8
01E6
FDBE
FA80
F9CB
FAEA
FBCE
FB6C
FA98
FA8D
FB46
FBBE
FB70
FAED
FAE6
FB3B
FB58
FB25
FB10
FB3F
FB49
FAE8
FA8A
FAC4
FB66
FB8E
FAD7
FA38
FB41
FE6F
026C
052D
05BF
04F4
045A
04A6
0545
0558
04D1
0466
0490
04FB
0511
04C9
049C
04C1
04E5
04B7
0478
04A6
052B
0562
04F9
047D
0495
04E0
0413
0177
FDF6
FB62
FAB5
FB41
FB9F
FB3C
FAAB
FAA4
FB16
FB62
FB45
FB20
FB51
FB9C
FB86
FB14
FADB
FB2F
FB99
FB78
FAF6
FADE
FB67
FBBD
FB27
FA6A
FB53
FEA1
02D0
056B
058B
0484
0425
04C6
055E
0525
0483
044D
04A5
04F4
04D4
048D
0494
04DB
04F1
04A8
0464
0487
04E0
04EA
048C
045B
04D3
0565
04A7
01CA
FDCB
FAC8
FA0C
FAE9
FBAD
FB77
FAD7
FAB2
FB18
FB68
FB58
FB3F
FB6E
FB9E
FB6D
FB08
FAF9
FB5D
FBA8
FB6C
FB00
FB0A
FB88
FBBC
FB3E
FADC
FBFA
FF01
02AF
0521
058A
04C3
0438
047F
050F
0533
04ED
04BF
04E2
0500
04CC
047A
0470
04A9
04B9
047C
0461
04CF
0566
0563
04B1
0433
0496
051C
041C
00F3
FD0C
FA99
FA67
FB46
FB96
FB0B
FA91
FAD2
FB5A
FB64
FAF8
FACD
FB32
FBA2
FB88
FB1A
FB06
FB6A
FBA1
FB39
FAA8
FAB7
FB55
FB96
FB09
FAAA
FC05
FF5F
032D
0579
05BC
050B
04B3
04F4
0538
051A
04DF
04ED
0527
0526
04D5
0496
04BA
0506
0505
04AE
047C
04C2
0527
0517
049E
0474
04F2
053E
03ED
00A3
FCC9
FA63
FA2A
FB0B
FB81
FB1F
FAA0
FAAF
FB16
FB35
FAE9
FAAD
FAE0
FB3E
FB4E
FB13
FB05
FB5A
FBA7
FB73
FAF3
FAD3
FB43
FB9B
FB47
FAEB
FC09
FF40
0335
05A7
05B4
049D
0433
04E2
059D
0583
04F7
04DD
054B
057D
050D
0489
0498
0501
0507
0489
0440
04A9
053B
051F
047A
0457
0519
058B
0400
0062
FC96
FAAB
FAD6
FB98
FB98
FAEE
FA84
FAB9
FB0B
FAFE
FAC7
FAE1
FB42
FB6C
FB32
FB05
FB4F
FBC9
FBD3
FB55
FAEF
FB1B
FB76
FB3F
FA81
FA6C
FC29
FF8B
0302
0503
0549
04C6
0488
04D0
0531
0548
0526
0512
0521
0525
04FD
04C4
04A7
04A2
048F
0469
0466
04A6
04EA
04DE
04A6
04CD
056F
05A0
041A
00B8
FCFB
FACB
FAA6
FB5D
FB90
FB13
FAB6
FAED
FB45
FB2A
FAC3
FAB0
FB19
FB81
FB82
FB58
FB69
FB97
FB6C
FAEB
FAB7
FB2E
FBB2
FB58
FA4D
FA14
FC0D
FFD2
036E
0530
051F
0490
048D
0502
0548
0524
04EC
04EB
04FC
04DF
04AD
04AA
04D5
04D5
0487
0448
048A
0522
055F
04F2
0477
04BF
0598
059A
0389
FFCC
FC43
FA92
FAB3
FB53
FB62
FAF7
FAC3
FB06
FB5A
FB62
FB41
FB47
FB68
FB56
FB0D
FAF2
FB47
FBB6
FBA8
FB17
FAA8
FADC
FB52
FB3E
FA9A
FA9B
FC8A
003C
03EB
05CF
05B7
04ED
04A9
04F4
051B
04D2
0484
0492
04C5
04B1
046C
046D
04CD
050C
04CA
0467
0483
0512
054F
04D2
0446
049E
059B
05A6
036B
FF71
FBCA
FA22
FA5F
FB1D
FB48
FAF5
FAC5
FAF9
FB44
FB5A
FB56
FB71
FB97
FB8A
FB4C
FB2B
FB4F
FB71
FB3B
FAD9
FAE1
FB78
FBE8
FB6D
FA67
FA6E
FCC0
00C3
0455
05C5
0554
049D
04C2
056E
05A3
0516
0472
0461
04C3
04FD
04CE
048D
0492
04C1
04C8
04A5
04A7
04E4
04FC
04A6
0445
0484
054C
055E
036F
FFB5
FC05
FA33
FA62
FB2E
FB54
FAE1
FAAC
FB03
FB5B
FB39
FAE4
FAEE
FB56
FB8E
FB51
FB0D
FB3B
FBA3
FBA8
FB3D
FB09
FB70
FBDE
FB70
FA63
FA46
FC74
0072
042F
05E9
05AB
04DE
04A9
0502
053C
0510
04D4
04D6
04F2
04DD
04A8
04A2
04D3
04E0
0492
0440
0463
04D6
04EE
0468
0401
049B
05CE
05D6
0358
FF1A
FB83
FA4F
FAFD
FBB2
FB5B
FA91
FA69
FB02
FB91
FB85
FB29
FB07
FB28
FB31
FB11
FB1C
FB75
FBBE
FB97
FB34
FB29
FB90
FBCA
FB4B
FA8F
FAE8
FD37
00D7
0405
0569
0530
049D
04A6
0523
0552
04EF
047E
048E
04F7
051F
04D4
048A
04A4
04E5
04CB
0466
044C
04BA
0522
04EE
0475
0491
0539
0509
02BA
FEDA
FB8C
FA6A
FB05
FBB2
FB80
FAEC
FACF
FB29
FB56
FB1A
FAE9
FB24
FB87
FB9B
FB63
FB4E
FB7C
FB89
FB2A
FABD
FADD
FB7E
FBCD
FB3D
FA78
FAF9
FD8A
0148
0452
0572
0510
047E
0494
050B
0532
04E0
048D
049C
04E3
04F4
04C1
0499
04AA
04C3
04AD
0494
04BD
0507
04FC
047A
0415
046B
0526
04FA
02DC
FF3F
FBE0
FA45
FA7E
FB51
FB92
FB28
FACD
FB06
FB86
FBA3
FB38
FAC6
FACC
FB2D
FB70
FB6B
FB62
FB82
FB8C
FB47
FAF8
FB0A
FB4F
FB2C
FABA
FB37
FDC2
01B2
04D7
05A4
04C0
040D
0472
0525
052A
04AE
048A
04EB
0532
04FF
04B7
04C6
04F0
04C4
046D
0479
04E2
0501
04A2
0478
04FB
053C
03AE
0024
FC6A
FA7F
FA95
FB43
FB5E
FB0D
FAFB
FB37
FB50
FB24
FB06
FB16
FB18
FAF7
FAFD
FB53
FB90
FB4B
FAD7
FAF2
FB9C
FBE2
FB35
FA93
FBB3
FEF6
02BE
0510
057D
0521
0504
0517
04DD
046F
045C
04C0
0511
04EF
04B0
04D0
0533
054B
04F9
04B4
04CF
04ED
04A6
0455
04AE
056C
050E
026E
FE5E
FB26
FA3C
FAF1
FB89
FB43
FAC1
FAC1
FB1C
FB42
FB23
FB20
FB42
FB2B
FAD1
FAB8
FB1D
FB72
FB26
FAA4
FAD9
FBB2
FBF7
FB0D
FA60
FC11
0042
0475
0628
056E
046D
0492
0542
0542
049A
044E
04BF
0534
050E
04B4
04D1
053F
0552
04F0
04B5
04EA
050C
04BB
0483
050A
05A2
048D
0118
FCDD
FA4A
FA20
FAF4
FB31
FACC
FAB8
FB44
FBBB
FB93
FB2F
FB2A
FB60
FB41
FACB
FA98
FAE8
FB39
FB18
FAE0
FB23
FB99
FB6D
FAB8
FAF3
FD66
015F
04A8
05D1
057D
0531
0574
0598
051E
0482
0470
04C9
04F1
04C2
04A7
04CF
04E6
04BA
04AE
0514
0576
0525
045D
0439
0512
057E
03AD
FFB3
FBD7
FA40
FACE
FB9B
FB54
FA77
FA38
FAD8
FB84
FB92
FB3A
FB02
FB03
FB01
FAF5
FB0B
FB39
FB3D
FB17
FB20
FB72
FB89
FAFD
FA8B
FBB3
FF01
02FA
0562
0581
04AB
0481
051E
0571
04F5
0465
048A
051C
053C
04C8
047A
04C5
0536
053C
0501
04F9
0509
04B9
043F
0470
0546
052E
02A1
FE56
FAED
FA24
FB12
FB9E
FB17
FA8C
FAD4
FB5E
FB4A
FAD9
FAF3
FBA0
FBEC
FB66
FAD3
FAF7
FB62
FB38
FAAB
FABA
FB77
FBB5
FADD
FA5D
FC39
0057
043A
05BA
053D
04AC
04F0
0551
051C
04C3
04F6
056C
0552
04A0
0430
047A
04F1
04F2
04C2
04FB
0564
0533
046E
0430
0517
05EF
04BB
0115
FCEB
FA8F
FA71
FB24
FB4D
FAEA
FAB8
FAF4
FB33
FB23
FAF6
FAFA
FB27
FB47
FB55
FB67
FB61
FB0D
FA9F
FAA8
FB47
FBBF
FB49
FA65
FABE
FD6F
0188
04BE
05B1
0517
049B
04E9
055A
053F
04D7
04BE
04F9
050F
04E0
04CD
04FE
050C
04AF
0458
049F
0541
0563
04DF
0498
0516
0547
0382
FFBD
FC04
FA61
FABC
FB60
FB33
FAB5
FAC4
FB38
FB4B
FADC
FA98
FADA
FB31
FB1D
FADD
FAF7
FB5A
FB73
FB2B
FB10
FB65
FB88
FAE9
FA55
FB7C
FEEF
0319
05AA
05D6
04DF
046A
04D5
0557
0554
0509
04F9
052C
054B
0532
0509
04F1
04DD
04CC
04DA
04F9
04DD
0468
041D
0496
056E
0520
0285
FE65
FB08
FA01
FAB7
FB62
FB24
FAA7
FAC4
FB3B
FB3B
FAB3
FA6F
FADC
FB6B
FB6D
FB07
FAD7
FAF7
FAFE
FAE3
FB1F
FBB6
FBD3
FB09
FA90
FC4C
0056
0459
05FD
0560
048D
04CB
056E
055C
04C7
04A9
052B
056E
0506
0499
04CC
0536
051F
04B5
04BF
0537
0533
046E
03F9
04B8
05A4
048E
00DA
FC92
FA45
FA60
FB3D
FB6B
FB05
FAD8
FB07
FB28
FB1A
FB26
FB4E
FB2E
FAB7
FA7C
FAE3
FB70
FB63
FADE
FAC8
FB71
FBF4
FB71
FA87
FB02
FDDE
01F4
0507
05E7
054A
04AA
04B6
050D
051E
04DF
04AC
04BD
04F7
052A
053E
0528
04E7
04A5
04A6
04ED
050B
04A9
042A
045C
0544
0584
038A
FF7C
FB84
F9D5
FA81
FBAB
FBC5
FB09
FAA3
FAFA
FB69
FB58
FAFC
FACD
FACE
FAC1
FABD
FB0D
FB87
FBA2
FB4D
FB2C
FB93
FBD5
FB3A
FA7B
FB71
FEE4
0336
05D6
05E4
04D0
0465
04DA
0536
04FA
04AE
04D5
052D
0533
04FB
04F9
0532
0535
04DA
0495
04B9
04E6
04A3
0442
0485
053A
04E4
024D
FE3D
FAFB
FA08
FAB9
FB58
FB26
FAC3
FADE
FB38
FB38
FAF1
FAF3
FB4C
FB69
FB05
FAAB
FAE5
FB5B
FB52
FAD9
FAC4
FB56
FBB2
FB2F
FAD1
FC70
004A
043F
05FA
056F
0487
04A2
0548
0567
0500
04E4
0547
0571
04F8
0471
0485
04ED
0500
04CF
04F6
056D
055F
0485
03E7
0484
0581
04B2
0139
FCE3
FA5B
FA5D
FB5A
FBA1
FB1A
FAB2
FACC
FAF6
FAD9
FABE
FAF3
FB3B
FB3A
FB11
FB19
FB3B
FB0F
FAA5
FAA9
FB60
FC04
FBAD
FAC6
FB0D
FDAC
01AC
04BF
058F
04E3
0465
04C2
0554
0560
0500
04C4
04D4
04E9
04DF
04E3
0504
0502
04C2
04A6
04FA
055A
051F
0473
044E
0507
055D
039C
FFCD
FC08
FA60
FAC7
FB83
FB5F
FAC3
FA9D
FAFF
FB4D
FB4B
FB49
FB63
FB46
FAD7
FA9C
FAF9
FB7C
FB6E
FAF1
FAE7
FB87
FBDB
FB24
FA5F
FB77
FEF5
030C
0566
057B
04B4
0483
04F7
0548
0523
04E0
04C1
04A2
0469
0459
04A8
0512
052A
04F1
04D4
04FF
0517
04CB
046F
0497
0510
04A6
0257
FEA3
FB59
F9FB
FA6D
FB54
FB94
FB37
FAED
FB06
FB3F
FB4F
FB49
FB55
FB65
FB58
FB43
FB43
FB3B
FB02
FAC7
FAF5
FB7E
FBB2
FB3B
FB10
FCB1
0046
0401
05D5
058C
04B2
0490
04EC
04E8
0476
0453
04C1
0526
0500
049C
0483
049D
048B
046F
04C3
055A
0558
047D
03D6
0466
0558
047C
00ED
FC85
FA08
FA3F
FB7E
FBF5
FB8D
FB48
FB80
FB9A
FB38
FADC
FB11
FB8E
FBA4
FB4F
FB26
FB63
FB8C
FB45
FAF5
FB27
FB95
FB7F
FB00
FB73
FDFA
01E6
0515
0603
0528
0428
040C
0496
050A
051D
04F2
04AD
045B
042E
0462
04D3
0509
04CD
0482
0499
04E9
04E7
0489
046D
04D5
04D2
030E
FF81
FBEC
FA3C
FAA3
FBA3
FBD5
FB3F
FAC5
FAE1
FB43
FB87
FBB1
FBD9
FBD2
FB7B
FB1B
FB13
FB40
FB2A
FAD3
FAD7
FB77
FBF2
FB81
FACC
FBA6
FEF6
0342
05F7
0608
04C9
0423
0486
04FF
04D6
0462
043E
046A
0481
0477
0490
04D1
04EC
04D7
04EB
053D
0543
04A5
0406
0460
0561
0539
027E
FE12
FA90
F9AF
FABB
FBC1
FBC4
FB53
FB42
FB89
FB9E
FB60
FB2E
FB3D
FB59
FB4C
FB33
FB36
FB36
FB0F
FAFF
FB50
FBB7
FB88
FAC8
FAB8
FCAF
0073
0413
05BF
0578
04B2
0488
04C5
04B8
0466
0462
04CA
050D
04CA
0468
0478
04E0
050E
04DF
04CD
050F
052D
04C9
0469
04BF
0540
0446
0111
FD0D
FA82
FA34
FAEF
FB4E
FB38
FB49
FB88
FB70
FB09
FAFF
FB7E
FBC2
FB4A
FABA
FAE7
FB7D
FB71
FAB4
FA72
FB3B
FBE9
FB37
FA03
FABC
FE48
029F
0510
052D
049C
049F
04E9
04D8
04A6
04D6
0526
04F6
0473
0466
04EE
0539
04E0
049A
0507
0583
0520
044D
044A
050B
04B7
01EE
FDD6
FB07
FA96
FB33
FB43
FACC
FAC3
FB47
FB9A
FB62
FB12
FB0C
FB22
FB19
FB15
FB35
FB3A
FAFA
FADD
FB48
FBBC
FB66
FABC
FB89
FEBF
02E0
0568
058D
04BD
0492
051A
0562
050A
0499
048D
04C3
04E5
04E8
04D4
04A1
047E
04C6
054C
0556
04B5
045D
050E
05C6
047B
00A6
FC51
FA13
FA4E
FB30
FB2F
FA9E
FA8B
FB17
FB94
FBA3
FB77
FB3E
FB09
FB11
FB79
FBD0
FB79
FAA6
FA57
FAEE
FB6B
FADB
FA3E
FBC7
FFF0
0453
0642
05AD
04AF
04B8
0553
057D
0527
04DD
04C2
0493
0468
0498
04F3
04E3
0472
0465
04F6
055C
0519
04E9
056C
058C
0376
FF32
FB37
F9CB
FA91
FB66
FB2C
FAB1
FADE
FB4C
FB35
FAD1
FAD7
FB3E
FB67
FB3B
FB2E
FB5C
FB59
FB13
FB05
FB49
FB27
FA62
FA5B
FCD2
0152
0517
0613
0528
0494
050F
0585
0532
04B3
04CD
053C
0545
04E4
04B4
04E0
04FD
04E6
04F0
0512
04CE
0444
046A
055B
055F
02C4
FE5B
FAF4
FA41
FB24
FB80
FAE4
FA7E
FAF6
FB83
FB57
FADB
FAC8
FB03
FB09
FAF0
FB12
FB33
FAE2
FA70
FAAA
FB76
FBC3
FB44
FB77
FDF3
0202
0505
0583
04B1
0480
0520
0570
0505
04A3
04CD
0510
04F0
04B4
04D8
0530
0539
04F6
04E0
0506
0502
04E1
051F
0564
043D
00F6
FD0F
FAD5
FAD3
FB84
FB7A
FAED
FAD2
FB3B
FB61
FB00
FAB3
FAE9
FB40
FB48
FB2A
FB21
FAFB
FAAB
FAB7
FB54
FBB0
FB0B
FA51
FB85
FF3C
037A
05B4
058E
04CA
04BD
0503
04D2
0473
0493
0505
0524
04F5
04F6
0521
04FB
0495
049A
052A
056E
04E8
0477
0511
05BC
043F
002F
FC00
FA42
FAB6
FB3A
FAD4
FA75
FAF5
FBB3
FBB3
FB22
FAE6
FB28
FB42
FAFF
FAED
FB3F
FB5B
FAFD
FAD8
FB51
FB8F
FADE
FA69
FC2F
0045
0441
05D9
0554
04AE
04EC
054E
0511
04A7
04B5
04F2
04D0
048E
04B6
0512
0509
04B8
04C0
0522
0529
04B2
04A0
0553
0566
0315
FED3
FB4D
FA5A
FB0F
FB6B
FAF9
FABA
FB1F
FB7A
FB4D
FB08
FB2F
FB77
FB63
FB1D
FB23
FB50
FB22
FACB
FB04
FB99
FB67
FA5F
FA78
FD63
01F5
052B
0598
04B0
047D
0524
056B
04ED
048C
04CB
0502
04A3
043A
046E
04E1
04E7
04B5
04E2
0534
04FD
047A
04AE
0588
052F
0224
FD9A
FA88
FA52
FB6F
FBC0
FB12
FA99
FACE
FB1A
FB1B
FB1F
FB5B
FB80
FB60
FB4E
FB7F
FB8C
FB25
FAD1
FB36
FBCD
FB74
FA7F
FB02
FE3E
02A5
056B
05A7
04D9
0498
04E8
0508
04E4
04F7
0536
051C
04AA
0488
04E4
0515
04BC
0475
04BF
050E
04BC
044F
04A2
0524
040C
00B7
FCE8
FAEA
FAF9
FB66
FB14
FAA5
FAED
FB7D
FB81
FB20
FB17
FB5E
FB50
FAE6
FAD3
FB4A
FB9A
FB46
FAE0
FB12
FB63
FAFE
FA8F
FC03
FFDE
03F7
05BE
0525
0440
0473
052C
0556
04EE
04A5
04A8
049A
0474
049D
050E
0530
04CC
0476
0493
04BD
049E
04BA
056A
05A1
03C4
FFD8
FBFD
FA42
FA91
FB40
FB4A
FB16
FB3C
FB7A
FB63
FB34
FB55
FB8B
FB62
FB07
FAFC
FB3C
FB4E
FB2A
FB44
FBA0
FB82
FAB5
FA8A
FC9F
00A2
0437
0588
051E
04AE
04DE
050F
04D6
048F
048F
049A
0476
046E
04C6
051F
04F9
0499
04AC
051B
0513
0481
0469
0526
0534
02DC
FEB4
FB58
FA82
FB4E
FBC7
FB57
FAF2
FB39
FB98
FB6F
FB18
FB2F
FB87
FB8F
FB50
FB41
FB65
FB53
FB0D
FB02
FB34
FB15
FAA6
FB28
FDD2
01E8
050C
05BD
04DA
043F
0486
04E4
04B9
045D
0458
049F
04D4
04D8
04CB
04B4
048B
0473
0491
04B6
04A0
0493
050A
0591
04B0
019C
FD90
FACB
FA4D
FB13
FB8F
FB4F
FAEF
FAF9
FB4C
FB89
FB8E
FB65
FB21
FAFD
FB30
FB86
FB83
FB30
FB31
FBBA
FBF8
FB3E
FA76
FB88
FF05
031C
0564
0558
0483
0458
04C1
04FF
04F2
04FD
051D
0503
04BF
04B9
04F4
0504
04BE
0481
048A
048D
044F
0444
04DC
0545
03DE
004C
FC66
FA61
FA86
FB58
FB98
FB63
FB57
FB7D
FB6C
FB16
FAD7
FADC
FAF4
FB00
FB1C
FB3D
FB33
FB26
FB84
FC1F
FC0E
FB11
FA8B
FC44
0026
0402
05C3
0573
04B7
04AC
0502
0502
04A8
0464
0463
0494
04EC
0540
052F
04B6
0471
04C9
052F
04D0
03F7
03E0
04D8
053A
0328
FF16
FB93
FA72
FAFB
FB69
FB30
FB00
FB33
FB5E
FB43
FB3D
FB77
FB7C
FB02
FA99
FAE9
FB92
FBA1
FB15
FAF0
FB88
FBD9
FB49
FB29
FD49
015B
04EA
0610
0553
048A
0490
04D4
04C4
0499
049F
049F
0474
0480
04FD
055F
051F
0497
047D
04C1
04C1
047D
04A5
052F
04B5
01FC
FDE7
FADC
FA23
FABC
FB0B
FAD2
FACE
FB31
FB74
FB64
FB62
FB9E
FBB9
FB75
FB23
FB1D
FB33
FB19
FB13
FB7C
FBD4
FB49
FA64
FB1E
FE7C
02DA
0590
05CF
0513
04E4
0538
0544
04F6
04D8
04F0
04BB
0437
040C
046C
04A9
0461
0437
04B4
0531
04D6
0427
0460
0541
04B6
0160
FCC5
F9E6
F9EB
FB22
FB7C
FAE3
FA88
FADE
FB47
FB56
FB4A
FB69
FB94
FBAF
FBD8
FC02
FBDC
FB5F
FB1C
FB70
FBBF
FB4A
FAB8
FBDA
FF60
038D
05FA
060F
052C
04AD
04BA
04DC
04EF
0505
04F6
0499
0434
042C
045F
044A
03F8
03FF
0478
04B3
0469
045F
0514
056A
03A8
FFCB
FBEE
FA15
FA2E
FABF
FAEB
FB08
FB68
FBA1
FB5C
FB09
FB22
FB65
FB6D
FB78
FBE2
FC44
FBF6
FB43
FB29
FBC9
FBF6
FB06
FA6B
FC4C
0096
049D
061D
059B
051E
0567
0598
0514
0473
0470
04CD
04DE
0494
046A
047E
0479
044A
0450
0492
049C
0465
0491
052E
04E8
0272
FE7B
FB44
FA34
FA8D
FAC5
FA76
FA5F
FAE0
FB67
FB6A
FB2E
FB2C
FB51
FB63
FB84
FBCF
FBE0
FB6F
FAFF
FB3D
FBD2
FBB9
FAFC
FB49
FE0C
024C
0566
05F3
0520
04CC
0545
058F
0536
04C9
04C4
04E7
04D3
04A4
0499
0499
0472
0452
047E
04BA
0497
0453
0495
050D
0436
012F
FD46
FACB
FA8D
FB3E
FB5C
FAE0
FAB4
FB13
FB52
FB09
FAB3
FAD9
FB4F
FB9A
FBA7
FBA7
FB91
FB57
FB43
FB8D
FBC7
FB6E
FB05
FC03
FF16
02EF
0559
058D
04C2
0477
04D2
0512
04EC
04C6
04DD
04F1
04CE
0498
0477
045B
0445
046A
04CD
04F1
0483
040E
045E
0500
0435
0102
FCC4
FA08
F9DD
FAFC
FB97
FB53
FB09
FB37
FB69
FB30
FAD8
FAE7
FB4D
FB96
FBA2
FBA2
FB9A
FB5C
FB14
FB33
FBB1
FBC9
FB04
FA50
FB68
FEDE
0317
05B8
05EA
04E0
0446
0493
051A
053C
050E
04F0
04F3
04E0
04A6
0471
0462
0472
049C
04E9
0531
051A
0494
042C
047C
0527
04CF
026A
FE9C
FB5E
FA28
FAA2
FB55
FB53
FAEE
FAD2
FB0D
FB29
FAFC
FADC
FB10
FB6B
FB96
FB80
FB52
FB1E
FAE7
FAE3
FB4C
FBD9
FBD4
FB18
FAB6
FC20
FF7E
0336
0566
05AB
052A
0505
0537
0520
04B4
048B
04F1
0565
054E
04C9
0478
049A
04D6
04E2
04E7
050B
050A
04A9
045F
04D4
059C
0511
0218
FDC9
FAA6
FA07
FADF
FB55
FAF1
FAA6
FB0C
FB82
FB49
FAB5
FAA2
FB1C
FB61
FB23
FAFC
FB54
FB9E
FB3C
FAA6
FAD0
FB84
FB7A
FA67
FA14
FC83
0129
0514
0619
0507
0438
04A8
0554
0533
04A3
0494
0510
055C
052C
04F8
050D
0510
04B9
0473
04B8
0520
04E8
043E
043E
0542
05D6
041B
0025
FC39
FA80
FAE4
FBA3
FB8C
FB0D
FB07
FB6C
FB7B
FAFF
FA91
FAAB
FB01
FB0C
FAE0
FAF2
FB4B
FB6F
FB36
FB25
FB94
FBE4
FB50
FA6D
FB0E
FE26
024F
0508
0557
048D
0458
04D4
0503
04A0
0479
0505
058F
054F
04AF
04A6
0538
056A
04D4
044E
04A5
0543
0508
042B
041B
0537
05A7
0368
FF09
FB5F
FA68
FB5B
FC11
FBA7
FAF9
FAE2
FB15
FAEC
FA8B
FA8C
FAF2
FB25
FAF6
FAE1
FB2D
FB65
FB1C
FAB9
FAF8
FBA7
FBAF
FAB9
FA31
FBEE
FFE0
03C8
0575
04F5
041A
043C
0500
055D
0521
04F5
053D
0588
0556
04DE
04B5
04F1
0526
051C
0514
052D
0519
04AE
0478
0502
05A4
04BA
0187
FD80
FB00
FAD0
FB83
FB78
FAB1
FA53
FAC1
FB2B
FAEC
FA86
FABD
FB5C
FB79
FAE2
FA68
FAA3
FB15
FB0A
FABB
FAE3
FB6C
FB6D
FABC
FAC4
FCFF
00E9
043E
0565
0501
04C3
0547
05C2
0589
0504
04E3
0511
04FB
04A3
04A5
0534
05AB
0578
04F2
04DC
0532
0537
04B4
0476
050F
058C
0433
00A7
FCB4
FA8A
FA86
FB2F
FB2C
FA99
FA55
FAA0
FAF6
FB03
FB0A
FB3C
FB4B
FAF1
FA86
FA94
FAFF
FB22
FACE
FA9F
FB03
FB65
FAFB
FA47
FB0B
FE40
0297
058D
05F3
04E7
0447
04B0
0558
0577
0526
04F0
04F5
04F8
04E3
04E3
0505
051C
0518
052B
055E
0561
0500
04AE
050E
05CF
0572
02BD
FE66
FACE
F9C6
FAD3
FBEF
FBCF
FAF8
FA9C
FAF5
FB3F
FAFA
FA99
FAB9
FB2B
FB44
FAD9
FA76
FA86
FACE
FAF2
FB02
FB21
FB0B
FA93
FA8A
FC51
0016
03FC
05C2
0530
042C
044F
052E
056C
04D7
047F
04F9
0586
0549
04A2
0495
0535
0595
0538
04CB
04F8
0551
0518
0495
04B5
0545
04A1
01AF
FD9F
FAE7
FA95
FB6D
FBBA
FB44
FAF1
FB1F
FB3D
FAEC
FA9D
FAC8
FB21
FB13
FABB
FABA
FB2B
FB64
FB09
FABA
FB2B
FBE7
FBCB
FACB
FA95
FCC7
00DB
046E
05AC
04FD
042E
0450
04F5
0540
051A
0503
0531
0556
0538
0502
04ED
04E5
04C2
04A7
04C1
04D6
0482
03FE
0422
0530
05E3
0473
00AE
FC9D
FA8B
FAC4
FB99
FB99
FAFD
FACC
FB2F
FB5B
FAEA
FA7A
FAB3
FB42
FB5B
FAE7
FA9E
FAF1
FB7B
FBB6
FBB9
FBCA
FBA4
FAE1
FA28
FB10
FE4B
0259
04D7
04FA
0438
0449
052F
05AC
0533
048B
0488
04EC
0501
04CD
04EC
056E
0597
04F9
0432
0414
047B
04A4
0480
04D5
05B9
05BA
0356
FF1D
FB8C
FA74
FB2A
FBAF
FB32
FA99
FAD0
FB70
FB84
FB08
FACA
FB1C
FB63
FB1E
FAB7
FAD3
FB4B
FB71
FB2F
FB23
FB7C
FB7D
FAB7
FA3D
FBC4
FF6C
033A
051E
0515
04BB
0508
055A
04D6
03EF
03E5
04F9
0601
05E6
04EF
043A
0449
04A4
04C8
04CC
04EF
050D
04EC
04DB
0551
05D9
0506
0200
FDE4
FAF0
FA52
FB22
FBB6
FB80
FB30
FB4E
FB74
FB1B
FA9C
FAB5
FB63
FBD0
FB84
FB0C
FB17
FB71
FB68
FAF1
FABE
FB05
FB0F
FA6F
FA44
FC3F
0059
044F
05E0
051F
03FE
03E4
0483
04EE
0506
0538
0572
052F
047A
0418
0472
04EC
04D4
0472
048F
0522
054E
04CF
0497
055A
0605
049F
00CC
FCAE
FABF
FB3A
FC3F
FC39
FB5D
FAC3
FACB
FAFC
FB02
FB20
FB7E
FBBA
FB79
FB0E
FB14
FB84
FBB5
FB5D
FB00
FB17
FB43
FADA
FA3D
FAEC
FDD6
01E6
04D4
0562
047C
03E5
0447
04EC
0510
04D5
04BF
04D9
04CD
0493
0486
04C1
04E2
04A8
046A
0491
04E0
04C7
0466
048A
0552
056A
0357
FF71
FBEA
FA92
FB17
FBBF
FB8B
FAFE
FAEE
FB4C
FB7C
FB5C
FB51
FB81
FB98
FB64
FB2F
FB3F
FB63
FB51
FB3E
FB8E
FBFE
FBBA
FAB3
FA4C
FC17
FFDF
0385
051D
04C2
0416
043D
04D9
0503
04A7
0477
04C6
0519
04E7
0460
0422
045E
04B9
04E9
0501
050E
04D2
043F
03EC
047A
0552
04B7
01A3
FD5C
FA82
FA5F
FBAF
FC56
FBC0
FB09
FB22
FBA1
FBAA
FB43
FB15
FB45
FB4A
FB01
FB04
FB96
FBF7
FB73
FAA0
FAAD
FB90
FBE2
FB07
FA9F
FCCF
0150
053F
0643
0502
03E6
0421
04D3
04E3
047D
0466
04A5
04AB
046B
047B
04FC
0543
04DF
0459
0468
04C7
04B2
0445
047D
058D
05EE
03F2
FFF0
FC3A
FAAF
FAF7
FB6D
FB41
FAFA
FB2F
FB92
FB8B
FB2D
FB0D
FB55
FB8E
FB60
FB18
FB25
FB6E
FB8B
FB7C
FB9E
FBE6
FBB0
FAC3
FA2E
FB7B
FEE4
02B3
04DD
04FE
0466
0457
04C4
04EC
04AC
0494
04E3
051C
04DE
048C
04B1
0519
0516
0496
0458
04BB
0503
046A
038C
03D0
053C
05B7
0347
FEA3
FAC5
F9C9
FAEE
FBEC
FBAB
FAFA
FAE8
FB5C
FB92
FB55
FB17
FB12
FB0A
FAEE
FB0F
FB83
FBC0
FB56
FAC0
FAE8
FBCA
FC3D
FB88
FAC1
FBE4
FF79
03A8
0605
05F6
04F7
04A4
051A
0569
0516
04A1
0497
04D1
04D2
0497
048F
04DB
0519
04FA
04B2
0495
0494
047C
047D
04E7
0546
0451
014C
FD4E
FA7E
F9F5
FAC8
FB58
FB21
FAC8
FACF
FAF5
FAE6
FAE0
FB36
FB9B
FB82
FB11
FB01
FB7C
FBC2
FB51
FAC4
FAF2
FB87
FB6F
FAB0
FAFA
FDAD
01D2
04DF
0588
04E9
04C1
054C
0588
0510
04AA
04F4
056E
0551
04CB
04A5
04FA
050A
0473
03E5
041C
04BB
04D7
0469
046C
0541
05AF
0410
0060
FC87
FA78
FA67
FB07
FB33
FAE2
FAA8
FACA
FB0A
FB18
FAF0
FAC9
FACE
FAFF
FB46
FB89
FBB5
FBB7
FB8C
FB4F
FB34
FB4D
FB5A
FB03
FA72
FA9C
FC90
0033
03E8
05D6
059D
0490
0439
04D3
0572
0561
04F2
04D7
0522
0548
04F8
0486
045E
0474
047A
046E
049D
050C
0545
04F2
047D
04A1
054C
054D
036E
FFE0
FC4D
FA64
FA5E
FB15
FB62
FB20
FAE4
FB04
FB42
FB4A
FB34
FB4D
FB90
FBAA
FB7E
FB55
FB6D
FB84
FB32
FA98
FA68
FAFE
FBBB
FBB5
FAFB
FAE2
FCB8
0044
03CF
05B7
05CA
0514
049D
0492
0499
0489
0493
04CD
04F4
04C2
045C
043A
0496
0515
053A
04FF
04D8
0506
0531
04E2
044D
0436
04CC
04F2
0331
FF88
FBD9
FA32
FAC9
FBF9
FC32
FB86
FB0E
FB44
FB8A
FB43
FAC5
FACC
FB57
FBAB
FB60
FAF3
FB02
FB5B
FB53
FAD8
FAAB
FB47
FBFC
FBB9
FAAF
FA8E
FCCB
00D4
0465
05B4
050A
041D
0421
04C9
052B
0506
04DB
0503
052E
04F6
0493
048D
04E7
0507
0498
0422
045F
051E
0563
04C3
0425
04A5
05DF
05EA
035D
FF14
FB82
FA50
FAF4
FBAE
FB81
FAE4
FAB2
FB03
FB42
FB1D
FAE2
FAF6
FB39
FB38
FAE4
FAB9
FB1E
FBC2
FBF5
FB8B
FB16
FB1B
FB4F
FAFB
FA41
FA77
FCD0
00C1
0432
0581
050A
0475
04B9
054E
054B
04C0
0480
04E6
055E
054C
04EF
04EF
0551
056C
04E2
0436
0424
0498
04D2
047C
0445
04EB
05F2
05BB
032E
FF1D
FBB5
FA78
FAF8
FB98
FB62
FAC8
FAB3
FB30
FB7C
FB2A
FAB6
FAC5
FB34
FB51
FAEE
FAAE
FB18
FBBB
FBC3
FB2F
FAE5
FB5A
FBC7
FB33
FA1C
FA5E
FD23
015C
04A7
05A4
0507
046C
048F
04FC
0519
04F8
04FA
0520
0514
04BD
047C
04AD
051D
0541
04E2
046C
0464
04C1
04FF
04DA
04B4
0502
0566
04B2
0220
FE72
FB81
FA90
FB26
FBC4
FB86
FAD6
FA91
FAE6
FB4C
FB58
FB3A
FB47
FB6A
FB4D
FAF9
FADF
FB3E
FBB8
FBC0
FB52
FAF3
FB03
FB32
FB05
FABD
FB6C
FDDB
0169
0459
0563
04E7
045B
04AF
056D
0593
04F1
0454
0467
04E0
050C
04CC
04A7
04E3
0512
04BF
043B
043B
04C9
051E
04C1
0452
04B3
0588
0534
0298
FE93
FB56
FA45
FAD0
FB6E
FB54
FAF2
FAF3
FB4C
FB72
FB2F
FAE3
FAF6
FB4C
FB6F
FB31
FAE3
FAE4
FB2E
FB6F
FB83
FB9C
FBC9
FBAC
FAF4
FA30
FABD
FD79
0189
04D4
05E0
0524
0448
0453
04DE
050F
04CA
04A6
04E9
0528
04F6
0493
0490
04F5
0537
0500
04A3
0495
04BB
049B
0438
043E
0514
05EA
0534
0241
FE2E
FB16
FA35
FAFB
FBD1
FBBA
FB05
FA9A
FAD7
FB52
FB84
FB63
FB40
FB3E
FB3B
FB26
FB2B
FB5D
FB78
FB37
FAD1
FACC
FB3D
FB7C
FB05
FA6F
FB23
FDE7
01C9
04D5
05D4
053E
047D
0473
04E8
0529
04F2
049C
0491
04CF
04F7
04D1
048E
048D
04D8
051F
0520
04FA
04F1
0508
050A
04F8
0513
0538
047F
0206
FE48
FB21
FA19
FAD7
FBA5
FB78
FAE5
FAF7
FB9B
FBCE
FB29
FA81
FAB6
FB72
FBAC
FB22
FAA5
FADE
FB63
FB68
FAF4
FAD0
FB3F
FB7E
FAEC
FA49
FB31
FE44
0232
04EB
0589
04E5
0466
049F
0517
0531
04EE
04BB
04D4
0504
0505
04E5
04E8
0517
0524
04D7
0475
046F
04BF
04E5
04A7
0484
04FF
058A
04B3
01BE
FDCF
FB0D
FA86
FB46
FBA9
FB2B
FA9A
FAB7
FB3E
FB74
FB2E
FAEB
FB06
FB42
FB3C
FB05
FAF9
FB2C
FB4F
FB39
FB2A
FB6D
FBCC
FBB4
FB00
FA84
FB85
FE73
0238
04FA
05AE
04FB
0467
04BE
056B
0571
04C1
0440
048E
053A
0567
04F0
0479
0476
04AA
04B1
04A9
04E2
051B
04BD
03E2
0398
0488
05AA
04F8
01AF
FD64
FA90
FA28
FB07
FB84
FB2D
FABD
FAD0
FB34
FB64
FB40
FB0C
FAFB
FB02
FB1B
FB5E
FBC3
FBF7
FBAD
FB12
FAC9
FB3E
FC08
FC3F
FB7F
FAAA
FB54
FE40
0256
056D
0638
0557
0481
04A4
0538
0545
04B5
044D
0491
0519
053B
04E8
049B
048A
0473
0433
0422
048B
050B
04EF
0445
03FE
04B1
0575
048B
0157
FD49
FA97
FA1E
FAD6
FB47
FB10
FAE2
FB32
FB9D
FB87
FB0B
FAD5
FB31
FBAC
FBB6
FB62
FB3C
FB76
FBA7
FB70
FB1D
FB3C
FBB4
FBBF
FB02
FA73
FBA0
FEEC
02DC
0562
05CA
0525
04D7
051F
0543
04D5
0453
0464
04E2
0512
04A7
0429
0431
0499
04C0
0477
0442
048F
0504
0502
0498
048E
0536
0598
043B
00DB
FCFD
FA91
FA33
FAD9
FB39
FB0A
FAE4
FB2E
FB98
FBA8
FB5E
FB27
FB3C
FB68
FB6E
FB67
FB89
FBC1
FBB7
FB55
FAFE
FB1A
FB77
FB6D
FAC9
FA68
FB9D
FECD
02BE
0584
0627
0560
04A1
04A0
04EB
04D8
0475
0452
04A7
04FF
04ED
04A4
04A2
04E8
04F9
049B
0448
0481
04FC
04F9
046A
042F
04DF
058E
047E
0125
FD1B
FAA0
FA67
FB2E
FB71
FB07
FACC
FB32
FBB2
FBA5
FB31
FAFE
FB44
FB8D
FB6B
FB0D
FAEC
FB1D
FB48
FB34
FB22
FB59
FBA1
FB78
FADF
FAC3
FC43
FF74
0302
0537
0579
04B0
043B
0491
0514
0513
04AD
0480
04C0
04FA
04CB
047B
0491
0506
054C
0516
04CC
04DF
0513
04D6
0441
042E
04F5
0578
0411
0084
FC94
FA62
FA62
FB3D
FB91
FB47
FB21
FB6C
FBA4
FB5A
FAE1
FADB
FB4D
FB9A
FB5B
FAE9
FADD
FB39
FB6D
FB2F
FAF1
FB3F
FBD5
FBCA
FADC
FA3B
FB9C
FF4B
0384
05F9
0603
04FA
0482
04D9
0517
04B6
0447
0482
052F
0569
04E0
0443
0451
04E0
0533
0503
04BD
04BC
04C1
0478
0437
04AA
05A1
05BD
03B8
FFE8
FC36
FA61
FA7B
FB34
FB65
FB12
FAF4
FB54
FBB9
FB98
FB16
FAC9
FAF5
FB3C
FB34
FAF8
FAFD
FB58
FB94
FB5B
FB06
FB25
FB94
FB8C
FAD5
FA92
FC44
FFFA
03D9
05D2
0596
049A
044B
04B1
04F3
04B0
0462
0479
04C0
04CE
04BA
04F5
057D
05AB
050F
0429
03ED
0498
0553
0542
04A2
0474
050C
054C
03AC
000F
FC38
FA2E
FA56
FB4F
FBA1
FB31
FAE5
FB3B
FBB1
FB9F
FB25
FAF0
FB3B
FB82
FB53
FAEC
FAD6
FB17
FB3D
FB1F
FB1D
FB75
FBAC
FB25
FA3F
FA6A
FCB9
0093
040D
05AC
0594
0508
04F1
0522
04F6
0451
03D4
0412
04D6
0565
0559
0505
04F3
052C
0545
0506
04BC
04AB
049C
043E
03ED
0466
0587
05D3
03D0
FFDC
FC19
FA56
FA60
FAB6
FA83
FA59
FAED
FBE4
FC48
FBD5
FB34
FB0A
FB35
FB35
FADF
FA79
FA50
FA79
FADF
FB52
FB7F
FB3F
FAF1
FB1B
FB9C
FBA8
FB05
FAEA
FCE3
00D3
0498
061B
056B
0464
0464
0508
0532
04AE
0441
0476
04FF
054A
052F
04EA
04BD
04C4
0506
0562
058D
055B
0505
04E0
04DA
04A2
0454
0479
04FF
04B5
0274
FEBB
FB88
FA5D
FAD1
FB5A
FB30
FAD0
FADD
FB30
FB4E
FB3F
FB5B
FB9A
FB9A
FB4B
FB0B
FB13
FB28
FB0E
FAEE
FB02
FB20
FB0A
FAFB
FB62
FBF5
FBD0
FAF2
FAEB
FD48
0179
0500
0606
051D
0442
047E
0530
0563
0516
04D9
04D6
04D0
04B5
04B1
04BF
04B1
0493
04A8
04E8
04F2
04A4
0473
04BC
0516
04DD
0455
0471
0531
04FE
026C
FE49
FB13
FA51
FB24
FBA7
FB32
FA9E
FAB6
FB33
FB6F
FB58
FB43
FB40
FB25
FB0A
FB2E
FB79
FB8F
FB65
FB4C
FB68
FB67
FB25
FB13
FB8A
FBF2
FB69
FA63
FAC5
FDBD
0205
050C
05AA
0500
04AF
04F6
0510
04BC
048D
04D7
0520
04FB
04B6
04C7
04FB
04D7
0478
0471
04D5
050A
04B8
0454
045D
048D
0466
043F
04E0
05DF
0567
0249
FDD3
FAB5
FA30
FB11
FB85
FB24
FAC7
FAF9
FB53
FB5A
FB2F
FB20
FB1B
FAFF
FB03
FB5A
FBAC
FB85
FB13
FAFB
FB5C
FBA4
FB77
FB50
FBA8
FBEF
FB44
FA32
FAB3
FDE9
0262
056D
05ED
0525
04CB
0521
054F
04F0
0485
0482
04B4
04C4
04CA
04F2
050A
04D7
0497
04A8
04EB
04ED
04AD
04A1
04DC
04D0
043C
03EA
04AA
05B8
0508
01AF
FD53
FA8B
FA35
FAF4
FB3B
FAEF
FAD9
FB31
FB6E
FB3D
FAF9
FAFE
FB28
FB33
FB35
FB54
FB62
FB30
FB01
FB2C
FB7B
FB69
FB09
FB15
FBC3
FC1E
FB4F
FA44
FB23
FEB9
0322
05AD
05A6
04A6
045D
04E3
054D
0531
04F0
04E2
04E9
04E4
04F3
0515
04FB
0495
0457
0498
04F8
04E4
0482
047A
04DD
04FC
0488
0449
04F5
05A5
0469
00BE
FC96
FA60
FA7A
FB45
FB61
FAFC
FADB
FAFE
FADF
FA84
FA8C
FB24
FBA7
FB8A
FB22
FB11
FB5A
FB8A
FB7B
FB6C
FB6C
FB47
FB10
FB36
FBAE
FBA8
FAB0
F9EC
FB55
FF53
03CE
0631
05FD
04E1
0486
0504
0582
058D
055E
052E
04F1
04B6
04B8
04EA
04E7
0492
0458
048D
04D9
04BE
0469
046E
04CD
04E8
0491
0487
0540
05A9
0402
0023
FC1C
FA1B
FA36
FACD
FAC2
FA6C
FA82
FAE9
FB10
FAEA
FAEA
FB2C
FB49
FB18
FB02
FB52
FBAD
FBAC
FB7B
FB7C
FB8A
FB3B
FACA
FAEB
FBA1
FBDA
FAFF
FA5C
FC0A
003D
0485
0653
05AA
04A7
04C5
0581
05AA
0523
04BF
04E8
052B
0513
04C8
04A3
04A0
0496
049A
04C2
04D8
04AD
048B
04C7
0517
04D8
042C
0414
04FA
0582
03C1
FFB0
FBA4
F9E9
FA65
FB36
FB20
FA9D
FA98
FB07
FB34
FAE9
FAA2
FAC2
FB17
FB4D
FB60
FB5A
FB24
FAD7
FAD8
FB4C
FBAB
FB77
FB0C
FB36
FBDD
FBED
FAFA
FA70
FC3D
0050
0449
05F9
0595
04E9
04FE
0557
0547
0504
0513
054E
0530
04C1
0499
04E7
0520
04E6
049F
04CA
052B
052A
04C1
0475
0472
0467
044D
04AD
058F
05AA
037B
FF54
FB7F
F9F7
FA75
FB35
FB2C
FAC9
FABC
FAED
FAE7
FAB6
FAC3
FB18
FB4D
FB36
FB1E
FB35
FB39
FAFF
FAD5
FB07
FB4E
FB4B
FB33
FB79
FBDC
FB86
FA80
FA5D
FCAE
00E5
048E
05DE
0568
04EC
051C
0553
0505
049B
04A7
04FE
0517
04E3
04CE
04F0
04F8
04D0
04D9
0532
0563
0517
04B6
04C5
0500
04CB
045D
04A2
059A
059C
030F
FEAD
FB21
FA2B
FAE4
FB49
FABB
FA3A
FA8D
FB36
FB68
FB2C
FB14
FB3D
FB42
FB0A
FAFA
FB33
FB41
FAE2
FA87
FAB6
FB3A
FB80
FB79
FB82
FB86
FAFB
FA19
FA5C
FD0E
0167
04F3
0605
054E
04A2
04D3
054C
0563
052F
0513
050C
04E6
04AD
0497
049E
0493
048F
04D2
0533
0536
04D6
04AA
04F6
051E
04A1
0427
04C0
0602
05D9
02D9
FE40
FAE1
FA24
FADD
FB38
FAE3
FAB3
FAFC
FB30
FB03
FAF2
FB5B
FBC5
FB90
FAFE
FAE2
FB68
FBD2
FB99
FB1E
FAF5
FB0B
FB07
FB0B
FB5A
FB8C
FAF9
FA19
FAAC
FDCB
0236
054D
05D1
04F7
049A
0516
0578
052C
04A5
0479
0495
049B
048A
0498
04BE
04C2
04AE
04B6
04CA
04A5
046E
04A8
0548
057E
04DC
043D
04B8
05C1
0540
01FF
FD72
FA62
FA00
FAFC
FB7F
FB2C
FAD3
FAEC
FB25
FB3E
FB64
FBAF
FBCE
FB93
FB50
FB62
FB93
FB74
FB1F
FB1A
FB6B
FB77
FB0E
FADB
FB57
FBD1
FB5C
FA92
FB5B
FE9A
02B6
052C
0548
0493
049B
053A
056B
04FE
04A6
04BA
04C6
0475
0420
0431
0476
0478
044A
045E
04B9
04E2
04B0
0492
04C2
04CD
0469
0432
04D4
058F
0491
0128
FD05
FAA2
FAA7
FB82
FB90
FADB
FA77
FACE
FB56
FB90
FB8F
FB8E
FB87
FB72
FB7C
FBAF
FBB7
FB59
FAF2
FB0E
FB88
FBAD
FB52
FB21
FB77
FBA3
FAF8
FA4F
FB7A
FF04
0320
0571
057D
04C4
04AB
0511
052B
04E1
04B1
04B9
049D
044D
0436
0486
04DA
04D1
04A4
04BB
04F5
04DB
047B
045F
04A6
04BF
046C
045C
0510
058A
0415
0071
FC90
FAA2
FACE
FB74
FB5D
FAE0
FACE
FB23
FB4F
FB44
FB67
FBB3
FBAB
FB35
FAE7
FB31
FBA6
FB9F
FB31
FB05
FB4A
FB79
FB44
FB19
FB49
FB56
FAD4
FAA0
FC46
FFFC
03DE
05BB
055B
046D
045D
04F9
0541
04EC
0482
0476
04B1
04F4
0522
051B
04C7
0459
0442
049C
04EF
04CF
0482
0493
04EA
04EA
0489
0495
0558
0597
03B1
FFC6
FBF0
FA29
FA64
FB1C
FB49
FB29
FB3A
FB56
FB29
FAEA
FB02
FB54
FB6B
FB42
FB46
FB9B
FBCE
FB8E
FB34
FB38
FB6C
FB4F
FAFB
FB0D
FB89
FB91
FACD
FA89
FC74
0066
0423
05A4
0523
046D
04A2
0541
0568
0515
04E0
04F2
04F4
04BD
0488
047D
047B
0470
0481
04B7
04CB
048D
044D
0473
04D5
04EB
04B3
04CC
0550
0521
0305
FF5B
FC12
FABA
FB0C
FB84
FB34
FA85
FA54
FAD6
FB89
FBE1
FBAE
FB1D
FA9A
FA92
FB0F
FB9C
FBCC
FBB6
FBBB
FBD9
FBAA
FB23
FAE7
FB64
FBF5
FB8C
FA6B
FA68
FCF3
012D
0497
059B
04E9
0441
0476
0505
053A
050D
04D8
04BA
04A4
04A6
04D1
04F9
04DF
0491
045C
045C
0472
0492
04D8
0520
04F7
0442
03C2
044C
0568
054E
02BE
FE9D
FB39
FA0D
FA93
FB4E
FB7C
FB67
FB7D
FBA1
FB89
FB45
FB1F
FB28
FB35
FB3C
FB57
FB85
FB91
FB64
FB35
FB41
FB78
FB8A
FB59
FB29
FB4B
FBA8
FBCB
FB65
FADC
FB31
FD3C
00BE
043B
060E
05D4
04AE
0412
0462
04EA
04F8
04A9
047C
048A
0483
045A
046B
04DD
0543
0524
04AE
0473
049C
04C1
049A
0473
04A4
04F3
04E8
049F
04B7
0536
04F8
02CF
FF1B
FBB4
FA2C
FA65
FB18
FB5C
FB4F
FB5F
FB86
FB7C
FB4F
FB58
FBA0
FBBA
FB5F
FAE4
FACF
FB21
FB55
FB18
FACB
FAFB
FB91
FBDB
FB7C
FAFA
FB09
FB80
FB75
FAA3
FA4B
FC24
004C
04AC
06D0
0645
04C8
0438
04C8
055A
0538
04C1
048C
0480
0439
03E2
041E
0503
05CD
05CA
053F
04F6
0522
0535
04D6
0476
049D
0508
0502
048B
0478
051B
054E
037A
FF96
FB98
F9A0
F9F0
FB06
FB72
FB25
FAE7
FB0B
FB31
FB10
FAF5
FB38
FBA0
FB9E
FB1D
FAA4
FAA5
FAE9
FAF0
FAB5
FAB2
FB21
FB8F
FB7D
FB1F
FB1D
FB95
FBD5
FB6B
FB28
FC89
FFE6
03AB
05C5
05AE
04C2
0487
051E
0595
055C
04E0
04BD
04E8
04F4
04D4
04DE
0525
0546
04FF
04A8
04B7
0509
0517
04CE
04BE
052F
0583
04F9
03F3
03BD
04CC
05A2
042A
002D
FBE4
F9D1
FA4B
FB8B
FBDD
FB3D
FAB5
FAC0
FAE6
FAB9
FA86
FAC4
FB46
FB6F
FB19
FACC
FAF6
FB4D
FB44
FAE9
FACB
FB1D
FB5F
FB23
FAC8
FAFC
FB9B
FBB0
FADC
FA55
FBE0
FFB3
03DD
060F
05D6
04BC
0460
04E1
054D
0523
04DE
0512
0589
059C
0525
04B1
04BB
0519
054F
053F
0528
0521
04EF
0486
0456
04BF
0569
0590
0516
04C8
053B
0594
0429
0074
FC21
F99A
F9AB
FAF0
FB9A
FB43
FACF
FAE7
FB3D
FB3F
FAF5
FACC
FAE3
FAF1
FAD8
FAD2
FAF1
FAE3
FA86
FA52
FACD
FB9E
FBC6
FAF8
FA2E
FA79
FB7F
FBCB
FACC
F9FD
FB6B
FF50
03A1
0610
0634
056A
050F
053F
054D
04EA
0470
0445
045B
0477
0498
04E7
0556
0596
057A
053C
053A
0576
0591
0550
04F8
04E6
0508
04EF
0496
0497
054C
05D2
048A
00E9
FC8C
F9E8
F9E2
FB16
FB9A
FB0B
FA80
FACA
FB77
FBAB
FB52
FB09
FB1B
FB30
FB0B
FAEB
FAFE
FAE8
FA59
F9CD
FA1C
FB33
FBF2
FB8D
FAAD
FA8D
FB3A
FB74
FA94
F9E4
FB5E
FF3D
036F
05A6
058D
04A9
0472
04FF
0583
0585
0540
050E
04F3
04C6
048A
046C
0481
04B3
04EA
052A
0577
05AE
059D
0549
0501
0508
0533
0522
04D5
04D3
056A
05D5
049B
0127
FCE2
FA25
F9F8
FB27
FBC9
FB4C
FAA1
FA9D
FAF1
FAEA
FAA5
FAD9
FB9E
FC22
FBC5
FAFF
FAB0
FAEE
FB0C
FABD
FA7F
FABD
FB10
FADB
FA5B
FA74
FB4C
FBD7
FB3B
FA4B
FAF7
FE1E
026A
0592
067A
05D9
0512
04CE
04D9
04E1
04E5
04FC
0510
04FB
04BF
048A
0483
04AC
04F0
053E
057A
0577
051B
0493
0450
0493
0518
054C
0502
04C1
0518
0597
04DB
01F2
FDC1
FA79
F98F
FA6B
FB48
FB2F
FAA6
FA99
FB12
FB63
FB37
FAF1
FB04
FB4E
FB6B
FB46
FB14
FAE7
FAA9
FA83
FAD3
FB90
FC19
FBE1
FB3B
FAF9
FB42
FB46
FA77
F9BD
FAD3
FE4C
02A0
0580
0600
0532
04B6
0515
05A0
05A0
052D
04D7
04DC
04F1
04CF
048F
047E
04AF
04F4
0522
0538
0539
050A
04AD
046D
0498
0504
0523
04BF
0465
04BB
055D
04DB
0229
FE0B
FAA4
F97C
FA2B
FB13
FB2F
FAC8
FAA3
FAE7
FB21
FB0C
FAE5
FAF8
FB34
FB61
FB7A
FB9D
FBB2
FB7F
FB11
FAD3
FB03
FB52
FB4A
FAF9
FAEC
FB64
FBD5
FB9C
FB1A
FBA9
FE35
01F9
0503
0600
0567
04B8
04D5
0550
0551
04BE
0446
0470
04FD
0554
0534
04D6
0480
0447
0433
045A
04AD
04E2
04C5
0495
04B6
050B
0500
0466
03F0
0462
0546
04F9
025B
FE44
FAE8
F9C1
FA52
FB11
FB29
FAFA
FB24
FB93
FBBC
FB76
FB29
FB34
FB75
FB8C
FB62
FB33
FB2B
FB37
FB3F
FB5C
FBA0
FBD4
FBAD
FB43
FB1C
FB7B
FBDF
FB88
FAA2
FA99
FCC9
00D9
04B3
0665
05E5
04D4
0493
0509
0543
04E1
046C
046A
04AE
04C2
0499
0486
04A3
04B7
04AD
04C3
0512
052E
04B8
0408
03E5
0471
04E4
04A5
043D
04AC
05C1
05D0
036E
FF3F
FB8D
FA12
FA72
FB10
FAF2
FA7C
FA7B
FAFD
FB6C
FB65
FB2E
FB35
FB7B
FBA4
FB7D
FB3B
FB1F
FB1E
FB09
FAEE
FB0B
FB64
FB9F
FB7A
FB3A
FB52
FBA3
FB7D
FABA
FA80
FC57
0040
0440
062E
05D9
04F3
04F2
0594
05B5
050D
0478
04A2
0520
052A
04C1
0482
04AC
04D8
04C0
04B6
0508
055D
0525
048A
0458
04D5
053A
04CA
03FF
0407
0502
0565
038D
FFB1
FBDE
F9F7
FA11
FAD0
FB12
FADB
FACA
FB14
FB5D
FB4D
FB03
FADC
FAF4
FB0F
FAFB
FADE
FAF1
FB23
FB2C
FB06
FAFE
FB3D
FB79
FB55
FB09
FB28
FBB8
FBED
FB4F
FAE9
FC80
0060
047E
0662
05C0
048D
0488
055D
0599
04DD
043C
048F
0548
0569
04FA
04DB
0554
05B1
055D
04C8
04AE
04FC
04FE
0485
043B
0492
0501
04D3
0455
047A
054B
0559
0337
FF4A
FBA2
FA05
FA5F
FB34
FB55
FAD4
FA7D
FAC0
FB4C
FB95
FB6C
FB12
FACF
FAA0
FA66
FA36
FA4E
FAB6
FB2B
FB72
FB9B
FBC7
FBD5
FB91
FB2E
FB2A
FB89
FB8D
FAC6
FA38
FBB8
FFB4
0425
0663
05E5
049D
0486
0583
060F
0581
04C4
04C9
0539
0529
04A0
0487
053A
05E9
05B7
04E5
0464
0486
04B8
0491
046D
04B4
0504
04B7
0408
03FD
04EF
059C
0450
00D4
FCE2
FA78
FA13
FAA4
FAFD
FAD9
FAA4
FAAB
FAD1
FADD
FACF
FACF
FAEC
FB10
FB22
FB29
FB33
FB43
FB51
FB64
FB85
FB9C
FB7C
FB21
FAE3
FB24
FBB6
FBD2
FB0F
FA57
FB5D
FEC2
0309
05CC
0614
051C
04B0
052C
0592
0538
04AE
04C1
0542
0561
04E7
0483
04B7
051A
04FF
0474
0432
048B
0504
0510
04D1
04C1
04E5
04DE
04A9
04CC
0567
058B
03F6
0092
FCDD
FA9C
FA45
FAD7
FB2B
FB0D
FAFD
FB3F
FB81
FB64
FB0E
FAEC
FB23
FB66
FB68
FB37
FB1A
FB24
FB2F
FB23
FB16
FB18
FB12
FAF9
FAFF
FB49
FB97
FB69
FAC2
FA88
FBEA
FF26
0304
05B2
0638
0531
0418
03F4
049C
0531
051D
0499
0443
046B
04DD
053C
055E
0545
04FF
04AD
0489
04A8
04DE
04F2
04F1
050C
0529
04E4
043B
03EE
04A2
05A2
051A
020A
FDAB
FA68
F990
FA55
FB22
FB57
FB67
FBB2
FBE3
FB9C
FB22
FAFE
FB3A
FB63
FB3C
FB08
FB1C
FB61
FB76
FB2A
FAB7
FA82
FABE
FB3A
FB8E
FB72
FB11
FAEA
FB3B
FB99
FB61
FABE
FAE7
FCF7
0095
0409
05C2
05A7
04D9
0461
0465
047F
0479
0473
0490
04BF
04E0
04ED
04EE
04EA
04E9
04F7
050F
051D
051F
052D
054B
054A
0501
04A0
0485
04B3
04BF
0478
045F
04FF
05C4
050F
01EB
FD8A
FA77
FA1A
FB6E
FC58
FBEF
FB07
FABB
FB17
FB5A
FB22
FAD4
FAF1
FB64
FBAE
FB77
FADC
FA48
FA2A
FA9D
FB39
FB6B
FB23
FAE6
FB18
FB66
FB44
FAD1
FAC1
FB47
FB9F
FB36
FAF1
FC78
0012
03DB
05AF
055C
047B
0464
04F3
054F
0530
04F2
04D7
04C6
04B6
04D6
0521
0541
0512
04E6
0507
0539
0527
04F5
0507
054B
054C
04EE
04AC
04D3
04FE
04B7
0460
04B5
055F
04C0
01D3
FDB6
FAC2
FA27
FB00
FBB3
FB9F
FB44
FB26
FB35
FB25
FAF5
FAD8
FAE9
FB26
FB7A
FBA2
FB4F
FAA1
FA35
FA75
FAFF
FB1B
FABD
FA97
FB0A
FB88
FB65
FAEB
FAFB
FBA2
FBDC
FB26
FAB8
FC5D
0024
03F8
05C1
0569
0481
0440
0486
04B3
04B6
04E2
052E
0535
04E0
0492
049C
04E0
0514
052D
0544
054E
0533
050B
0501
0504
04DB
04A1
04B2
0503
04FA
0455
03D4
045A
055E
04FC
0205
FDB5
FAA9
FA3A
FB51
FC05
FBB3
FB22
FB10
FB5B
FB84
FB67
FB36
FB17
FB06
FB02
FB02
FADF
FA96
FA7A
FADD
FB79
FBA6
FB47
FB00
FB41
FB90
FB45
FAB5
FAD3
FBA9
FC0D
FB4D
FAA7
FC24
FFF6
03E1
0595
051A
0441
0444
04BB
04D2
0495
04A0
0513
0569
0544
04E0
049F
0498
04B8
04FD
0548
0549
04E8
048F
04A5
04F2
04F1
04A5
049F
050F
0556
04F4
0476
04CD
05A1
052E
0249
FE11
FAFD
FA51
FB1F
FBBA
FB8F
FB33
FB2D
FB51
FB42
FB0F
FAF6
FAFB
FAFB
FAFA
FB0C
FB14
FAF4
FAD4
FAF7
FB3B
FB2F
FABF
FA75
FAC2
FB4A
FB60
FB06
FAE7
FB34
FB33
FA84
FA41
FC0F
FFF8
03E5
05B1
0557
0493
04A5
0527
052A
04B6
048C
04F4
0566
056A
0526
04FB
04F0
04D9
04C4
04E0
051C
052E
0509
04F1
04FF
04FE
04E2
04F9
055A
0587
0515
0481
049F
052F
04A3
01E0
FDEA
FB15
FA87
FB30
FB67
FAE3
FA8A
FAD2
FB2A
FAFD
FA90
FA88
FAF6
FB61
FB7E
FB70
FB51
FB01
FA98
FA87
FAF9
FB72
FB68
FAFF
FAC6
FADD
FAE7
FAC7
FAD9
FB30
FB31
FA95
FA76
FC7A
0099
048E
060F
0537
041B
0439
0515
0571
0519
04D4
050D
054E
0526
04DA
04DB
050D
050E
04E1
04DC
050B
0521
0507
0503
0539
0561
053D
0509
0512
0521
04D9
0486
04DA
0583
04E3
01DF
FDA2
FAB3
FA4B
FB36
FB91
FB00
FA91
FAE9
FB6D
FB5F
FAF0
FABD
FAD1
FAD0
FAC2
FAFE
FB6D
FB7D
FAFA
FA77
FA85
FAE3
FAF0
FAA6
FA93
FAEC
FB3D
FB47
FB63
FBBE
FBBD
FB01
FA99
FC37
FFFC
03D0
057A
04F6
0424
0458
051D
056B
053B
0538
057F
0589
0523
04CA
04DE
0517
050D
04E1
04FA
0545
0546
04E3
0497
04BE
050A
0513
04ED
04DA
04C1
0478
0460
04F3
059F
04CE
01A5
FD79
FABD
FA7E
FB7A
FBE1
FB60
FAE0
FAE6
FB05
FAD0
FA96
FAC9
FB31
FB46
FB02
FAE8
FB23
FB40
FAF9
FAB0
FADB
FB46
FB67
FB34
FB17
FB37
FB4D
FB3E
FB5B
FBAD
FB91
FAB7
FA40
FBF4
FFF6
040B
05D4
0546
0451
0465
051A
0560
051B
04F3
051E
0522
04D1
04B2
0510
0563
0517
047D
0453
04B1
04FC
04E1
04B8
04D5
0508
0506
04EC
04F3
04E2
0476
042F
04CF
05D0
054B
021D
FDAC
FAA7
FA34
FB14
FB8E
FB5D
FB47
FB86
FB84
FB08
FAB2
FAF5
FB59
FB3E
FAD2
FAB2
FAEB
FB05
FAEE
FB11
FB8A
FBCD
FB79
FB02
FB0A
FB6B
FB77
FB1D
FB10
FB7D
FB8D
FAC4
FA56
FC0C
FFF1
03DE
05AA
054E
0472
044F
04B2
04ED
04ED
0502
0524
050B
04C6
04B8
04F7
0528
050B
04D4
04C8
04D7
04CA
04AE
04B9
04DE
04D1
0491
0479
04A5
04B0
0464
044D
04FE
05D6
0527
0219
FDF9
FB1E
FA8D
FB38
FB99
FB5E
FB26
FB2C
FB05
FA8D
FA56
FAD2
FB8E
FBB6
FB3B
FAD1
FAE2
FB12
FAFB
FADB
FB11
FB6D
FB78
FB35
FB16
FB37
FB42
FB21
FB4A
FBDE
FC1C
FB62
FAA9
FBE1
FF8C
03A9
05C2
0589
04AF
0491
04EC
04F1
04A9
04B2
0514
0532
04D8
0495
04C9
0518
0512
04EC
0501
051D
04E4
0494
04B6
052D
0549
04D6
047D
04B4
04EA
0471
03D7
043F
0548
04D5
01A7
FD56
FABD
FABB
FBA2
FBB3
FB14
FAF1
FB7A
FBC7
FB63
FAF1
FB07
FB43
FB07
FA8C
FA82
FAF6
FB4E
FB40
FB21
FB33
FB3C
FB09
FAE6
FB20
FB6D
FB53
FB0C
FB4E
FC0E
FC3D
FB59
FAB4
FC3E
0018
0408
05C0
052B
0417
03F8
049C
050F
0504
04EC
0519
0555
0554
051C
04DC
04AF
04AB
04E6
0539
0539
04B8
042F
043E
04D6
0542
0523
04E7
04F6
04F1
0455
039F
03E1
04FE
050D
026A
FE0C
FAD6
FA6B
FB8A
FBF9
FB3E
FA9A
FADB
FB60
FB5A
FB08
FB1B
FB72
FB58
FAC9
FA94
FB10
FB86
FB53
FADF
FAD8
FB18
FB12
FAE1
FB18
FB9A
FB97
FADF
FA6F
FB0A
FBE5
FBCD
FB51
FC7F
0009
03DC
0579
04E6
042C
0486
0535
0527
0494
045C
0499
04AD
0472
0476
04E3
0527
04F3
04D7
0539
0586
051D
0470
0465
04E7
0511
04B0
04A8
056B
05FD
0547
03F9
03CD
04DA
04E9
022C
FDC8
FAA0
FA13
FAF1
FB79
FB4B
FB0D
FB11
FB1F
FB2F
FB85
FC05
FC19
FB92
FB17
FB3D
FBA4
FB89
FAEE
FA93
FAD6
FB40
FB49
FB14
FB05
FB13
FAF3
FACF
FB1E
FBC0
FBD1
FAFE
FA85
FC2F
0017
042A
0621
05B5
0489
042A
04A7
0527
0536
050D
04EF
04CA
048C
046F
04A3
04FA
051B
04EB
049C
045D
0446
0481
0519
05A6
0592
04EA
0473
04A8
0503
04C4
0433
0451
051D
04F0
0247
FDF1
FA93
F9CE
FABC
FB76
FB57
FB0C
FB10
FB19
FAEE
FADE
FB1D
FB3D
FAD5
FA54
FA7F
FB45
FBBE
FB78
FB0F
FB1F
FB56
FB21
FAB7
FABB
FB29
FB5E
FB2A
FB16
FB6E
FBB1
FB7C
FB90
FD2F
005F
038F
0545
0588
0547
0503
04B0
046B
048A
0502
0562
0577
057E
0598
057D
0500
048D
04A2
0501
04F9
0481
045D
04E7
0568
0530
04B5
04D8
0571
056F
0477
039C
03F5
04F4
04BD
023F
FE71
FB4D
F9F2
FA06
FA85
FABB
FA99
FA87
FADE
FB7D
FBD2
FB8A
FAF3
FA9B
FAA9
FAD9
FAF7
FB11
FB2E
FB1B
FAC3
FA87
FADB
FB97
FC04
FBBB
FB1F
FAD3
FAF6
FB45
FB9A
FBEC
FC00
FB99
FB1C
FB90
FDAB
00F2
03F7
0599
05CD
0554
04DF
04A9
04AA
04CD
04FB
0516
0511
04F8
04DE
04D5
04E3
04FB
050D
051D
0536
0541
0518
04BE
047A
0481
04A3
0485
0425
03F3
0441
04BC
04D0
047D
0470
04F5
0533
03D9
009D
FCCD
FA44
F9D9
FAC8
FB9D
FB90
FB06
FACA
FB0F
FB57
FB3E
FAF7
FAE9
FB0B
FAFC
FAB5
FAB8
FB56
FC0B
FC14
FB79
FB06
FB2D
FB75
FB5E
FB2E
FB63
FBC0
FBA2
FB1B
FB08
FBBC
FC42
FB98
FA73
FAE4
FDF3
0236
0534
05DE
0527
048B
04A2
0516
055D
0545
04FF
04D7
04E7
0502
04F0
04C1
04B9
04E9
0501
04C6
047D
048E
04CF
04B4
043F
0420
04A8
052C
04FF
047A
046F
04D9
04E7
0468
0444
04F7
053A
0332
FF0C
FB46
FA00
FAB7
FB5E
FB0A
FA8A
FAB0
FB26
FB34
FAF1
FAF9
FB62
FB90
FB33
FAC8
FADE
FB44
FB6C
FB3F
FB26
FB4F
FB6A
FB36
FAEF
FB06
FB8F
FC10
FBFA
FB4C
FAB2
FACB
FB65
FB9C
FB07
FA9B
FBFA
FF99
03D1
063D
061A
04E0
046A
0501
0590
055C
04E2
04E9
0560
058B
0517
0484
0471
04D4
0520
0518
0505
0527
053F
04E9
0448
03F4
043D
04BB
04D2
0484
0464
04BA
050A
04DC
0494
04E6
056C
0497
017A
FD4D
FA69
F9DF
FA92
FADB
FA73
FA47
FAD5
FB75
FB6A
FAEC
FAB4
FAEA
FB1E
FB10
FAFB
FB13
FB34
FB30
FB32
FB76
FBD8
FBE4
FB74
FAF6
FAF1
FB5E
FBAD
FB73
FAE9
FAB0
FB0F
FB8F
FB70
FACF
FB09
FD7A
01AA
054D
0678
058B
0493
04D6
05B0
05DA
0537
04C3
0502
055B
0526
04B1
04AA
0505
051C
04B7
045D
0479
04C5
04C1
0479
0471
04D9
0540
052B
04BE
0486
04B4
04E5
04C0
047C
049E
0521
0513
0351
FFD6
FC2A
FA26
FA2D
FAF6
FB20
FAA6
FA6F
FADF
FB57
FB32
FAB2
FA98
FB12
FB8E
FB9E
FB74
FB5F
FB42
FAEE
FAA6
FACB
FB32
FB4A
FAEE
FAA8
FAF3
FB87
FBB1
FB48
FAEA
FB2A
FBBC
FBCF
FB2B
FAC2
FBE8
FF03
02E5
05A2
0630
054E
0498
04D4
0560
055A
04D3
0484
04AE
04E1
04C5
04AB
04F7
055E
0541
04AB
0458
04A9
0516
0508
04BA
04CA
052F
0540
04C2
044F
047A
04FA
050E
04A3
047E
0513
0598
04A5
01BC
FDF3
FB0A
F9F9
FA59
FAFF
FB1A
FAC9
FAA4
FADD
FB10
FAF0
FABE
FAE5
FB54
FB8A
FB46
FAE4
FADF
FB2A
FB55
FB38
FB18
FB2D
FB4E
FB54
FB64
FB9D
FBB4
FB51
FABC
FAAC
FB55
FBF4
FBAE
FACC
FABE
FCBF
0073
0419
0611
0624
0562
04F9
0532
0585
056B
0501
04C5
04E2
0515
0529
0539
0558
054A
04E3
0471
046D
04CB
04F8
04A2
0434
043C
0499
04AF
0467
0461
04ED
056A
051B
045B
0445
051A
0588
03FB
006D
FC95
FA4A
F9E7
FA64
FAAA
FA89
FA78
FAC0
FB20
FB2F
FAE5
FAA8
FACC
FB22
FB39
FAFE
FAD7
FB0A
FB63
FB88
FB7A
FB75
FB78
FB51
FB0C
FB0B
FB6B
FBA9
FB45
FAA2
FAA6
FB6E
FBEC
FB57
FA8D
FB63
FE8A
029C
0573
062B
0594
04F3
04D3
04FD
0527
0543
0543
050C
04BB
04B0
051A
05A2
05AB
0504
043A
0412
04B1
0565
0575
04FA
04AA
04DA
051C
04FA
04AD
04C0
0520
051F
0487
042B
04D7
05E0
0570
0291
FE6C
FB31
F9FB
FA39
FAC7
FB1A
FB41
FB4F
FB33
FAF7
FACE
FACC
FAD5
FAD4
FAE3
FB0F
FB2B
FB13
FAF1
FB08
FB52
FB87
FB70
FB1F
FAD2
FABF
FAED
FB27
FB2C
FAFE
FAF3
FB43
FB95
FB49
FA79
FA67
FC6A
0046
040C
05E3
05BF
0509
04E6
053B
0562
052D
04F9
04FD
0507
04E9
04D0
04FD
054E
0560
0517
04C6
04C2
04FC
051B
04E7
048C
0464
0494
04E4
0512
0522
053C
054E
0518
04B3
04AF
0553
05C5
0480
00FB
FCB1
F9F9
F9C5
FADF
FB7D
FB23
FAA8
FAB8
FB03
FAF8
FAAB
FAA6
FB00
FB3E
FB15
FADD
FB03
FB59
FB57
FAF3
FABA
FB00
FB61
FB4F
FAE9
FAD4
FB44
FB92
FB1B
FA49
FA2E
FB0F
FBD3
FB5E
FA4F
FAAD
FDAB
020F
054C
060B
0541
04B6
050E
058D
0581
0529
0514
0540
0539
04F0
04D2
0517
055A
052E
04BF
049F
04F4
0541
0518
04B7
04B0
0519
056D
0543
04E0
04CF
051C
053E
04DF
0476
04BD
0580
0563
0338
FF80
FC2F
FAC9
FAFC
FB4C
FAE5
FA47
FA3A
FAA8
FAE0
FAB5
FAAE
FB15
FB67
FB1B
FA7E
FA58
FADD
FB69
FB71
FB33
FB37
FB7B
FB7E
FB1D
FADC
FB28
FBA5
FBA1
FB0E
FAA5
FAF0
FB83
FB7C
FAB4
FA43
FB95
FEE4
02B6
0515
055B
04A1
0467
0507
05A6
0591
051D
050E
0566
0576
04F7
0483
04B3
0535
054C
04E4
049B
04C6
04F9
04BF
0461
0472
04DC
04E9
0467
040B
046C
050D
0503
0468
0461
057A
0679
056E
01E7
FDA5
FAF7
FA96
FB49
FB87
FB00
FA7A
FA91
FAFC
FB1C
FADE
FACB
FB37
FBB6
FBA5
FB0A
FA92
FAAC
FB01
FB0D
FAE1
FAF9
FB70
FBC7
FBA9
FB6E
FB9A
FBFF
FBEA
FB39
FAB4
FB05
FBA6
FB8A
FAC4
FADE
FD32
0123
047C
05A7
051E
0487
04C1
0535
050C
0473
0446
04D4
057A
0587
051B
04D5
04EC
0505
04E1
04CA
050B
0550
0512
0472
0431
04A3
051E
04E3
0435
0400
0483
04EC
048B
03EC
042B
0531
0559
032C
FF35
FBA2
FA2A
FA9F
FB87
FBC0
FB58
FAFC
FB02
FB21
FB03
FACD
FAE0
FB36
FB5B
FB08
FA99
FAA2
FB23
FB74
FB29
FAB3
FACB
FB6A
FBC9
FB84
FB24
FB49
FBB3
FBB6
FB56
FB4A
FBC7
FBFC
FB49
FA99
FBB6
FF22
0328
0589
05BE
0514
04D9
0514
0517
04BA
047D
04B7
0512
0511
04BF
049D
04E6
054A
0562
0532
0511
0520
0523
04DB
046E
0442
0471
04A5
0497
047C
04AC
04F8
04CE
042C
03ED
04AE
059A
04EA
01E1
FDE0
FB2D
FAA9
FB38
FB5A
FAD5
FA84
FAE7
FB7F
FB98
FB39
FAF6
FB1C
FB5D
FB52
FB08
FAE8
FB20
FB65
FB61
FB21
FAF8
FB09
FB1A
FAFA
FADA
FB15
FB9A
FBE8
FBA9
FB35
FB1D
FB58
FB59
FB12
FB6F
FD60
008E
037F
050A
0558
0558
057C
0577
0510
04A7
04B4
050B
051D
04C2
0470
0494
0504
0533
04E3
0468
043C
0476
04C0
04CD
04B5
04BD
04E5
04F1
04D1
04CD
0512
0541
04CC
03E8
03A1
0485
056C
0455
00BD
FC94
FA4C
FA5F
FB2C
FB34
FAA7
FA8C
FB07
FB4A
FAF5
FAA3
FADD
FB39
FB0C
FA93
FAA0
FB50
FBC6
FB69
FAC9
FAD2
FB77
FBC7
FB4C
FABA
FAEA
FBA1
FBE4
FB61
FADC
FB11
FBB7
FBF4
FB94
FB36
FB4A
FB75
FB4B
FB61
FCF5
0049
03DF
05C8
05A7
04E9
04FA
05C2
061F
058D
04B6
0474
04C7
0519
0531
054B
0573
0550
04CA
0462
048C
04EC
04CE
0431
03E1
0468
054B
05A3
053E
04BB
049E
04BC
04B6
0490
0487
0495
0490
04A4
0516
057D
04B2
01FB
FE2A
FB1D
FA03
FA5D
FAD1
FAB1
FA68
FA85
FAEE
FB20
FAF5
FAC2
FAC5
FAD5
FABD
FAA1
FAD0
FB3F
FB84
FB68
FB34
FB42
FB6D
FB4C
FAE5
FABA
FB14
FB8B
FB98
FB48
FB0F
FB10
FB02
FADD
FB13
FBBE
FC0B
FB3F
FA3B
FB16
FEB2
0349
060E
0614
04EF
0487
0517
0597
057C
053E
0549
0557
0520
0508
0577
05FF
05C6
04CD
040E
0448
050E
0574
053E
04F6
0502
051D
04ED
04AC
04C6
0526
054B
050C
04D7
04FB
0526
04E2
0462
045F
04FB
051F
036E
FFE7
FC48
FA74
FAA5
FB6D
FB75
FAD5
FA89
FAF6
FB76
FB54
FABA
FA5E
FA86
FADC
FB16
FB54
FB9E
FB9D
FB20
FA99
FA9E
FB0F
FB38
FACE
FA61
FA8A
FB0B
FB2F
FADB
FAA4
FAE1
FB31
FB3C
FB55
FBD6
FC35
FB98
FA5C
FA49
FCBC
00E4
0468
05BF
0571
04F9
04FE
0520
050B
0502
0543
057A
053D
04C3
04AD
051D
0577
052A
0478
0429
048D
052A
0570
055F
054D
054B
051E
04CC
04B0
04ED
051D
04E6
048F
04A7
0519
0528
048A
0416
04AA
0598
04F6
01DB
FDBB
FAFF
FA86
FB14
FB2A
FAB2
FA8B
FB01
FB6E
FB46
FAD9
FAB8
FAE3
FAEE
FAC1
FAAB
FACB
FADD
FAB2
FA8B
FABA
FB22
FB59
FB3D
FB17
FB27
FB41
FB1D
FAD2
FAC6
FB1B
FB7D
FB98
FB8A
FBA5
FBDA
FBB0
FAFA
FA87
FBAF
FEE7
02E0
057F
05CE
04CA
042A
049A
0568
05B4
0578
0539
0529
050E
04E3
04FF
0575
05C8
0593
0523
050C
054E
0559
04E8
046D
0464
04AD
04CA
04A7
04A2
04DC
04F7
04BC
0483
04A3
04D1
0495
0431
046B
0542
055E
0360
FFA4
FC2D
FAAA
FADE
FB45
FAF1
FA50
FA37
FAB2
FB21
FB22
FAF8
FB00
FB1E
FAF7
FA8A
FA4B
FA8E
FB17
FB6C
FB69
FB56
FB70
FBA0
FBAF
FB92
FB5E
FB1E
FAD9
FABB
FAEB
FB3F
FB4E
FB0A
FAF2
FB62
FBD9
FB85
FAAD
FAF4
FD9C
01C0
04DD
055E
0436
0397
047A
05E1
066C
05FC
0571
0553
0554
051F
04E6
0500
053D
0522
04A8
0452
047F
04E0
04E4
0479
0420
0440
04B1
050D
0532
0540
0538
04FA
0498
0468
0494
04D8
04E1
04DA
0518
0541
0437
0156
FDA4
FB1C
FAAB
FB51
FB7B
FAD2
FA36
FA42
FA8B
FA81
FA60
FAB9
FB51
FB4F
FA93
FA26
FAD4
FBFB
FC4A
FB85
FAC8
FB01
FBC2
FC00
FB78
FAD6
FAA3
FAAF
FAB3
FAD7
FB42
FB9A
FB77
FB2B
FB58
FBDD
FBCA
FAD5
FA4B
FBEA
FFBF
03C0
05CC
05AE
04E9
04CA
0542
0591
056A
051D
04FE
050D
0536
057F
05C7
05AA
04FE
043F
042A
04D5
0575
054C
0492
042B
0488
0529
0562
0530
0514
0536
0536
04D4
046E
0478
04BF
04B6
0465
0476
050D
0501
02F3
FF15
FB66
F9D0
FA52
FB4F
FB71
FAD2
FA58
FA6B
FAB3
FACD
FAC2
FAC9
FAE8
FB00
FB0A
FB0B
FAFA
FAD6
FACC
FB0E
FB76
FB9A
FB51
FAF8
FAFD
FB47
FB54
FAF9
FAB2
FAF3
FB78
FB96
FB33
FAF7
FB56
FBD2
FBA2
FB0D
FB87
FE1A
01EB
04E3
05C7
054C
04F4
0555
05CF
05C6
0571
055C
0585
0570
04F4
047E
047D
04D7
0525
053A
0530
051F
050C
050B
0527
052D
04DB
0453
0423
048E
051A
0514
0490
0462
04E7
055F
04E2
03C6
0365
0450
053F
0445
0102
FD25
FAB7
FA2F
FA7E
FA92
FA64
FA73
FAD0
FB0C
FAE6
FAA9
FAB0
FAE0
FADA
FA92
FA71
FABE
FB2F
FB43
FAF2
FABE
FB02
FB80
FBB4
FB7A
FB29
FB10
FB27
FB42
FB5E
FB85
FB91
FB5D
FB22
FB45
FBA9
FBAE
FB28
FB1A
FCE4
0088
043B
060F
05D9
0513
04FA
055E
056F
0517
04F8
054C
057E
051A
048F
049C
0533
058A
053A
04C9
04D8
0531
0524
04A0
0458
04B8
0539
051D
0487
044B
04BF
0547
053B
04CB
0495
04B0
04A9
0471
048E
0514
04E2
02A9
FEBD
FB2F
F9CC
FA57
FB1E
FB07
FA77
FA48
FA84
FA9C
FA69
FA66
FADE
FB68
FB84
FB4B
FB30
FB45
FB30
FAD3
FA98
FAD8
FB4E
FB75
FB48
FB40
FB88
FBA7
FB33
FA7D
FA40
FAA6
FB26
FB51
FB63
FBB4
FBF5
FB97
FAED
FB5B
FDE7
01CD
04FD
0620
05BB
0547
0576
05CB
05AE
0544
0516
0534
053C
050B
04FA
0548
059D
057C
04F4
048C
048C
04AB
049B
0486
04C1
0538
057A
0557
051D
050E
0502
04BD
0476
0493
04F6
050B
04AF
0491
0529
0599
043F
00A9
FC7F
FA09
F9F0
FAD6
FB23
FAA6
FA3A
FA62
FABA
FACA
FAB1
FACD
FB17
FB34
FB12
FAF8
FB04
FAF6
FAA4
FA5F
FA91
FB19
FB69
FB3E
FAF1
FAEB
FB14
FB10
FADE
FAD7
FB15
FB3B
FB13
FAF8
FB55
FBD9
FBC3
FB12
FB02
FCDE
006D
03E8
05A6
0595
04E9
04AA
04E5
0528
0544
055D
0578
0561
050D
04C8
04D9
0524
0554
0551
0553
0582
05A7
0579
0508
04B9
04D1
052A
056C
056E
0543
0506
04C2
0494
04A0
04D2
04D6
0484
043F
0485
050A
049E
0251
FEB0
FB86
FA36
FA7E
FB0C
FB06
FAAC
FA92
FABF
FAD5
FAC2
FACD
FB06
FB18
FACF
FA8B
FABF
FB44
FB7A
FB2C
FADD
FB0A
FB6E
FB63
FAD2
FA5F
FA81
FAE8
FAFD
FABE
FAA8
FAE8
FB1F
FB0D
FB10
FB83
FBFF
FBD1
FB46
FBD0
FE7B
0262
0552
0601
0531
048D
04C9
054D
056F
0550
0562
059D
05A2
056A
0548
054E
051F
049B
0447
04A1
0550
057C
04F2
0472
04A6
0533
054B
04D7
0497
04F2
0556
0518
0481
0468
04E9
0531
04C1
043E
0473
04CA
03A4
006B
FCA8
FA8C
FA95
FB4B
FB36
FA78
FA24
FA91
FAFE
FAC8
FA54
FA65
FAFD
FB67
FB35
FAC0
FA92
FAB3
FACE
FAD2
FAFB
FB52
FB89
FB72
FB44
FB3B
FB35
FAF9
FABB
FAEE
FB88
FBEA
FBBD
FB7A
FBB5
FC0D
FB99
FA78
FA55
FCA8
00BD
042A
0553
04F3
04CE
057C
0611
05D0
0542
0551
05DE
05FB
054F
0491
047F
04E7
0515
04DC
04AD
04CE
04F1
04C8
048D
04AA
050C
053B
0504
04B0
0489
0485
0488
04A8
04EF
050B
04AB
0416
03FD
0483
04EA
049D
0422
0473
0556
0519
026A
FE31
FADE
F9ED
FA8F
FB02
FAA9
FA4F
FAA0
FB32
FB42
FAD8
FA9F
FAD7
FB07
FAD0
FA8A
FABC
FB48
FB8D
FB4C
FAEF
FAE3
FB05
FAF5
FAC1
FACF
FB33
FB82
FB62
FB05
FADE
FB0E
FB5D
FB99
FBB6
FBA5
FB58
FB14
FB48
FBE2
FC18
FB54
FA60
FAFB
FDF6
0206
04E7
059D
0523
04F6
0562
05AA
055F
04FD
051A
0584
0599
0538
04E3
0500
054A
0544
04E6
04A2
04C5
051F
0550
0537
04FF
04D1
04B2
0499
0487
0484
0490
04AC
04D0
04E5
04DA
04CA
04F2
054C
0572
0510
047E
0485
054A
05AC
042E
00AB
FCC8
FA7F
FA3C
FAC3
FACC
FA53
FA29
FA9E
FB22
FB1F
FAC1
FA97
FAC5
FAE9
FAC3
FA96
FABC
FB21
FB62
FB4A
FB01
FAC0
FA9D
FA9B
FAC1
FB01
FB2C
FB28
FB0E
FB07
FB0C
FB03
FB02
FB34
FB74
FB54
FAC3
FA5E
FABA
FB76
FB8D
FAC7
FA76
FC37
FFFD
03D0
05BC
05A3
04F9
04F3
0577
05C4
0594
0541
051D
0514
04FE
04E8
04E8
04DF
04B0
047F
0491
04DB
050D
04FF
04EC
0514
0554
055C
052B
0515
053C
0559
0521
04BF
048E
0495
0493
0483
04B6
0531
055D
04C4
03F3
03FF
04F0
0539
0340
FF5C
FBB7
FA1E
FA58
FADF
FACA
FA7B
FA96
FB09
FB52
FB57
FB5F
FB77
FB56
FAF5
FAC1
FB03
FB6B
FB6F
FB0E
FAC8
FADF
FB03
FAE5
FAB2
FAC3
FB01
FB07
FACA
FABA
FB0E
FB69
FB5E
FB19
FB21
FB80
FBAF
FB6C
FB2C
FB5D
FB99
FB2C
FA71
FAF8
FDD8
021C
056F
0662
05A3
04E2
04E0
0514
04D7
0458
042D
046D
04AE
04B8
04BE
04EA
04FF
04C2
0469
0463
04BE
051F
0546
054F
0561
055B
0518
04D2
04E8
0545
055D
04EF
0467
0450
0491
04A7
047B
047C
04E1
0528
04DB
045F
0479
04E7
0432
0159
FD5A
FA78
F9E8
FAC5
FB58
FB0C
FAA2
FAD3
FB5D
FB95
FB62
FB38
FB5B
FB8D
FB84
FB51
FB2C
FB1F
FB13
FB0F
FB22
FB2A
FAF4
FAA0
FA9A
FB0A
FB85
FB87
FB29
FAF8
FB33
FB7A
FB6C
FB34
FB40
FB87
FB95
FB4F
FB31
FB87
FBD3
FB7A
FAFD
FBD8
FECB
02A7
054B
05C2
0508
04A1
04F3
0546
0513
04AD
04A4
04FA
0547
054F
0530
0509
04CE
048D
0481
04BB
04EC
04C7
0472
0454
0485
04B1
049B
0474
047E
04A4
049B
0469
0461
0499
04B3
0470
0423
043B
0491
0490
042C
0420
04D4
0555
0408
0092
FCA1
FA5A
FA4C
FB29
FB7A
FB0E
FAA3
FAAF
FAEB
FAFB
FAF1
FB05
FB24
FB1D
FB09
FB36
FBA4
FBEA
FBBC
FB4B
FB08
FB1C
FB52
FB75
FB84
FB87
FB72
FB54
FB64
FBB0
FBEB
FBCB
FB7E
FB75
FBBC
FBCF
FB62
FAF1
FB25
FBC4
FBD1
FB03
FAA3
FC57
0017
03E2
05B9
0589
04E0
04F9
0592
05C4
0552
04CA
0499
048C
0453
040F
0420
0493
050A
0531
0512
04E4
04C8
04C2
04D4
04F2
04F9
04D6
04AC
04A2
049F
0460
03EC
03AD
03EB
0455
0467
0426
0421
0496
04F9
04B8
043C
0477
0564
0573
0318
FECD
FAF3
F985
FA39
FB2C
FB1F
FA7D
FA59
FAEC
FB86
FB96
FB50
FB32
FB58
FB7F
FB77
FB4F
FB29
FB12
FB15
FB31
FB3F
FB19
FADA
FADA
FB38
FB97
FB84
FB12
FACA
FAF5
FB47
FB61
FB66
FBAE
FC19
FC1F
FBA2
FB3E
FB73
FBCC
FB76
FAB5
FB17
FDCD
01F4
0533
0601
0513
0444
0491
0567
05C3
056E
04F3
04BE
04BF
04BF
04B9
04C4
04D9
04DA
04BF
048F
0456
042F
044A
04BD
0542
0563
04FE
047E
0462
04AD
04F6
0500
04F4
04FF
04FA
04AF
044A
0431
0462
0468
0416
03F7
0491
054C
04A4
01CE
FDE6
FB09
FA48
FAD5
FB39
FAF7
FAA7
FAD0
FB2D
FB32
FADD
FAA8
FADB
FB40
FB7D
FB82
FB6F
FB54
FB35
FB2B
FB4B
FB79
FB7D
FB54
FB2D
FB24
FB1A
FAFE
FAF8
FB30
FB74
FB6E
FB27
FB16
FB72
FBCE
FBA7
FB2F
FB16
FB83
FBBF
FB44
FAD6
FBFC
FF2C
02F8
055C
05B4
051B
04E4
0544
0590
0560
0507
04EB
04F9
04E0
04A1
0480
0499
04B9
04B7
04AC
04C6
04F5
0507
04EE
04C9
04B5
04B8
04DC
0527
056D
0559
04DC
0463
045A
049A
0497
042D
03EB
0446
04DB
04DB
0443
0404
04A2
0520
03D0
005B
FC6B
FA14
F9D3
FA79
FAC4
FAA2
FAB1
FB23
FB89
FB87
FB44
FB0E
FAEC
FAC0
FA9C
FABA
FB13
FB55
FB47
FB09
FADE
FAD6
FADA
FAE5
FB07
FB39
FB5B
FB6E
FB8F
FBBA
FBB1
FB5E
FB13
FB38
FBAC
FBDC
FB8A
FB3E
FB85
FC06
FBD2
FAD4
FA7A
FC5C
004D
0436
0615
05D4
04FC
04D0
0539
0573
0540
0505
0503
0506
04DA
04B9
04EA
054D
0579
054C
050E
04FC
04FF
04E3
04B0
0497
04A1
04A8
04A2
04A7
04B5
04A5
0475
0469
049F
04CB
0499
0444
045C
04E8
052F
04AE
03F9
0411
04CA
0488
0207
FE18
FB06
FA3B
FAFC
FB90
FB3D
FAAB
FAA1
FB04
FB38
FB14
FAEF
FAFF
FB0D
FAE6
FAB6
FACC
FB2B
FB81
FB8F
FB5C
FB16
FAE5
FAE3
FB17
FB5A
FB69
FB35
FB03
FB19
FB5F
FB79
FB51
FB39
FB6A
FB9F
FB75
FB1C
FB32
FBD7
FC3F
FBB1
FAD5
FB6B
FE66
028F
0587
0621
0556
04DB
053A
05A5
055E
04B6
046E
04A9
04E2
04C5
0490
049A
04C7
04CE
04B1
04B4
04E7
0505
04E2
04A2
047F
047A
047D
048B
04B1
04CC
04AF
047E
0494
04F1
0518
04C4
0462
0482
04EC
04DA
042B
03D3
0488
0556
044F
00D3
FCA2
FA2D
FA19
FAF3
FB28
FAA5
FA57
FAA3
FB07
FB0A
FAE0
FAF8
FB44
FB5F
FB37
FB2A
FB6F
FBC5
FBCF
FB8B
FB3E
FB18
FB13
FB2B
FB66
FBB2
FBDF
FBDB
FBCA
FBC1
FB91
FB1B
FAAE
FAC3
FB50
FBAD
FB6B
FAFB
FB16
FB9E
FBA3
FACE
FA63
FC25
0028
044D
064A
05EF
04FD
04F4
0591
05B1
050F
0485
04BE
0552
0571
0503
04A7
04BC
04ED
04CB
0475
0455
0480
04A4
048F
0471
047E
04A1
04A5
048B
047D
0488
049D
04C4
050D
054D
0538
04E3
04CC
0527
055E
04CB
03D2
03A9
04A4
053F
0382
FF6E
FB61
F9B4
FA60
FB66
FB4A
FA79
FA31
FABD
FB4E
FB49
FB02
FB12
FB6D
FB95
FB65
FB3E
FB65
FB9F
FB91
FB46
FB16
FB2C
FB5F
FB79
FB70
FB5C
FB4C
FB49
FB59
FB5F
FB2D
FACC
FA98
FAD8
FB4B
FB69
FB1D
FAF4
FB51
FBB7
FB61
FA93
FAD8
FD6E
01A3
0530
0666
05AD
04BE
04AB
0511
051A
04B0
0473
04B8
051A
0513
04AE
045E
045F
047F
0485
047F
0498
04C6
04D3
04B2
048E
0497
04C6
04F8
0513
0514
04FD
04DD
04D4
04ED
0502
04DE
0492
046B
0489
04A8
0482
0442
0451
04A4
04B3
043E
03E1
044B
04FC
045B
0179
FD72
FA88
F9EB
FAC3
FB73
FB61
FB21
FB39
FB6C
FB4A
FAF1
FACF
FAFB
FB20
FB15
FB11
FB3C
FB60
FB3E
FAFB
FAF2
FB2E
FB5B
FB43
FB15
FB0D
FB15
FAFC
FAD9
FAED
FB39
FB72
FB76
FB7F
FBB7
FBE1
FBAC
FB40
FB24
FB7F
FBD7
FBB9
FB6A
FB7D
FBDC
FBC7
FB02
FA9E
FC1B
FFA3
038D
05D8
0601
0530
04BE
04EE
0529
0513
04F2
051B
0565
0564
0503
049C
0478
047C
0470
0465
0492
04F0
0534
0531
0513
050D
050C
04E0
0498
0478
0499
04C1
04B8
0499
049A
04B3
04AF
0487
0465
0451
0424
03E3
03E7
0454
04B2
047D
03FC
0407
04BB
04C8
02BC
FEDD
FB48
F9D6
FA5B
FB38
FB58
FB09
FB07
FB53
FB60
FB07
FABF
FAE5
FB3C
FB4F
FB16
FAE2
FADA
FAD2
FAAC
FA91
FAB4
FB04
FB49
FB64
FB64
FB5C
FB49
FB2E
FB1B
FB19
FB1B
FB1A
FB30
FB6F
FBB3
FBC7
FBB1
FBB7
FBF9
FC31
FC0C
FBAD
FB93
FBE1
FBFE
FB5A
FA7D
FAF6
FDBE
01E0
051A
05FF
0539
0483
04B0
051B
04E9
044D
0424
04B6
0552
054C
04D9
04A9
04EF
0539
0525
04DE
04C4
04E3
04FE
04F9
04F1
04FE
0501
04E5
04C2
04B7
04B7
04AD
04A2
04A7
04A3
0475
0441
0451
04A4
04CF
048B
0424
0419
045F
046B
041C
0418
04D7
0581
046E
010B
FCE5
FA55
FA38
FB4A
FBC4
FB3C
FA9D
FAB1
FB2A
FB4C
FAFC
FAC9
FB15
FB90
FBAE
FB52
FADD
FAA8
FAAE
FABF
FACB
FAE2
FB08
FB29
FB33
FB21
FAFC
FAD7
FAD7
FB0E
FB5E
FB8D
FB8D
FB8A
FBA1
FBA4
FB63
FB0E
FB10
FB7C
FBD2
FBA6
FB3F
FB39
FB8F
FB8B
FAED
FAC8
FC94
0056
042A
0601
05A0
049A
0467
04FD
0562
0524
04C0
04C9
0523
054E
0522
04EC
04EB
0501
04F2
04BA
048E
048A
04A5
04C7
04E3
04ED
04DC
04C0
04BC
04D0
04D2
04B0
0494
04B1
04E8
04E2
048C
0447
046C
04CA
04DC
0487
0440
045D
048B
044E
03E8
041F
04EE
04F5
02C8
FED0
FB42
F9F9
FAAB
FB84
FB57
FA9F
FA5D
FAB1
FAEF
FAC6
FA9F
FAE0
FB4B
FB64
FB23
FAF2
FB0A
FB39
FB48
FB4B
FB64
FB74
FB56
FB2B
FB32
FB5C
FB60
FB2B
FB05
FB26
FB5E
FB63
FB47
FB5A
FB9E
FBB0
FB60
FB08
FB11
FB55
FB5B
FB1D
FB1B
FB85
FBC4
FB42
FA96
FB4C
FE42
0262
0576
063A
0566
049F
04B5
052E
0547
04FB
04D1
0509
054D
053E
04FA
04DD
04F8
0502
04D1
0499
04A1
04D9
04FF
04F7
04E8
04F4
0504
04F6
04D2
04C1
04CA
04D6
04D7
04D4
04CB
04AE
048C
048B
04A5
049D
045D
0433
046C
04CC
04C9
0469
0467
0526
05A9
044D
00B7
FC9D
FA3B
FA27
FB10
FB7E
FB38
FAF1
FB0C
FB39
FB29
FB06
FB19
FB4D
FB52
FB1E
FAF3
FAFA
FB14
FB1C
FB18
FB1F
FB2E
FB38
FB3B
FB37
FB14
FAC8
FA89
FAA1
FB08
FB5B
FB56
FB2D
FB3E
FB81
FB97
FB60
FB39
FB70
FBC1
FBA4
FB1B
FAD1
FB32
FBB3
FB73
FA99
FA9D
FCCF
00B9
044E
05D1
0562
0483
0456
04B4
04DD
04A8
0490
04E1
053F
0536
04DC
04A3
04AE
04B5
0481
044D
0475
04F2
0563
0582
0560
0525
04DE
049B
0482
04A1
04C6
04BF
04A5
04BA
04F4
0500
04B9
0470
0472
0499
0485
044A
045A
04BF
04DE
045D
03E9
0469
0572
0535
0270
FE2B
FAEE
FA2E
FB08
FB9B
FB36
FAA4
FAB4
FB2A
FB56
FB26
FB26
FB93
FBFD
FBE4
FB6D
FB24
FB45
FB85
FB8E
FB62
FB37
FB23
FB16
FB10
FB1E
FB37
FB3C
FB24
FB0D
FB0D
FB12
FB03
FAF8
FB1F
FB70
FBAC
FBAE
FB96
FB89
FB6E
FB22
FAE1
FB17
FBB1
FBEC
FB45
FA8B
FB70
FEAF
02E6
05B2
0600
04EF
0449
0494
04F6
04BA
0449
046D
051A
057C
051D
0474
042E
0452
0465
043C
042F
0481
04F1
0515
04E9
04C9
04E4
050C
050B
04ED
04D9
04CE
04B1
048B
047F
0493
04A8
04B2
04C2
04D2
04BA
0477
0456
0490
04D7
04B0
0441
044F
0517
056D
03B8
FFE2
FBE8
F9FE
FA66
FB71
FB99
FB01
FAB8
FB1C
FB87
FB66
FB07
FB02
FB5A
FB8A
FB51
FB09
FB10
FB44
FB48
FB12
FAF4
FB19
FB4A
FB43
FB08
FAD3
FAD1
FB00
FB41
FB72
FB74
FB48
FB18
FB19
FB45
FB63
FB5F
FB6C
FBB2
FBED
FBB6
FB21
FAD0
FB26
FBA0
FB68
FAA1
FAB9
FD07
0116
04BC
0621
057B
0489
048C
052A
055D
04F1
049F
04E1
0547
052C
04B2
0490
0503
0580
057C
0526
0504
0526
0525
04CF
047E
0490
04E3
050E
04EC
04B5
049E
049D
04A3
04BB
04D0
04B3
0468
0447
0482
04C8
04B5
0471
0485
04F4
050E
0473
03E1
0455
0562
0525
025D
FE1B
FAD8
F9EE
FA85
FAFC
FAC3
FA80
FABE
FB27
FB27
FAC9
FA96
FAD2
FB30
FB55
FB43
FB32
FB38
FB3E
FB34
FB28
FB28
FB32
FB37
FB31
FB20
FB09
FAF9
FB01
FB23
FB43
FB49
FB47
FB68
FBA8
FBC5
FB8C
FB35
FB2E
FB8E
FBE6
FBC6
FB5B
FB39
FB81
FB91
FAFB
FA8E
FBD2
FF3A
033B
05A2
05C1
04E2
049B
0522
058E
055A
04F8
04F9
0531
0527
04DC
04C1
04F6
0520
04FA
04BA
04AD
04BF
04AC
0480
048D
04E0
051C
0506
04DB
04E8
0509
04F0
04A8
048A
04A7
04A5
045A
0424
0461
04CE
04D6
0474
044B
04B1
0519
04DE
045D
0487
055F
056B
033B
FF41
FBA3
FA22
FA7D
FB27
FB1F
FAAB
FA7B
FAA2
FABA
FAAA
FAC0
FB1E
FB72
FB6A
FB2A
FB0F
FB26
FB2A
FB05
FAFA
FB3D
FB90
FB90
FB46
FB13
FB22
FB30
FB08
FAE1
FB00
FB43
FB4C
FB1F
FB21
FB79
FBC3
FB9A
FB39
FB1D
FB3D
FB18
FAA0
FA88
FB39
FBF2
FBA7
FAB1
FAE4
FD91
01C2
0508
05F2
0546
04B0
04D5
051C
04FD
04BD
04D7
052B
053B
04EB
04AB
04C8
050B
0513
04E7
04DC
050B
0528
0500
04C6
04C8
04F8
04FE
04C0
0487
0496
04CB
04DC
04C6
04C9
04F1
04F6
04B0
0472
049C
0505
0526
04DE
04A0
04B6
04CA
0480
0440
04AF
0561
04B6
01A0
FD4B
FA3F
F9D3
FAF0
FBA1
FB46
FAC1
FADC
FB4E
FB65
FB1C
FAF7
FB31
FB73
FB6A
FB39
FB2B
FB37
FB22
FAEE
FAD0
FAE1
FAFE
FB09
FB0D
FB1A
FB2B
FB34
FB31
FB25
FB10
FAFD
FB05
FB37
FB7A
FBA0
FB95
FB6A
FB34
FAFB
FAD3
FADB
FB12
FB53
FB7E
FB92
FB8A
FB62
FB49
FB85
FBFE
FC18
FB78
FAE2
FBD5
FEE8
02CA
0552
05A8
04E0
047F
04D2
0523
0502
04CA
04E6
0535
0556
053A
0522
052E
0532
050F
04E7
04ED
051C
0546
0552
053D
050D
04DA
04C8
04D1
04C0
0486
0463
048E
04E1
0510
050D
050D
0522
0518
04D6
04A1
04C2
0500
04E6
046E
0416
0428
045E
0473
0490
04D5
04F0
049E
0454
04AF
052D
0435
00F3
FCCB
FA30
FA14
FB1B
FB87
FB22
FADE
FB1B
FB48
FAFD
FAA2
FABE
FB22
FB3E
FAF2
FAB2
FAD1
FB16
FB22
FAF8
FAE0
FAFB
FB2E
FB5C
FB72
FB5E
FB27
FAFC
FB02
FB23
FB39
FB47
FB61
FB7A
FB73
FB57
FB4E
FB62
FB64
FB3B
FB13
FB1E
FB38
FB25
FB06
FB30
FB81
FB7A
FB1C
FB17
FBB7
FC32
FBBC
FB19
FC26
FF8D
038B
05B1
0582
04AA
04AA
053C
0558
04ED
04CA
0533
0583
053D
04C3
04BA
051C
055F
053C
0502
0506
0530
0536
050D
04D8
04B0
049E
04B0
04DE
04F1
04D2
04B3
04C5
04EE
04ED
04C8
04BF
04EC
051D
051E
04F5
04C8
04A5
0487
0489
04BD
04F0
04E2
04BE
04DE
051A
04E2
043C
0412
04DA
0566
03D9
FFFC
FBE9
F9EA
FA25
FAE5
FAE9
FA9F
FAE1
FB7E
FBA5
FB3A
FAEF
FB20
FB5D
FB2B
FABF
FA9F
FADF
FB15
FAFB
FAC3
FAC0
FAF7
FB35
FB59
FB5C
FB3E
FB15
FB12
FB3B
FB51
FB30
FB0A
FB1D
FB4E
FB54
FB28
FB0E
FB29
FB4B
FB3C
FB0D
FAF7
FB05
FB13
FB21
FB46
FB66
FB50
FB30
FB73
FBF3
FBE8
FB1D
FACB
FC88
0042
03F4
05A3
0556
04A5
04B1
0523
053C
0502
04FA
0531
0536
04E5
04A3
04BE
0509
0532
052C
0525
0531
0534
0517
04E9
04BF
049F
0493
04A9
04CE
04D6
04C6
04D3
0501
0509
04C8
0489
049C
04E2
04F8
04D3
04C2
04F0
051E
050F
04E7
04E9
04FE
04DA
048F
047D
04A6
04A3
0474
04BC
05A0
05E0
03E7
FFD2
FBC4
F9DB
FA20
FAED
FB08
FAB6
FAC0
FB25
FB4C
FB0C
FAD4
FAF4
FB36
FB43
FB16
FAE3
FACB
FAC8
FAD2
FAED
FB16
FB3D
FB4D
FB42
FB21
FAFF
FB02
FB3B
FB7B
FB7E
FB45
FB18
FB1D
FB21
FAFF
FADF
FAEE
FB04
FAE5
FAB0
FAC2
FB2A
FB89
FB99
FB90
FBB0
FBC5
FB78
FB10
FB2B
FBAD
FBA8
FAD7
FA97
FC95
0097
0457
05DB
0562
04B1
04D7
054F
053F
04C6
0496
04DB
0516
04F9
04C6
04D1
050D
053E
0555
056C
0587
0583
0548
04EE
04A9
049A
04BD
04F1
050C
04F9
04D0
04C2
04CF
04CF
04B5
04A7
04B7
04C2
04B3
04B2
04E6
051F
0514
04C8
048A
0474
044E
0409
0407
048C
0519
04F7
0461
045D
051D
0528
02E2
FEC0
FB25
F9EA
FA8F
FB44
FB21
FAC8
FAF9
FB6A
FB69
FAF5
FAA0
FAA8
FABC
FAA5
FA9F
FADC
FB29
FB31
FB04
FAF9
FB33
FB6F
FB65
FB26
FAF3
FAE4
FAEB
FB01
FB25
FB45
FB4B
FB3B
FB2B
FB23
FB28
FB46
FB75
FB95
FB92
FB81
FB7D
FB79
FB62
FB55
FB8C
FBF1
FC0A
FBA4
FB40
FB76
FBE8
FB9D
FA9F
FA8F
FCF1
0121
04B0
05EC
056B
04EE
0534
058F
054D
04C0
0493
04CF
0504
0511
052D
0555
0546
0502
04EA
0534
058E
058E
0539
04ED
04D4
04C2
049B
0491
04C1
04F3
04EA
04C5
04C4
04E5
04F4
04EB
04EC
04F9
04EB
04B2
046D
0444
0438
043C
044C
045F
045B
0444
0460
04CE
0528
04F8
0494
04D6
05A8
0576
02D5
FE80
FAF8
F9F2
FABA
FB5A
FAFA
FA63
FA7C
FB05
FB3A
FAF7
FAB7
FAB4
FAB7
FAA5
FAB2
FAF7
FB3B
FB46
FB2E
FB2A
FB39
FB37
FB24
FB2D
FB59
FB75
FB62
FB48
FB45
FB3C
FB12
FAF3
FB09
FB34
FB3A
FB28
FB2B
FB42
FB3E
FB13
FAF1
FAF2
FAFB
FAFA
FB13
FB5C
FB91
FB77
FB61
FBBD
FC2D
FBCE
FACD
FAED
FDA7
0212
057C
0640
0551
04BA
0526
0596
053E
04A2
0499
0507
053A
050E
04FC
053C
056C
0545
04FD
04E5
04E8
04C2
047A
045C
0485
04BB
04CC
04D4
04F0
0501
04E7
04C6
04CD
04ED
04FF
0503
0510
0515
04F9
04D0
04C2
04C6
04B4
048C
0486
04B1
04D5
04C2
04A7
04B5
04A6
0431
03CD
044D
0555
0511
0230
FDCA
FA88
F9DD
FABD
FB41
FAE6
FA94
FAE3
FB4A
FB26
FABE
FAB6
FB0B
FB39
FB20
FB1B
FB51
FB74
FB4D
FB13
FB13
FB43
FB5E
FB56
FB50
FB56
FB42
FB12
FB01
FB2C
FB57
FB48
FB1E
FB0B
FB0C
FB09
FB19
FB49
FB6C
FB52
FB2A
FB44
FB97
FBC1
FB99
FB65
FB68
FB72
FB45
FB29
FB83
FBEC
FB91
FABB
FB28
FE1B
0277
059A
0627
0535
04A5
04FC
0562
053F
04FE
0527
0576
0560
04F3
04B2
04BF
04CD
04B7
04B3
04E8
0527
0534
050B
04CF
04A0
048F
04B2
0501
0545
053E
04F8
04BA
04A6
049A
048A
049C
04CD
04D9
04A8
048B
04B7
04E5
04B5
0455
0443
0496
04D4
04BB
04A0
04D3
04F2
0481
03F3
043E
051F
04C2
01D9
FD8B
FA7A
F9F2
FAD1
FB41
FAD5
FA6C
FA9B
FAF7
FAF6
FAC8
FAE0
FB2B
FB3B
FB01
FADF
FB03
FB30
FB22
FAE9
FAC7
FADF
FB20
FB59
FB67
FB46
FB1C
FB0C
FB19
FB28
FB29
FB35
FB5D
FB7A
FB5E
FB32
FB45
FB84
FB80
FB1D
FAD2
FAFB
FB4C
FB4D
FB1E
FB38
FB95
FBA3
FB35
FAF9
FB7A
FC19
FBCE
FB03
FB9D
FEB9
02F1
05AF
05F1
0504
049F
050C
0578
0565
0526
051E
052A
050E
04ED
050B
054B
0558
052E
0513
0526
053D
0531
050E
04F3
04E5
04DF
04DD
04DC
04DC
04DD
04E9
04F9
04FD
04EE
04E5
04F2
04F2
04BD
047D
0488
04DE
051F
0516
0501
0515
0511
04AE
043C
044A
04C6
04EC
0469
0404
048D
054D
045D
00ED
FC9C
F9F5
F9D8
FAEF
FB82
FB2C
FAAA
FA97
FACA
FADF
FACE
FACB
FADF
FADE
FAB3
FA7D
FA69
FA84
FAC6
FB0F
FB3C
FB44
FB3B
FB2F
FB11
FAE3
FACA
FADE
FB04
FB10
FB04
FB07
FB22
FB34
FB2C
FB2E
FB5C
FB8D
FB83
FB4B
FB2D
FB36
FB2D
FB11
FB30
FB94
FBB7
FB43
FAC8
FB29
FC39
FCA3
FBA9
FA8C
FB7F
FF0C
0343
05B9
05F4
0557
0525
0551
0544
0501
0508
0576
05CC
059F
0526
04E0
04EF
0518
052D
0541
0566
057C
055E
0518
04D9
04BD
04C1
04CF
04D8
04DF
04E2
04E1
04DD
04DF
04E7
04EA
04E1
04D7
04D4
04C7
049A
0467
046C
04BC
0505
04E2
047B
047B
0515
0544
038E
FFD4
FBDF
F9CE
F9FF
FAFA
FB42
FAD0
FA8B
FAD6
FB2D
FB17
FAD1
FACA
FAEB
FAD8
FA98
FA91
FAE5
FB3B
FB47
FB33
FB48
FB74
FB6A
FB2B
FB13
FB4F
FB99
FB9F
FB76
FB5E
FB54
FB29
FAEB
FAE6
FB2A
FB64
FB56
FB38
FB5C
FBA1
FB92
FB2A
FB01
FB77
FBFD
FBBD
FAF2
FB19
FD62
012D
0471
05BB
0567
04E0
04F3
0547
0546
0505
04FD
0545
0572
0548
050A
0503
0510
04E6
04A3
04B6
0531
0593
0567
04E4
04A2
04CA
04EF
04C3
0485
049A
04F0
0522
0507
04D7
04BE
04A5
0478
046A
049F
04D2
04AD
0457
0456
04B9
04EF
04A7
0477
050B
05C6
04FF
01E1
FDBF
FAED
FA65
FB0B
FB45
FAC7
FA65
FA9A
FAF0
FADC
FA93
FAA2
FB0B
FB4B
FB29
FB0D
FB53
FBB0
FB96
FB0C
FAB2
FAEB
FB5F
FB75
FB1E
FAD1
FADE
FB17
FB26
FB08
FAF1
FAFC
FB1D
FB54
FB9F
FBD6
FBC3
FB7C
FB63
FB9D
FBC6
FB7C
FB0D
FB23
FBB1
FBCD
FAFA
FA53
FBA7
FF4B
035D
058F
0579
04A6
0484
04F8
051F
04CF
04B3
051D
0589
056D
050A
0500
0554
0572
0516
04BA
04DE
0548
0554
04DB
0466
046C
04C1
04F0
04D6
04A9
0491
0481
0477
0490
04C9
04DF
04B4
048D
04B6
04FA
04E2
0478
0461
04F7
059D
057C
04C0
047F
0517
0539
033D
FF4E
FB9F
FA2B
FAB8
FB7A
FB58
FAD9
FAE6
FB5C
FB6E
FAF4
FAA0
FAE2
FB43
FB23
FAAE
FA92
FAF3
FB34
FAEC
FA8C
FABD
FB6A
FBE0
FBBC
FB54
FB26
FB3D
FB58
FB67
FB86
FBA6
FB92
FB55
FB46
FB7D
FB98
FB49
FADD
FAE0
FB4B
FB86
FB4F
FB23
FB74
FBCB
FB58
FA68
FAA2
FD49
0181
04ED
0605
056A
04CB
04EE
0544
0530
04EB
04FF
0554
0559
04F0
04A2
04D7
0539
0537
04DF
04C2
051D
0578
0553
04D5
048C
04B4
0502
0520
050F
04F1
04C7
0495
0488
04C7
051C
0524
04DC
04AC
04CD
04F1
04CA
0493
04BA
0516
0507
047B
0447
0501
05BC
04A8
0130
FCF5
FA4D
F9F3
FAB1
FB1E
FB0A
FB0A
FB42
FB3E
FAD5
FA89
FACC
FB4A
FB5A
FAED
FA9E
FAD1
FB32
FB3B
FAF5
FAD1
FB00
FB39
FB35
FB0F
FB08
FB1B
FB18
FB00
FB01
FB1D
FB18
FAE0
FAC1
FAF6
FB41
FB33
FADB
FAB9
FB03
FB4A
FB23
FAE5
FB2B
FBC6
FBC1
FADC
FA73
FC43
0035
0418
05D0
056D
04AC
04BB
052A
0518
049A
0481
0506
0579
054F
04E6
04E4
053D
0552
04EE
0492
04B2
0515
0534
0503
04E8
051B
0554
0546
0505
04D4
04BA
049D
0498
04DD
054A
056F
0524
04D0
04E0
052C
053C
04FE
04E2
0516
0520
04A1
0425
048A
0587
0561
02B4
FE4F
FABA
F9B8
FAAD
FBA4
FB93
FB0E
FAFD
FB56
FB6A
FB00
FA9C
FAAB
FAF7
FB15
FB0C
FB29
FB6A
FB74
FB1D
FABA
FAB0
FAF6
FB38
FB48
FB3F
FB33
FB14
FAEA
FAE4
FB0C
FB21
FAEE
FAB0
FACD
FB3C
FB83
FB63
FB2C
FB3B
FB59
FB14
FA9A
FAA8
FB6E
FC01
FB7E
FA97
FB37
FE5A
02A6
059B
060F
0516
0470
04AF
051E
051A
04D2
04BD
04DD
04E7
04D2
04DF
051C
0545
052B
0502
050F
0539
0534
04FC
04DA
04F3
0507
04DA
0490
047E
04AE
04E2
0503
0541
05A4
05D1
0579
04E5
04AC
04E9
0516
04D6
0482
049D
04F3
04D7
0441
0417
04D8
0575
041E
0074
FC53
FA15
FA44
FB68
FBED
FBA9
FB60
FB6F
FB75
FB28
FAD0
FAC7
FAEC
FAE1
FAAC
FAA4
FADD
FB00
FAD0
FA99
FAC2
FB30
FB66
FB2B
FAD5
FAC8
FB02
FB3B
FB55
FB62
FB58
FB10
FAA2
FA78
FACA
FB43
FB65
FB2C
FB05
FB1D
FB24
FAE5
FAC8
FB3E
FBE9
FBDE
FB0F
FADE
FCCB
008D
0412
0588
051F
046E
0485
0506
0521
04CD
049D
04CC
04FF
04F4
04EB
052A
0573
0550
04C9
046E
049C
0509
0539
051E
0506
0513
051A
04FF
04EB
0505
0531
0540
053B
0546
054A
050B
049A
0462
049C
04F2
04F2
04B8
04B8
04FC
04F2
045E
03F2
047F
0584
053D
0283
FE60
FB36
FA62
FB12
FB9A
FB5B
FB05
FB34
FB89
FB5A
FABF
FA6D
FAB0
FB07
FAE8
FA7F
FA65
FABF
FB22
FB35
FB24
FB3C
FB6B
FB68
FB2C
FAFF
FB0D
FB2F
FB33
FB21
FB11
FAF4
FAB5
FA88
FAB8
FB2D
FB70
FB4E
FB21
FB3F
FB6E
FB3E
FADC
FAF5
FBA5
FC08
FB65
FA93
FB73
FEBE
02DC
0563
0591
04C8
04A6
0547
05A5
0543
04C2
04DD
0563
0590
0523
04A7
04A7
050E
0564
0576
056B
0562
0540
04EF
0494
046F
0492
04DC
052A
0565
0571
053E
04EA
04BC
04CF
04EC
04DC
04BD
04DB
052B
054A
0512
04E3
0518
055F
0519
045C
0412
04AF
0512
037E
FFC2
FBDE
FA14
FA92
FB93
FB94
FAD7
FA7F
FADD
FB2E
FAE5
FA6D
FA72
FAE5
FB29
FAFB
FAB8
FABD
FAF1
FB10
FB17
FB2A
FB3D
FB22
FAE5
FACA
FAEC
FB0F
FB04
FAF4
FB19
FB4C
FB36
FADE
FAB3
FAF0
FB38
FB1F
FACB
FAC3
FB22
FB63
FB2F
FAEF
FB36
FBC2
FBB9
FB0C
FB1A
FD51
014C
04DD
0633
059F
04DD
04F8
0566
053B
0494
0453
04D1
0568
056D
0511
04F0
052B
054F
051B
04DA
04E0
0507
04F3
04AB
048C
04BB
04F5
04FF
04FE
0520
053C
051A
04E1
04F3
0546
055E
04FB
048E
04A7
0526
0568
052C
04E4
04EA
04EB
0482
0410
0448
04DE
0452
019A
FDAB
FAC9
FA30
FAF3
FB56
FAD7
FA59
FA9A
FB34
FB53
FAED
FAA9
FADE
FB20
FAFA
FA9F
FA9E
FB14
FB87
FB91
FB55
FB32
FB46
FB62
FB66
FB53
FB28
FADA
FA8C
FA87
FADF
FB40
FB4F
FB28
FB2C
FB74
FB9F
FB65
FB09
FAFD
FB3D
FB61
FB47
FB48
FB8E
FBA4
FB2E
FAE3
FC31
FF88
0372
05CA
05E4
0507
04BE
0535
058D
0551
0502
0528
057E
0563
04D5
047E
04C6
0551
057E
052C
04B6
0470
0465
0485
04C6
04FE
04F1
04A2
046C
0497
04F3
051A
0501
04FE
052C
0532
04C9
044D
0454
04DE
0543
051C
04C4
04BD
04DF
049F
0413
0401
04A3
04CF
030C
FF6F
FBE3
FA44
FA8C
FB30
FB11
FA80
FA5C
FAC1
FB0B
FADF
FA9C
FAB8
FB1A
FB57
FB4F
FB41
FB54
FB66
FB5B
FB57
FB7B
FB9E
FB90
FB71
FB86
FBC4
FBCA
FB6B
FB00
FAED
FB19
FB1E
FAF2
FAF9
FB56
FB90
FB36
FAA0
FA88
FB0A
FB75
FB55
FB29
FB9B
FC57
FC53
FB74
FB40
FD58
0162
0523
06B3
063D
0554
0508
0526
051B
04E8
04E7
0514
0511
04C9
0494
04AB
04D0
04B1
046C
0460
04A1
04DD
04D7
04B0
0497
0483
045C
044A
0483
04E2
0503
04D8
04CA
0519
0569
053C
04BE
04A6
0523
0583
052A
048F
0495
04FF
043E
0140
FD10
FA11
F98B
FA83
FB2C
FAEF
FA99
FAE0
FB6A
FB81
FB1B
FACE
FAEC
FB2E
FB44
FB44
FB66
FB90
FB84
FB4C
FB33
FB51
FB6C
FB5C
FB45
FB56
FB72
FB6B
FB55
FB6B
FB9A
FB88
FB29
FAF6
FB43
FBB0
FB9A
FB14
FADD
FB45
FB94
FB1B
FA98
FBC7
FF45
036C
05CA
05A8
048B
0448
0518
05DC
05C7
053B
04F9
0524
0553
0549
0524
0503
04D4
0499
0484
04A7
04C5
04A2
046A
047C
04DA
0520
0507
04BE
0497
048F
047D
0477
04BA
0525
0539
04CA
045C
0479
04D9
04BE
0425
03FE
04C9
0565
0403
0058
FC58
FA4D
FA91
FB83
FBA0
FAFE
FA9C
FADF
FB40
FB3A
FAF9
FAE2
FAFE
FB12
FB1D
FB4E
FB90
FB90
FB3D
FAFC
FB27
FB88
FBA8
FB72
FB3F
FB42
FB41
FB09
FAD4
FAF6
FB53
FB82
FB69
FB61
FB96
FBB1
FB6D
FB2A
FB70
FBF8
FBD4
FADE
FA82
FC62
004B
0407
059D
053E
04A7
04EF
058F
058D
04E8
046F
048F
04E0
04E9
04C2
04BC
04CB
04B1
047F
0485
04C7
04E1
04A3
046D
04A5
051B
053C
04E3
0487
0485
04A3
0484
0447
0454
04A7
04CA
0499
0482
04D1
0519
04D2
045D
04A4
0587
055D
02B2
FE53
FADB
FA07
FB0D
FBD5
FB70
FAB5
FAA8
FB1B
FB42
FAF5
FAC9
FB10
FB67
FB6D
FB51
FB6D
FB9F
FB7D
FB15
FAF0
FB48
FBA8
FB9E
FB5D
FB62
FB9C
FB89
FB0F
FAC5
FB22
FBC9
FC07
FBCA
FBA2
FBCA
FBD1
FB6E
FB1D
FB62
FBCE
FB82
FAC2
FB31
FDFD
021A
0512
059E
04D5
0492
0540
05D9
0596
04EC
04AD
04E1
04FD
04D0
04B9
04E6
0501
04C2
0471
047A
04BF
04CC
0494
0480
04C1
04F5
04C3
0475
048C
04F5
050D
049C
0432
045C
04D5
04F6
04B9
04B5
0516
0544
04D7
0469
04C1
054E
0459
0113
FCF7
FA73
FA5E
FB53
FB93
FAF3
FA7A
FABD
FB35
FB38
FAE7
FAC8
FAEF
FB08
FB02
FB23
FB71
FB7A
FAFF
FA75
FA82
FB1A
FB91
FB89
FB5C
FB73
FB9D
FB68
FAF3
FACF
FB2F
FB95
FB92
FB68
FB8C
FBD1
FB9C
FAF2
FA9F
FB0F
FB89
FB39
FABE
FBDE
FF54
0384
05F2
05E4
04E7
04BB
056E
05D5
0560
04B5
0495
04E4
0510
04FC
04F7
0515
050A
04CC
04C1
051A
0563
051F
0490
0473
04F1
055F
052C
04AF
049B
04FC
052E
04E0
047C
0471
0486
0455
0410
0442
04D7
0514
04B6
0477
04ED
052E
038D
FFD1
FBFD
FA54
FAE8
FBCB
FB7A
FA68
F9EB
FA62
FAFE
FB1B
FAFA
FB0E
FB37
FB1B
FADC
FAE1
FB19
FB07
FA93
FA52
FAB5
FB56
FB7C
FB23
FAF4
FB33
FB57
FAE3
FA44
FA49
FAFD
FB99
FB99
FB59
FB5D
FB87
FB68
FB1E
FB37
FBA9
FBB7
FB2A
FB31
FD33
00E6
0445
05A6
0566
0516
056A
05B2
053B
047A
045D
04FE
0590
058F
054C
0548
056B
054E
04F2
04BF
04D8
04EC
04C6
04B2
04FE
0570
058E
0552
0533
0564
0583
0533
04B9
04A0
04ED
0511
04C1
0461
0463
04A1
04B7
04C2
0527
058C
04B1
01CF
FDE7
FB07
FA3F
FAAE
FAD1
FA53
FA0C
FA88
FB3A
FB51
FADC
FA97
FAD8
FB32
FB31
FAF8
FAE7
FAF7
FAD5
FA81
FA61
FAA5
FAF7
FAF3
FABB
FAB9
FB00
FB2E
FB05
FAC2
FAB5
FAD0
FADA
FAE4
FB27
FB87
FB99
FB4B
FB21
FB70
FBB9
FB4E
FAAC
FB6C
FE76
0295
0572
05F6
0532
04D2
0534
057A
051C
04A9
04C8
053C
0551
04EE
04AE
04E3
0528
050F
04DD
0519
05AB
05E8
0581
04F6
04E2
052B
054E
052D
0526
0568
059D
0570
050C
04C9
04A9
0472
043F
0469
04DC
04FD
0499
0460
04EA
056F
043C
00CA
FCCB
FA8A
FA81
FB1B
FAE7
FA36
FA38
FB12
FBB0
FB55
FA9A
FA7C
FB02
FB5C
FB22
FACB
FAD9
FB18
FB15
FAE4
FAF5
FB4F
FB73
FB1F
FAB1
FAA0
FAD0
FAD4
FA9E
FA96
FAF2
FB5E
FB7D
FB60
FB48
FB30
FAFC
FAED
FB58
FBEA
FBC8
FAD9
FA86
FC77
007A
0447
05CD
0549
04B0
0537
0626
0633
0551
04A1
04DE
0587
05B6
0547
04C6
048D
0477
0459
045D
04AA
050D
0535
0521
051A
0538
0547
0522
04F2
04EF
0510
0527
0529
0520
04F7
0494
0433
043D
04B1
04F1
048A
0401
044E
0556
0578
0328
FEDF
FB00
F988
FA36
FB37
FB4D
FAD2
FAB6
FB17
FB4A
FAF6
FA8C
FA9B
FB11
FB70
FB77
FB54
FB36
FB0E
FACB
FA9B
FAB3
FAFD
FB2D
FB25
FB12
FB1F
FB3A
FB39
FB1A
FAFE
FAFC
FB19
FB5E
FBBE
FBF0
FBA8
FB14
FAD9
FB50
FBE6
FBC1
FB12
FB53
FDC5
01C0
050B
060D
054D
048D
04C6
0565
0573
04EA
0480
049D
04EB
0501
04ED
04F4
050F
0500
04CC
04BF
04F5
052E
052B
0505
04FA
04FF
04DD
0494
0473
04A5
04F2
0514
0513
0516
0510
04D8
048F
048B
04C3
04B9
043D
03F4
048A
0562
04BA
019C
FD4C
FA41
F9B4
FAA5
FB57
FB3E
FB0C
FB48
FB89
FB4C
FAD0
FAB9
FB17
FB5C
FB3A
FB08
FB2E
FB82
FB8C
FB39
FAE7
FAD0
FACC
FABC
FAD6
FB42
FBB5
FBC2
FB77
FB4A
FB71
FB93
FB5D
FB06
FAF9
FB2E
FB40
FB1F
FB36
FB9F
FBBE
FB23
FA9D
FBC0
FF0D
030B
0595
05F5
054C
0501
0549
0576
052B
04C9
04B3
04C4
04A8
0469
045C
0495
04D0
04D8
04CF
04E3
04FD
04EE
04BE
04AB
04C8
04EA
04F1
04F0
04FD
0501
04E0
04B6
04AF
04C0
04B0
0485
0496
0503
0557
050D
0462
0434
04CE
0525
03BC
005F
FC9B
FA54
FA0C
FAB8
FB24
FB11
FAF5
FB20
FB69
FB94
FBA3
FB9F
FB6F
FB0C
FAC3
FAEF
FB73
FBC9
FB9A
FB2C
FB07
FB48
FB8B
FB7A
FB2A
FAE9
FAD0
FAC2
FAB3
FABB
FAE3
FB11
FB33
FB5F
FB8E
FB83
FB1A
FAA8
FAB6
FB40
FBA0
FB82
FBAA
FD4A
0074
03A8
0543
0529
04AE
04E2
0573
0576
04CB
043C
045E
04D8
04FD
04B3
0467
0457
0452
0437
044B
04C4
0553
0578
052A
04E4
04F6
052A
0526
04F0
04CC
04C4
04A9
047F
048D
04E1
051A
04E7
0486
046F
04A2
04B7
049D
04CB
0552
052B
0311
FF38
FB91
F9FC
FA72
FB5B
FB7F
FB1D
FB18
FB9E
FC14
FC08
FBA8
FB4D
FB01
FABD
FAC1
FB3C
FBCF
FBD4
FB34
FA98
FA99
FB0C
FB55
FB3A
FB10
FB13
FB14
FAEA
FAE1
FB4D
FBE6
FC09
FB9E
FB41
FB5E
FB81
FB0F
FA7E
FB41
FE1A
01EB
04A4
0552
04D5
0496
04F1
053A
04F2
0477
0463
04BF
050C
0500
04C1
048D
0467
044C
0463
04BF
0514
04FB
0487
044C
04A8
053C
055B
04EE
0493
04C9
054D
0575
050C
047D
0430
0425
0448
04C2
0588
05BD
042A
00AA
FCCF
FA9D
FA96
FB64
FB81
FAD7
FA6E
FAD6
FB7D
FB96
FB2C
FAEC
FB1E
FB57
FB36
FAF4
FAFD
FB45
FB61
FB29
FAEE
FAFD
FB37
FB58
FB60
FB72
FB77
FB32
FAB9
FA7E
FAB2
FAFC
FB07
FB0F
FB77
FBF4
FBB9
FAC8
FA93
FCA5
00AC
0467
05D7
0527
041A
03E9
0443
045B
0430
0463
0515
05A0
0580
0501
04C1
04DB
04EF
04D0
04BB
04D6
04DF
0496
043B
043E
04A3
04F3
04E9
04C7
04E5
0528
053B
051A
050E
0518
04DE
045C
0436
04E4
05A1
04CC
01B2
FDA8
FAEC
FA72
FB2D
FB8D
FB30
FAD5
FB01
FB54
FB4A
FB13
FB32
FB9A
FBA7
FB10
FA6C
FA6F
FAFA
FB52
FB2D
FB0D
FB68
FBE8
FBDB
FB41
FADD
FB32
FBD2
FBF6
FB80
FB03
FAE4
FAF7
FB04
FB2B
FB7C
FB7E
FACF
FA2E
FB30
FE7E
02AA
0558
05A4
04D0
0493
0530
05A4
0555
04CB
04BC
0504
0503
04A4
0476
04BE
050D
04EC
0491
047D
04AF
04B7
047A
046D
04D7
0543
0517
047E
0437
0481
04C7
0485
041C
043E
04D6
0521
04E1
04C5
0542
056D
03C6
0026
FC58
FA61
FA83
FB53
FB8D
FB31
FAF0
FB04
FB0F
FADC
FAA7
FAB2
FAE2
FAFC
FB06
FB28
FB54
FB58
FB37
FB2A
FB44
FB4C
FB1B
FAE7
FAF8
FB34
FB3B
FAFF
FAE7
FB35
FB8A
FB62
FAEA
FAE5
FB96
FC26
FB9F
FA74
FA73
FCEB
010B
047D
05A9
050D
044F
0456
04B7
04C0
047E
0479
04D2
0517
0501
04DC
0510
0574
0580
050E
0493
048E
04E9
0535
053E
0530
0537
0540
0528
04F8
04CA
049E
0474
0479
04CC
0522
04F7
045A
041A
04C7
059A
04E2
01D9
FDD0
FB12
FAA0
FB6C
FBCD
FB57
FAE2
FB17
FB92
FB96
FB22
FAD2
FAE9
FAFD
FAB5
FA64
FA95
FB33
FB94
FB5B
FAEC
FAD5
FB0F
FB23
FAE0
FA99
FAA4
FAE5
FB19
FB3A
FB5F
FB6D
FB39
FAE8
FADB
FB0E
FAFB
FA6F
FA48
FBDB
FF58
0335
0580
05B4
04EF
0487
04BB
04FA
04E2
04AE
04AD
04CD
04DB
04DD
0500
0530
052B
04EB
04CA
0508
0568
0575
0520
04D5
04EC
053A
054E
0503
049B
0455
042E
041A
0439
049F
0503
050D
04EB
0532
05E1
05D6
03C9
FFEC
FC28
FA67
FABE
FBA0
FBBC
FB32
FAE1
FB0A
FB2A
FAF0
FABF
FAFF
FB71
FB7E
FB17
FAC5
FAE0
FB20
FB1C
FAF0
FB00
FB4B
FB5F
FB09
FAAA
FAB8
FB22
FB73
FB7C
FB75
FB81
FB76
FB3A
FB17
FB44
FB5B
FACF
FA05
FA76
FD2E
014E
048D
056C
049A
03E8
0436
04CE
04B9
041C
03E4
0475
0539
0583
0554
0522
0511
04EE
04B2
04AA
04F4
0540
0535
04F4
04DD
04F1
04D9
0481
0451
0493
04F0
04EA
0497
0489
04EC
0540
0528
050D
0572
05C6
049D
0161
FD5A
FA9F
FA14
FADA
FBA0
FBEB
FBF9
FBEA
FB8D
FAF4
FA9B
FAC9
FB25
FB34
FB02
FAF7
FB1F
FB13
FAAC
FA62
FAB8
FB74
FBD0
FB70
FAC8
FA7B
FA9D
FAD9
FB16
FB80
FBFB
FC03
FB66
FAC1
FAD2
FB61
FB64
FA76
F9D5
FB45
FF00
0325
057F
05A1
04E8
04B4
0513
0541
04EE
0491
049C
04E7
050A
04ED
04BF
0492
045A
0434
0468
04EE
0556
0550
0524
054C
05BE
05ED
058A
04F2
04AA
04AD
0497
0462
0474
04E8
052A
04C6
0443
049F
05B9
05E4
038E
FF3B
FB5C
F9F3
FAB6
FBB7
FBA3
FAE5
FAA2
FB21
FBA5
FB87
FAFD
FAAF
FAE8
FB6E
FBE6
FC13
FBD0
FB2A
FA88
FA74
FAFC
FB80
FB5F
FAC2
FA62
FA91
FAE3
FAEA
FAE3
FB39
FBB1
FB9F
FAF4
FA85
FAE1
FB66
FB1A
FA5A
FAE1
FDBD
01C8
04BE
0593
0537
0504
052D
0511
048E
044F
04C3
0571
059D
053D
04D9
04B7
049E
0465
044D
048B
04DD
04D6
0485
0467
04B5
0514
0519
04E6
04E9
051F
050E
0485
040E
0442
04E8
0536
04F1
04DA
0589
0629
04F8
0157
FCEE
FA3B
FA1E
FB31
FBA2
FB21
FAAE
FAF0
FB6B
FB67
FAF7
FAC0
FAFA
FB3E
FB37
FB13
FB12
FB18
FAFB
FAF1
FB46
FBBD
FBC3
FB38
FAB7
FAC7
FB24
FB33
FAFE
FB25
FBD2
FC4B
FBEC
FB29
FAFA
FB69
FB70
FA98
FA1A
FBC1
FFA6
03B9
05C3
058F
04B4
0492
050F
054F
0508
04B0
04A5
04BA
04A9
0489
0499
04CB
04E6
04E5
04F6
0513
04FC
04A9
0486
04D6
053A
0517
0489
044C
04B2
0514
04BF
040E
03FE
04BD
0548
04DD
0430
0475
056D
0537
028A
FE7A
FB71
FAA2
FB1B
FB57
FB00
FAC6
FB08
FB52
FB31
FAEC
FB06
FB74
FBAF
FB7C
FB2D
FB1D
FB46
FB73
FB94
FBB3
FBB2
FB67
FAF4
FAC1
FAFF
FB51
FB42
FAEE
FAE4
FB5B
FBCF
FBAC
FB2B
FB1A
FBB5
FC20
FB7E
FA6E
FACF
FDBE
0206
0521
05BD
04D7
044B
04BF
0570
0599
055F
0540
0530
04D5
044E
0428
0484
04D4
04B2
0480
04C9
054D
0543
047C
03C4
03DF
0490
0506
04EB
04A9
0496
0482
043F
0421
047B
04EE
04D4
0450
0454
053B
05D4
0467
00C0
FCB6
FA76
FA71
FB51
FBA5
FB37
FABB
FAB4
FAF8
FB22
FB15
FAF9
FAF0
FAFB
FB10
FB2C
FB44
FB4A
FB4B
FB65
FB91
FB9B
FB66
FB28
FB2A
FB6B
FB98
FB80
FB5F
FB83
FBD5
FBEE
FBB1
FB7F
FB9D
FBAF
FB24
FA42
FA55
FC7E
004E
03E7
059F
0568
0490
0459
04E5
0578
057C
0514
04D2
04FE
0557
055F
04E5
043A
03E0
0416
04A2
0519
053D
0513
04C6
047E
0459
0467
04A5
04EE
0505
04BC
0438
03E8
0424
04C0
0528
0508
04BF
04E1
0537
0494
0219
FE83
FBB6
FACF
FB1C
FB33
FAAE
FA53
FAA5
FB16
FAE8
FA58
FA4D
FAFC
FBA0
FB9F
FB5C
FB79
FBCC
FBAA
FB0B
FAB5
FB24
FBCF
FBE6
FB65
FAF7
FAF5
FB0A
FAEC
FADD
FB1F
FB66
FB4D
FB19
FB5C
FBE0
FBAF
FA7B
F99B
FAF0
FEB4
02EF
0551
0568
04AC
049B
0547
05C3
0589
0502
04DC
052B
0575
055D
050E
04E3
04E1
04C0
0465
041D
0439
049F
04E9
04E2
04C3
04D7
0510
0520
04F0
04BC
04B2
04BA
04BC
04E7
055E
05AD
04E3
0283
FF31
FC50
FACE
FA86
FAB1
FACF
FAE6
FB15
FB39
FB1A
FACB
FA99
FAAA
FAD4
FAE5
FAE7
FB06
FB3C
FB47
FB04
FAB0
FAA6
FAF5
FB57
FB90
FBA6
FBAA
FB85
FB2A
FADE
FAFF
FB81
FBD0
FB71
FAC4
FAE6
FCB4
FFE3
0320
0513
055D
04B9
0441
0478
04FC
052A
04EE
04CD
0520
0597
05A6
0549
0500
050F
0524
04E0
047F
0486
04EF
051E
04C6
0468
0494
0518
0551
0518
04E0
04E1
04C6
045E
0437
04D0
0564
0447
00DC
FCB9
FA3B
FA2E
FB3F
FBBD
FB4F
FACD
FADD
FB3D
FB57
FB10
FAC7
FAC2
FAE1
FAF2
FAFA
FB1F
FB62
FB90
FB78
FB2A
FAF5
FB0E
FB53
FB78
FB67
FB50
FB4F
FB47
FB2C
FB37
FB88
FBBB
FB4D
FA9A
FB0E
FDBA
01CE
0506
05E3
051F
0491
0501
059F
057E
04E0
04B3
0529
058A
054B
04D3
04CD
0529
0546
04ED
04A3
04DC
0545
053B
04B1
044B
047A
04E6
04EF
0486
043B
045D
0494
0476
0448
04A4
055C
0526
02E1
FF0B
FB9A
FA2E
FA9F
FB68
FB61
FAB4
FA3F
FA6E
FAE9
FB36
FB42
FB3D
FB3D
FB2D
FB08
FAE6
FAD4
FAC3
FAA7
FAA0
FADE
FB55
FBB4
FBB6
FB6E
FB2E
FB21
FB20
FB03
FAEF
FB30
FBA4
FBB1
FB21
FADD
FC54
FFCC
03AD
05DC
05CC
04D8
0497
052A
0592
0543
04CA
04DA
053E
0543
04CF
0483
04CC
054C
0560
04FA
049C
049F
04CE
04CC
04A1
049A
04C7
04E2
04C0
0497
04B2
04FC
0519
04EF
04E1
0546
0597
0495
0196
FD9E
FABA
FA18
FAEC
FB7D
FB12
FA71
FA8E
FB37
FB7B
FB07
FA83
FA90
FAF0
FB0E
FAEA
FAFF
FB63
FB98
FB4E
FAE8
FAF3
FB5C
FB8C
FB49
FB03
FB20
FB65
FB54
FAFD
FAE9
FB43
FB77
FAFC
FA54
FAD9
FD65
0136
0469
059F
0529
0476
0480
0508
0543
04FE
04C3
04FF
055D
0551
04E9
04BD
050C
0561
0542
04E1
04C4
04FA
0512
04D7
04A5
04D1
0514
04EF
0481
0470
04F2
055B
0508
0463
046D
053E
057F
03BB
0020
FC86
FAB6
FAD2
FB87
FB9E
FB16
FAB3
FADC
FB38
FB41
FAFB
FAD3
FAFA
FB28
FB0C
FAC5
FAAC
FAD4
FAF4
FAE0
FACE
FB02
FB56
FB6D
FB31
FAEB
FAD3
FACA
FAAC
FAB6
FB31
FBD7
FBE5
FB23
FA96
FBBA
FEE3
02A8
0521
059E
0513
04D0
052F
058C
055C
04E0
04AC
04DA
0501
04EA
04DD
0522
0575
055C
04DD
048B
04C5
0529
051F
04B3
0488
04E3
0548
052F
04CD
04B9
0502
0515
04B3
046F
04E0
057E
04D1
0207
FE12
FAEB
F9C9
FA3C
FAF8
FB26
FAEB
FAD3
FB0A
FB42
FB2C
FAE4
FABB
FAC8
FADA
FAD7
FAE7
FB2F
FB81
FB8C
FB51
FB2B
FB4F
FB79
FB57
FB10
FB0B
FB3F
FB39
FAE7
FAE7
FB91
FC2B
FBB1
FA79
FA61
FCE0
0126
04C0
0610
05A8
051F
0525
053C
04F0
0499
04BA
0535
0579
054A
0506
0514
0555
0556
04EC
046B
043C
0466
0494
047F
0443
043B
048F
04FB
0518
04DF
049E
0485
0478
046E
04A4
0521
0524
0397
004E
FCA0
FA57
FA06
FAB5
FB24
FB0C
FAE9
FB04
FB1B
FAF9
FAD2
FAE9
FB1C
FB1C
FAF2
FAFB
FB60
FBC3
FBBD
FB68
FB37
FB4E
FB5E
FB2B
FAFB
FB31
FBAC
FBD5
FB6A
FAFC
FB41
FC05
FC34
FB46
FA50
FB38
FE97
02D1
058C
05EB
051A
04B3
0514
0576
0548
04E6
04E0
0520
0517
04A1
0441
046F
04F4
0536
04F7
0496
0488
04C6
04E7
04B9
047F
0491
04E3
0516
04FC
04C6
04A9
0491
045E
0450
04C8
0571
0508
028B
FE9C
FB41
F9F6
FA54
FAD6
FAB2
FA63
FA8F
FAFE
FB0A
FAAF
FA90
FAFD
FB77
FB79
FB38
FB3D
FB8A
FB9F
FB49
FAF6
FB09
FB3F
FB13
FA91
FA58
FAC7
FB67
FB81
FB14
FAD8
FB41
FBCB
FB9A
FABB
FA81
FC59
0026
040E
0618
05FC
052A
0502
0585
05CA
056F
0500
0509
054C
0539
04D5
04B1
04FE
0534
04E0
0458
0445
04AD
04F9
04D8
04B2
04FF
058E
05BE
055F
04EE
04E2
0504
04D0
0450
0434
04D5
055E
045B
013B
FD2B
FA3E
F992
FA63
FB09
FAC0
FA26
FA1C
FA99
FAEE
FAD4
FABA
FB02
FB64
FB64
FB13
FAF5
FB35
FB67
FB41
FB13
FB4B
FBAE
FBA6
FB1F
FAAF
FAC7
FB17
FB16
FADC
FB01
FB9D
FBEB
FB47
FA67
FAF9
FDE4
0212
054E
0650
05BA
051B
0537
0587
0558
04DA
04CC
0552
05B2
0565
04D8
04CC
0537
0551
04C1
042F
045C
0501
0528
0492
0418
0477
0538
0555
04AB
041D
0452
04D9
04EA
0494
049D
0533
0536
034C
FF93
FBD6
F9EF
FA18
FAFD
FB41
FAC6
FA5F
FA95
FB07
FB14
FABA
FA85
FAB1
FAEB
FAEB
FAEB
FB34
FB8F
FB8E
FB43
FB36
FB95
FBD4
FB75
FADF
FAD6
FB4D
FB69
FAD8
FA78
FB1F
FC33
FC46
FB20
FA6A
FBF7
FFA4
0366
055B
056D
04E4
04CA
051C
054E
0527
04EE
04FD
054F
057E
0541
04CF
04A4
04DB
0510
04F0
04B5
04BF
04F5
04E0
046F
0438
04B0
0567
058A
0503
0498
04C6
0510
04D9
0477
04A9
0528
0474
0196
FD98
FABB
FA35
FB19
FBA9
FB45
FAB5
FAC2
FB36
FB54
FAF2
FA97
FAAC
FAF1
FAEF
FAB0
FAB3
FB25
FB8A
FB67
FAF7
FAE1
FB3F
FB78
FB26
FABF
FAE3
FB64
FB77
FAED
FA95
FB15
FBCF
FB97
FA91
FA89
FCF7
0121
04A8
05F2
0573
04B6
0496
04C7
04C2
0499
04BB
0536
0594
0577
0515
04ED
051E
0546
0510
04AB
0491
04D7
0504
04BF
046E
04A7
0538
0553
04C8
0468
04D4
0566
0515
0426
0417
0569
0650
0484
002E
FC0B
FA6A
FAE3
FB7A
FB47
FAFF
FB49
FBAB
FB73
FAD4
FA95
FAE3
FB21
FAE9
FA9E
FAC6
FB3E
FB7F
FB64
FB40
FB49
FB5F
FB51
FB24
FAF8
FADF
FAD6
FAD0
FACD
FAE4
FB2D
FB84
FB7F
FAEF
FA81
FB7C
FE77
0254
0506
058E
04D9
046D
04B6
04FF
04CC
0483
04A7
050A
051F
04DC
04C4
0516
0560
0522
048C
043F
0474
04C7
04DA
04CA
04E2
0517
051C
04E7
04D0
0514
0567
0550
04DE
04BC
053F
05A5
0499
01AC
FE08
FB71
FAB0
FB18
FB85
FB7A
FB42
FB34
FB3E
FB2F
FB12
FB09
FB07
FAE0
FA99
FA75
FAA1
FB00
FB4C
FB5E
FB51
FB58
FB75
FB6E
FB1C
FABE
FABA
FB13
FB52
FB22
FAD7
FB03
FB7E
FB6B
FA95
FA5E
FC81
00C3
04B8
0632
057A
0486
0486
04F1
04F3
04B5
04DB
0541
0533
04AE
0482
050B
0587
053D
049A
0480
04EB
0510
04A8
0455
049B
0519
052F
04E8
04C4
04CC
049F
0460
04AD
0556
04DC
0217
FDF3
FAC3
F9DE
FA8C
FB41
FB50
FB17
FB00
FB04
FB02
FB0D
FB28
FB1B
FADE
FAC7
FB0B
FB5E
FB62
FB37
FB3B
FB6B
FB71
FB41
FB33
FB69
FB8D
FB67
FB50
FBAC
FC0B
FB99
FA8E
FA85
FCD4
00C4
041F
0568
051B
04AC
04D1
0527
052C
04EF
04BF
04AB
0492
047F
049F
04EA
052A
0546
0555
0552
0516
04A9
0467
0489
04C1
049E
043A
0426
048D
04DE
04A3
0458
04C6
058A
04F0
01DB
FD7A
FA61
F9E8
FAF6
FB9D
FB45
FACA
FAE2
FB42
FB54
FB26
FB27
FB5C
FB6A
FB46
FB46
FB7E
FB81
FB17
FAA6
FAA4
FAEC
FB1D
FB3B
FB83
FBD0
FBBA
FB5C
FB57
FBCE
FBEC
FB2F
FABC
FC72
0066
0447
05D7
0550
04AB
04F3
0568
051D
046D
044C
04C6
050D
04CA
0491
04D9
053B
0520
04AF
047A
049C
04C2
04D7
0505
0534
050F
04A6
047A
04B8
04D4
045C
03E1
0441
0507
0467
0159
FD32
FA6F
FA19
FB07
FB91
FB52
FAFB
FB0E
FB52
FB65
FB4A
FB38
FB32
FB1E
FB08
FB0B
FB15
FB0B
FB04
FB21
FB44
FB36
FB08
FB07
FB43
FB68
FB45
FB32
FB9A
FC29
FC0C
FB2B
FAD6
FC9F
0074
045E
0654
0617
0512
0498
04BD
04DB
04B5
04A5
04E4
0522
050A
04C3
04BD
050A
054F
0548
0518
04FB
04F8
04F1
04E5
04DB
04CE
04BD
04BE
04CC
04AC
0449
0415
048C
0533
0480
0179
FD42
FA57
FA02
FB16
FB96
FB01
FA64
FA8A
FAF9
FAEC
FA85
FA7B
FAF1
FB4E
FB40
FB2D
FB6C
FBA4
FB63
FAE4
FABF
FB08
FB47
FB37
FB12
FB15
FB33
FB56
FB95
FBD9
FBB2
FB11
FB02
FCE7
00A4
043A
05BC
054D
04A5
04E8
05A1
05DB
0574
050D
0504
051E
0519
0510
0523
0520
04D6
0473
0449
045C
047C
04A0
04D3
04F4
04D6
04A3
04BC
0519
052D
04AF
0436
0487
0536
04A4
01C7
FDA3
FA7F
F9A6
FA5B
FB0A
FAFF
FAAD
FAA0
FACB
FADD
FADC
FB08
FB56
FB74
FB47
FB17
FB30
FB7C
FBA8
FB8B
FB48
FB18
FB1A
FB48
FB78
FB65
FB09
FAD0
FB2E
FBD8
FBE9
FB1E
FABA
FC72
0059
0450
0612
058F
04AF
04E3
05B1
05DC
053E
04C4
04F7
0559
0543
04CD
0475
0458
043B
0429
046F
04F5
0531
04EC
049D
04A9
04D6
04C4
04A4
04D1
0510
04DF
046E
0483
0511
049A
01D2
FD9C
FA83
F9FA
FAEB
FB64
FAEB
FA71
FA8B
FAC4
FAA7
FA82
FACE
FB56
FB8C
FB66
FB53
FB6B
FB57
FB0E
FB0F
FB7C
FBB7
FB53
FAE1
FB1E
FBC1
FBD6
FB3B
FAE2
FB50
FBB3
FB36
FAC4
FC4C
0020
040D
05BC
0541
048A
04C6
055C
0562
0506
0507
0567
0578
04FD
0483
0489
04DA
051A
054F
0588
0563
049D
03C1
03AE
0465
04FB
04DB
0483
049F
04E9
04B0
0430
0461
052B
04D0
01F9
FDC2
FAD5
FA72
FB49
FB73
FABE
FA5C
FADB
FB7A
FB7A
FB2C
FB2C
FB51
FB18
FAA6
FA9D
FB10
FB5B
FB28
FAF0
FB2F
FB91
FB79
FB09
FAF0
FB4A
FB75
FB34
FB29
FBA8
FBEC
FB50
FAD9
FC65
0028
03F3
058D
051E
0497
04FC
057A
0524
047B
0478
04F9
051D
04C5
04B1
0523
0561
04DF
0435
0447
04E9
0528
04C7
048A
04E6
053C
04F1
0479
0491
04F3
04CF
0448
045D
0516
04C4
01F9
FDBD
FAC4
FA60
FB3A
FB6B
FAD9
FAB5
FB58
FBCB
FB5A
FA9E
FA84
FB07
FB6C
FB64
FB4D
FB5A
FB45
FAF0
FAC5
FB0F
FB6F
FB73
FB47
FB54
FB75
FB3D
FAE0
FB0F
FBC3
FBED
FB0B
FA79
FC36
0036
03FC
055D
04D8
0480
0525
05AA
0519
0426
0419
04EB
056B
0509
0488
04B1
0529
052E
04CB
04B2
0515
0565
0542
04F2
04D7
04D6
04AF
0482
0493
04B7
049A
047A
04E8
058C
04E5
01FE
FDFB
FB22
FA7C
FAFA
FB1F
FABD
FAA5
FB21
FB8B
FB66
FB19
FB34
FB8A
FB90
FB40
FB10
FB2C
FB46
FB2A
FB05
FB02
FAF7
FAC4
FAB2
FB08
FB79
FB78
FB22
FB24
FB91
FB8A
FAA7
FA32
FC08
002C
043E
05E2
0533
0446
0485
0555
0574
04D0
0461
04A8
0513
04FD
0490
046A
04B3
0505
050A
04DC
04C1
04CA
04E4
04FD
0509
04FC
04F4
0520
0561
054A
04BB
044F
04B0
0564
04E0
022D
FE43
FB42
FA4C
FAA2
FAF4
FAEF
FB0E
FB6D
FB81
FB0A
FA95
FAC0
FB58
FBA4
FB70
FB36
FB45
FB54
FB18
FAD8
FAF9
FB51
FB61
FB11
FAC9
FAC8
FAE3
FAFE
FB46
FBB1
FBA7
FADD
FA5B
FBD6
FF96
03AF
05D3
05AA
04C9
049D
0512
0554
0523
04EF
04EF
04DC
048B
0449
0458
0488
0499
04A5
04E0
0529
0542
0541
0563
0587
0550
04CC
048F
04DD
0527
04DA
0469
04B8
057F
0508
022D
FE11
FB22
FA85
FB2B
FB73
FB00
FA99
FABA
FB0B
FB28
FB39
FB7A
FBA9
FB6C
FAFF
FAF5
FB63
FBBC
FB95
FB22
FAD3
FAC2
FABA
FAAE
FABE
FAE0
FAE4
FAD9
FB05
FB52
FB30
FA83
FA5A
FC1C
FFC1
0377
0559
054B
04BC
04C3
0517
0505
04A6
04A6
0528
058F
0567
04F6
04B9
04B4
049A
0471
048B
04E8
051E
04FC
04D5
04F1
051A
050A
04EF
0513
053A
04FE
04AE
050F
05F3
05A5
02B5
FE1F
FABA
FA32
FB5C
FBFE
FB77
FAE2
FB09
FB5F
FB23
FA95
FA78
FAD4
FB0B
FAF1
FB03
FB6B
FB94
FB1E
FA98
FAB0
FB2C
FB59
FB29
FB27
FB6D
FB72
FB02
FAB2
FAF1
FB23
FA9F
FA3E
FBCD
FF96
0378
0529
04C3
0437
04A7
0559
054D
04C5
04B1
052D
0579
0532
04DC
04EB
0515
04EF
04B2
04D1
052B
0544
050F
04ED
04F2
04D1
0488
0492
0516
0563
04E2
0433
0485
059F
0581
02A4
FE24
FACF
FA2D
FB27
FBC1
FB60
FAE0
FAF2
FB3F
FB33
FAED
FAEA
FB27
FB35
FAF4
FAC0
FADD
FB16
FB26
FB1C
FB2B
FB3F
FB21
FAEA
FAEC
FB2E
FB54
FB39
FB24
FB37
FB07
FA5F
FA35
FC0D
0012
0443
0643
05C5
04A3
047F
051D
0559
04F6
04B2
04EC
051A
04C5
0459
047B
0502
0538
04F8
04D8
0522
0557
0504
0490
049A
0508
053D
050D
04D2
04BD
04A0
0486
04E1
058B
052C
0278
FE1F
FA97
F99B
FA76
FB3E
FB1F
FAB8
FAB4
FAEE
FB09
FB21
FB6B
FBA7
FB76
FB08
FAF4
FB53
FB99
FB67
FB09
FADC
FAC8
FAAF
FADB
FB75
FBEE
FBA0
FAE6
FAC5
FB68
FBB0
FADB
FA19
FB8A
FF8C
03EA
061F
05F1
051C
04F7
0546
053F
04DE
04B9
0501
0543
050E
048C
0435
043B
0478
04BB
04F2
050E
04F9
04C3
04A7
04C7
0500
0501
04A6
0447
0476
0544
05B4
046A
0116
FD25
FA9E
FA4C
FB2B
FBAB
FB49
FAB3
FA98
FADB
FAF7
FAD1
FABA
FAE1
FB1E
FB49
FB76
FBB2
FBD4
FBB7
FB85
FB87
FBB0
FB94
FAFE
FA6B
FA8E
FB54
FBC4
FB3A
FA90
FB8C
FEDD
0305
059E
05B6
0493
0409
047E
04F8
04C9
0474
04B3
0550
0581
0515
04AE
04C5
050D
0502
04B0
0489
04A4
049F
0450
041D
0460
04C5
04B7
0454
0468
0548
05FF
04F7
01A5
FD6B
FA98
FA53
FB91
FC47
FB9A
FA83
FA58
FB19
FB9D
FB3E
FAB2
FAF1
FBC5
FC1D
FB9F
FB17
FB2F
FB7D
FB54
FAF1
FB0E
FBA9
FBEE
FB91
FB47
FB9B
FBDB
FB17
FA02
FAB2
FE1F
028D
053B
054F
045A
0426
04D6
0564
053F
04D8
04D0
051A
053A
04F7
048A
043E
042B
0446
047E
04B6
04C9
04B1
048E
048D
04B9
04DF
04B6
044E
0434
04D3
058C
04E9
0216
FE19
FB1C
FA56
FAFF
FB7C
FB3B
FAFD
FB59
FBCE
FB94
FAD6
FA7B
FAE8
FB85
FBA2
FB4F
FB1D
FB48
FB81
FB7D
FB5F
FB65
FB82
FB80
FB71
FBA2
FC00
FBF6
FB2C
FA55
FAEB
FDBD
01CE
04F3
05CA
04FB
0450
04A7
054C
0546
04B7
0481
04E7
0536
04DE
044F
044A
04C9
050E
04D4
04A2
04DE
0515
04B8
0420
041A
04A8
04E7
0465
03EF
0476
056A
04F3
0210
FDFF
FB16
FA71
FB29
FBAF
FB6A
FAD7
FA92
FAAB
FAE3
FB1A
FB5B
FB92
FB92
FB5D
FB3D
FB5B
FB7F
FB62
FB2B
FB49
FBC8
FC0F
FBA1
FAE6
FACD
FB8C
FC19
FB76
FA4A
FA97
FD88
01E3
051C
05DD
0511
047F
04D0
0548
051F
0487
0449
04AD
0533
054B
04FC
04B7
04BD
04E6
04F0
04CE
049F
046C
0430
0409
0432
049D
04CF
047D
0426
0495
0595
0591
0322
FEE0
FB31
F9EE
FAA4
FB66
FB26
FA94
FAB1
FB5E
FBBB
FB7A
FB22
FB1C
FB24
FAE6
FAA3
FACE
FB4D
FB8E
FB64
FB48
FB92
FBE1
FBB0
FB3B
FB45
FBED
FC51
FBA6
FA82
FA99
FD06
00FB
045B
05AA
0540
0493
0491
04EE
04F9
04A6
0490
04FD
0570
0553
04C8
0479
04A3
04D4
04AE
0474
048D
04CF
04C1
046B
0457
04B5
04EE
0484
0403
045D
055C
054F
02D6
FEAE
FB2F
FA01
FAB1
FB96
FBAA
FB3F
FB19
FB66
FBAD
FB8C
FB2C
FAF2
FB05
FB3A
FB5D
FB64
FB62
FB66
FB6D
FB78
FB8C
FB92
FB5E
FB05
FAF5
FB73
FC08
FBDA
FAEC
FAA9
FCA5
00B4
04AC
0663
05C9
04A7
0475
04F9
0526
04B6
0457
0484
04E0
04D8
0479
0444
0467
0496
049C
04AC
04F4
0530
0506
049F
047F
04BD
04CE
0454
03D5
0426
0520
0548
033C
FF5D
FBBE
FA2D
FA92
FB5A
FB55
FAC1
FA86
FAE5
FB4C
FB45
FB0F
FB21
FB6E
FB85
FB44
FB10
FB3B
FB88
FB91
FB64
FB67
FBA8
FBBC
FB66
FB0F
FB3A
FBA9
FB91
FAD0
FA9A
FC67
0027
03F7
05DB
059C
04B3
0486
0516
057A
0544
04E4
04DB
0501
04E7
0496
0486
04E1
053D
0538
04FB
04D8
04BB
045B
03E5
03F1
04A0
0531
04EA
043B
044F
055A
05D5
0400
0001
FC04
FA1C
FA5E
FB32
FB3F
FAA4
FA5B
FAD6
FB89
FBB9
FB53
FAE4
FAD8
FB19
FB49
FB41
FB27
FB25
FB2E
FB29
FB20
FB28
FB2B
FB1A
FB27
FB8C
FBF1
FB9B
FA7B
F9EE
FBA8
FFBB
040D
0637
05E3
04C8
0482
04FD
0536
04E4
04AC
04F5
054A
051E
04AB
048F
04D1
04E1
0486
0448
04A4
053E
055C
04EC
049D
04D5
051E
04E2
0468
0493
0583
05EF
0447
0084
FC84
FA5E
FA7B
FB7B
FBCE
FB34
FA8F
FA90
FAF5
FB15
FAD1
FAAA
FAF1
FB5D
FB81
FB59
FB30
FB22
FB10
FAFD
FB1F
FB70
FB89
FB2E
FAD4
FB16
FBBA
FBC2
FAD2
FA2A
FB8E
FF32
032E
0555
0547
0476
0444
04B3
0500
04E6
04D5
0513
0548
0510
04A5
0495
04F9
055B
055A
0526
051D
0535
0518
04BB
0481
04A0
04C6
048D
0430
045F
0536
05A8
0452
0108
FD43
FAE7
FA91
FB48
FBB4
FB70
FB0D
FB10
FB4E
FB56
FB26
FB22
FB62
FB7F
FB2A
FAB0
FA98
FAE3
FB0D
FAD2
FAA4
FAFB
FB90
FBAE
FB46
FB14
FB7E
FBD2
FB44
FA75
FB38
FE70
02A9
0562
0596
0494
042D
04B9
053F
050D
048C
046D
04BD
0500
04F8
04D7
04CB
04C2
04B5
04CF
0518
0538
04E3
0465
045F
04E8
054D
04F3
043E
0438
0530
05F9
04E7
0195
FD7E
FABA
FA2A
FAF4
FBA7
FBA0
FB47
FB2A
FB3F
FB2A
FAE4
FAD2
FB2A
FB90
FB8D
FB2C
FAEA
FB0C
FB4B
FB4E
FB28
FB29
FB4F
FB4E
FB19
FB14
FB6B
FB96
FB04
FA46
FAF1
FDF4
0234
054F
05E9
04E1
041A
046D
0526
054E
04E9
04A7
04D3
050A
04EE
04AA
0496
04AD
04AD
0495
04A9
04F6
0521
04EE
04A0
049C
04C5
04A6
0443
0457
0549
062C
0551
0216
FDE6
FB06
FA77
FB38
FBA4
FB30
FA9B
FAAC
FB3D
FB9A
FB77
FB2E
FB22
FB47
FB51
FB35
FB25
FB35
FB3A
FB1B
FB06
FB2A
FB5D
FB4F
FB11
FB0E
FB63
FB88
FAF8
FA3F
FAD3
FD94
0196
04C2
05CF
0551
04BF
04CC
0502
04D9
0486
048B
04DF
04FB
04BB
049A
04F0
055A
0542
04BD
047B
04C8
051A
04E2
0469
046E
04FE
054E
04EB
0481
04EF
05C7
0558
0295
FE86
FB67
FA7B
FB0B
FB8F
FB64
FB0B
FB16
FB5B
FB52
FAE7
FA8A
FA99
FAF6
FB44
FB55
FB3E
FB1E
FAFC
FAE6
FAFF
FB44
FB74
FB55
FB11
FB14
FB71
FB98
FB00
FA24
FA83
FD2A
0149
04A5
05AB
04E5
0427
047A
0543
056D
04EE
04A1
04F3
0554
052C
04B5
0495
04D7
04F2
04B3
0497
04FB
0565
052B
0489
046C
0513
0591
0518
0446
0465
0568
057C
030B
FED0
FB46
FA17
FAA2
FB2E
FB02
FABC
FAFE
FB78
FB83
FB25
FAFA
FB44
FB98
FB7C
FB13
FAD6
FAEA
FB08
FB05
FB14
FB54
FB77
FB1C
FA7B
FA4A
FADB
FB8E
FB81
FAD6
FAEC
FD0A
00DB
0477
061C
05B1
049B
0432
049E
051F
052B
04EA
04C8
04D7
04D8
04AC
0488
04A8
0504
0558
0571
054F
0512
04DC
04CD
04F0
051A
04FE
048F
043A
0482
0530
051E
032B
FF8A
FBF1
FA2C
FA79
FB77
FBB5
FB19
FA99
FACD
FB4D
FB6B
FB29
FB0D
FB46
FB6E
FB3D
FAFD
FB0B
FB33
FAFB
FA7E
FA64
FAE3
FB55
FB1E
FAA7
FACF
FB8A
FBCA
FB23
FAE7
FCD8
00DC
04AE
062C
0579
046C
044E
04CC
04FC
04AC
046A
0494
04F3
0528
0519
04E0
04A3
0495
04DC
0540
0550
04FE
04D0
0521
057F
053A
0481
0447
04CE
04D2
02D7
FF26
FBCA
FA69
FAB0
FB2D
FB2A
FB04
FB25
FB53
FB43
FB25
FB3C
FB5F
FB38
FAF3
FB06
FB63
FB76
FB16
FADF
FB36
FB91
FB44
FAA9
FAAE
FB4D
FB70
FAB9
FAB1
FD23
018D
0533
061F
052A
048E
0511
059A
0533
0468
0444
04D0
052F
04F0
0483
046B
0494
04BB
04E3
051B
0524
04E2
04AE
04D4
04FA
04AB
0448
04AE
05AB
057C
02AD
FE32
FAC2
F9F8
FAD1
FB5B
FB0B
FABE
FAFA
FB37
FAF7
FAA5
FADD
FB6E
FBA7
FB6E
FB4A
FB6D
FB64
FAFA
FAB7
FB02
FB63
FB37
FACE
FAFA
FBA4
FBC1
FB15
FB29
FDA4
01E9
0556
0623
052B
0473
04B7
051E
0500
04C4
04FA
055F
0553
04DC
0492
04B7
04F1
04FA
04FE
0518
0504
04AC
0485
04E3
0550
0525
04AA
04BF
054F
04CB
01EF
FDAA
FA7B
F9CE
FAA5
FB30
FAF2
FABF
FB23
FB9E
FB8F
FB14
FABD
FACB
FB0C
FB4D
FB79
FB6D
FB1B
FAD7
FB07
FB71
FB61
FAC0
FA6D
FAFE
FBAE
FB58
FA6C
FAF2
FE22
028C
0575
05C6
04ED
04B8
0545
0590
053C
04E9
04FD
0517
04D8
0496
04C6
0529
0523
04B0
0473
04BD
051C
051B
04E6
04D3
04BE
0479
0474
0520
05C3
04B4
014A
FD1D
FA97
FA74
FB41
FB63
FADC
FAA4
FB00
FB48
FB0E
FAB7
FAC2
FB10
FB39
FB31
FB34
FB47
FB3A
FB1E
FB3B
FB7D
FB72
FB16
FB03
FB79
FBB3
FB02
FA3F
FB50
FEDA
0312
057D
0583
04B8
04A4
0529
0559
050B
04DE
050F
052B
04EB
04A7
04B6
04DB
04B8
047B
0498
04F4
0501
04A3
046D
04AA
04DF
04A9
048C
0522
05A7
0463
00D1
FCB5
FA68
FA60
FB10
FB19
FAB8
FACE
FB4A
FB69
FAFC
FAA9
FADD
FB3B
FB4D
FB38
FB5F
FBAA
FBAF
FB6E
FB52
FB72
FB66
FB18
FB0C
FB75
FB93
FAD1
FA27
FB80
FF56
03AF
0600
05D5
04E4
04BF
0540
056B
0512
04D1
04F4
051C
0505
04E6
04ED
04E7
04A6
046F
0491
04D0
04B2
0455
0454
04C1
04F1
04A1
048B
053D
05AA
0402
000B
FBE3
F9E4
FA40
FB36
FB6A
FB1D
FB12
FB35
FAFC
FA86
FA78
FAF4
FB63
FB5F
FB37
FB50
FB82
FB70
FB3F
FB54
FB95
FB81
FB1F
FB12
FB80
FB98
FAE8
FA9D
FC76
0073
0457
05F7
0570
0494
048E
04EE
04F3
04CB
04FD
055D
054F
04D7
0494
04C5
04F9
04D3
049C
04B0
04D6
04A3
044E
0469
04D9
04DE
045F
044F
051D
056E
0363
FF2A
FB40
F9E0
FAB3
FBA8
FB8B
FAF9
FAE2
FB2D
FB3F
FB1C
FB36
FB83
FB83
FB22
FAE5
FB19
FB65
FB64
FB3E
FB45
FB4A
FB02
FAC9
FB40
FC14
FC11
FB01
FAAA
FCF4
014C
04EB
05D9
04E5
0435
0497
0513
04DF
0480
04B7
0532
0526
04A1
046B
04C8
0519
04E7
0488
047D
04AD
04B6
04AC
04E3
051B
04C1
040E
0411
0500
0541
0315
FEEF
FB53
FA1C
FAB8
FB55
FB2C
FAE5
FB10
FB4F
FB31
FB05
FB3B
FB8A
FB63
FAF3
FAE2
FB48
FB7F
FB34
FAF2
FB43
FBC3
FBB9
FB4A
FB40
FB98
FB63
FA81
FA96
FD40
01B7
0538
0604
0513
0479
04DB
0545
0507
04B0
04E7
054D
052B
04A9
0483
04DE
051D
04E2
048F
048E
04A8
0485
045E
049F
050E
0507
049A
049A
0524
04DC
0267
FE69
FB23
FA1A
FAB3
FB55
FB4B
FB06
FAF3
FAF3
FAE8
FB15
FB89
FBBE
FB5E
FAE3
FAF3
FB65
FB7E
FB22
FAFC
FB62
FBB6
FB5B
FACF
FAFB
FBA5
FB9C
FABD
FAD2
FD84
01F8
0566
061A
050B
043D
046C
04D1
04C8
04A2
04CD
0506
04E4
0496
0492
04CE
04E4
04C5
04BF
04DF
04DF
04BA
04D9
054E
056D
04B9
03F0
043E
0548
04FF
0208
FDBB
FADB
FA94
FB84
FBD7
FB59
FB10
FB65
FBA9
FB54
FAD9
FAD8
FB2C
FB50
FB39
FB43
FB72
FB73
FB3A
FB1E
FB3B
FB39
FAFF
FB07
FB9D
FC09
FB69
FA57
FAC9
FDCF
01FC
04D1
0563
04DD
04A1
04C4
04AF
046F
0497
0521
0554
04E7
047F
04AE
0516
050E
04AF
0495
04D3
04E1
0494
046F
04B5
04D4
0458
03F0
0497
05B0
051A
01C2
FD5F
FAC6
FAD6
FBDC
FBFC
FB34
FAB6
FB00
FB72
FB7B
FB52
FB4B
FB41
FB02
FADA
FB18
FB71
FB6A
FB22
FB23
FB74
FB8B
FB40
FB2E
FBA9
FBE8
FB1A
FA24
FB25
FED8
0335
058A
055D
047D
0473
04ED
04E7
0466
044C
04D0
052F
04EE
0490
04AB
04F0
04C7
0455
0444
04B1
0509
04F6
04C9
04C4
04A1
043F
043E
051B
05D8
048E
00CD
FC9F
FA7D
FAAB
FB68
FB5C
FAEA
FAF9
FB6F
FB7D
FB03
FABD
FB0D
FB78
FB83
FB6F
FB9E
FBCD
FB8A
FB12
FB02
FB4A
FB45
FADC
FAD7
FB9B
FC3C
FBB3
FACD
FBAD
FF18
0322
0543
0527
048C
04C1
0552
054A
04D0
04B9
051A
0536
04C1
045D
0487
04CE
04A2
0447
0459
04BE
04D3
0484
0468
04B2
04C6
044B
0402
04AD
0563
0425
0077
FC70
FA83
FAD4
FB83
FB46
FAA8
FAAA
FB2B
FB54
FAFE
FAD0
FB18
FB5B
FB44
FB38
FB93
FBEC
FBB9
FB43
FB3E
FBA3
FBC5
FB77
FB5B
FBB8
FBCB
FAFB
FA67
FC04
0004
0415
05D7
0569
04C1
04FB
056A
052A
048E
0475
04E0
050D
04C0
0485
04B1
04DA
04B1
049C
04EE
051E
048C
03A8
037D
0425
049A
0455
0433
04F6
057F
03C0
FF9C
FB9E
FA30
FAED
FB93
FB0A
FA52
FA89
FB49
FB83
FB27
FB0F
FB7D
FBBE
FB5C
FAE2
FAF4
FB5B
FB8E
FB9F
FBEE
FC42
FC0C
FB76
FB57
FBD4
FBEB
FB0B
FA90
FC84
00D3
04D1
061C
052C
044E
04AA
0563
0565
04EC
04CE
0512
0512
04AF
0481
04CA
0507
04CA
0469
0451
0448
03FB
03C7
043A
04FB
050E
0459
0405
04B7
051B
0334
FF18
FB4E
FA02
FAB6
FB58
FAF9
FA75
FAAB
FB42
FB72
FB3B
FB26
FB48
FB39
FB00
FB29
FBC9
FC29
FBD2
FB52
FB6B
FBDF
FBE8
FB7E
FB5C
FBAB
FB9A
FAD4
FAB6
FCFA
0141
04F6
0613
0543
049E
04FD
0572
0522
0490
04A1
0532
055A
04CA
0433
0438
049A
04C6
04A9
0491
0494
048A
0477
047D
047E
044B
0424
0485
052F
04D8
026D
FE95
FB5C
FA2F
FA9E
FB37
FB36
FAE2
FAB0
FAB1
FAD6
FB2C
FB9E
FBCF
FB90
FB3B
FB44
FB8C
FB90
FB42
FB2E
FB98
FBFB
FBCF
FB65
FB61
FBA2
FB64
FAB9
FB15
FDBA
01D5
04F4
059A
04BB
044D
04EF
0598
055C
04A3
0469
04D6
052C
04E9
046A
0450
049E
04D7
04B3
0473
0462
046B
044E
0419
0435
04D1
055C
04B8
023D
FE98
FB7F
FA4D
FACC
FB8E
FB76
FABD
FA64
FAD0
FB65
FB73
FB1C
FAFB
FB39
FB69
FB4D
FB37
FB7C
FBD9
FBCE
FB72
FB68
FBE2
FC28
FB8A
FAAE
FB46
FE2E
0232
050D
059A
04C8
044D
04BF
054E
0520
0479
0446
04D1
0574
057D
0513
04DB
0502
0508
0496
041A
0431
04B4
04D5
044F
03EA
046E
053F
04A4
01B6
FDAB
FAD1
FA4E
FB30
FBC6
FB70
FADE
FAD1
FB2C
FB5A
FB31
FB0C
FB26
FB3E
FB09
FAB8
FAC1
FB32
FB87
FB5E
FB0E
FB42
FBF6
FC4C
FBA3
FAC0
FB5C
FE4F
0259
052C
05AD
04DD
0476
04FA
0585
0545
0492
0453
04B5
0511
04F3
04B7
04DA
052F
0523
04A9
0463
04B1
051C
04EC
043E
03FC
04A1
054D
0475
0189
FDB8
FAF8
FA45
FAF0
FB7B
FB26
FA73
FA53
FAEE
FB90
FB99
FB3F
FB19
FB45
FB52
FB06
FAC9
FB07
FB78
FB7A
FB19
FB17
FBBD
FC32
FB98
FAA0
FB31
FE3D
025E
0528
05A1
04F4
04B4
051A
0554
04FF
049E
04B3
0503
050D
04D2
04BF
04EF
0500
04B5
046C
0498
050D
051C
0485
03EC
0429
052D
05BF
0478
012E
FD4D
FABE
FA4C
FB15
FB9E
FB45
FAA3
FA87
FAF9
FB63
FB73
FB6D
FB85
FB77
FB03
FA8D
FAC1
FB99
FC33
FBE6
FB24
FAE4
FB4B
FB74
FACF
FA48
FB82
FEE7
02E8
0568
05B3
04E8
0483
04DF
053A
04F6
0469
0452
04D0
053B
0509
048A
0477
04F4
0557
0515
0487
0468
04C2
04DF
0468
0412
0497
054E
0480
0169
FD74
FAF3
FAB4
FB67
FB67
FA97
FA18
FA8E
FB63
FBB3
FB6D
FB28
FB34
FB4D
FB2B
FAFE
FB16
FB53
FB52
FB08
FAE8
FB49
FBDA
FBEA
FB57
FAFE
FC1B
FEFA
026D
04BC
0533
04B4
0498
0538
05C2
057C
04C2
0482
04EA
0539
04DF
0459
0471
0514
0563
04FB
048B
04CA
055A
0539
044E
03BF
0459
0526
0439
00F8
FD05
FAA6
FA88
FB67
FBBC
FB40
FAB7
FAAD
FAE0
FAE2
FAC4
FAE6
FB4D
FB87
FB49
FADC
FAC9
FB1D
FB57
FB1E
FAD2
FB0A
FBA8
FBCF
FB16
FA7C
FBAC
FF1E
0342
05D4
05FD
04E9
0445
048C
050B
0522
0507
052F
0581
057E
0508
0499
049A
04D6
04DA
04B2
04D8
0564
05B0
051F
0421
03E5
04D4
05AB
047F
00DD
FC89
F9EF
F9D5
FAF0
FB8C
FB46
FAE1
FAEC
FB0F
FAD2
FA71
FA85
FB06
FB46
FAF1
FA9C
FAF4
FBB2
FBDD
FB25
FA6B
FAA0
FB77
FBBE
FB11
FAB1
FC40
FFCE
0397
05B1
05C9
050F
04BD
04FD
0537
050F
04CA
04CB
0509
0535
053C
054E
0577
056A
04F1
0468
0473
051B
0595
052B
0449
041A
04EC
0565
03C4
FFF9
FBFE
F9F8
FA30
FB25
FB6A
FB04
FACC
FB19
FB66
FB36
FAC5
FAA4
FAEC
FB29
FB0B
FAD1
FAE5
FB3C
FB5E
FB18
FAD0
FAFE
FB72
FB77
FAE4
FABE
FC6E
0017
0406
0623
05F4
04EB
04A4
0535
058B
0515
0482
04AC
0558
058C
04F3
0452
0464
04E5
050F
04CB
04BC
0523
0558
04C3
03EB
03F7
0504
0590
03ED
002A
FC2A
F9E0
F9AA
FA75
FB10
FB27
FB0F
FB07
FAF8
FAC7
FAA3
FAD6
FB5A
FBCA
FBCD
FB76
FB26
FB0F
FB08
FAEF
FAFB
FB74
FC0A
FBFD
FB26
FAB0
FC33
FFE6
03FD
0634
05F5
04BD
0452
04F9
05A4
0586
04FC
04CF
051A
0540
04DF
0455
0439
0494
04EB
04F5
04E2
04ED
04EB
049B
043C
0463
050B
051C
0350
FFB8
FC07
FA20
FA51
FB42
FB89
FB05
FA90
FAB8
FB23
FB3F
FB0F
FB07
FB49
FB75
FB42
FAEE
FAE4
FB1D
FB38
FB1B
FB1F
FB7A
FBBB
FB4B
FA72
FA83
FCAC
008E
0448
0613
05C9
04C8
0467
04C3
0513
04E1
0492
04AD
0502
04F6
0479
043F
04CF
05B0
05EB
054A
049C
0497
04EA
04CF
044E
0443
04F9
0540
038F
FFE5
FC1D
FA26
FA3D
FB16
FB7D
FB62
FB55
FB87
FBA1
FB6F
FB2E
FB2D
FB5A
FB62
FB1F
FAC4
FA93
FA90
FA99
FAB1
FB06
FB9A
FBFC
FBB2
FAFC
FAFA
FCC8
003D
03BA
058B
0571
04A7
0463
04A7
04BA
0462
0435
049F
0532
0538
04B9
0470
04C0
0530
0527
04DA
04EE
056C
0593
04ED
0426
044A
053A
055E
0348
FF6A
FBE3
FA78
FAFD
FBDC
FBE9
FB64
FB38
FB9D
FBDC
FB60
FA9A
FA75
FB1B
FBB4
FB81
FACA
FA78
FAD7
FB4C
FB43
FAFF
FB10
FB56
FB20
FA77
FAA8
FCED
00C7
042C
0583
0512
044F
0426
045A
046A
046F
04C7
0544
0553
04D3
0464
04A2
0551
05A3
053F
04AB
0498
04FE
0539
04F3
04A8
04FB
059F
0544
02E2
FEFE
FB86
FA20
FABE
FBE1
FC38
FBBD
FB40
FB35
FB53
FB38
FB01
FB02
FB2A
FB1A
FACB
FAB5
FB1C
FB8D
FB5B
FAA0
FA40
FAC2
FB7E
FB66
FA93
FA9A
FCF0
0115
04BE
0606
0532
041E
0424
04E6
053D
04CF
0458
0485
050B
0531
04DF
04A1
04C5
04EA
04B7
0489
04EC
059B
05AF
04E6
0448
04DB
05FE
05AE
02C5
FE7A
FB3D
FA43
FAB0
FB0A
FAE8
FAE4
FB5B
FBCE
FBAB
FB1F
FAD2
FAFE
FB38
FB1A
FAD6
FAE0
FB42
FB7B
FB2D
FAA9
FA97
FB18
FB76
FB02
FA39
FAA5
FD59
018C
050F
064A
05A5
04C8
04B4
04FB
04DD
047B
048A
0520
0578
0511
0475
0484
0533
0597
0533
04A8
04C3
0544
0538
0474
040A
04DD
0613
059B
0263
FDC4
FA5F
F9A4
FABD
FBC9
FBD0
FB4B
FB0B
FB26
FB1D
FAC3
FA86
FAC7
FB3B
FB49
FAE4
FA9B
FAC8
FB12
FAFC
FAB8
FAEA
FB92
FBCB
FAFD
FA1B
FB03
FE63
02AD
0576
05D4
04ED
0465
04A7
04FD
04E2
04B0
04EF
0578
05A4
0537
04B4
04AE
0511
0553
0534
050B
053C
0590
0573
04D1
0465
04CE
056D
04AC
01B0
FD98
FAA6
FA0F
FAE9
FB77
FB21
FABF
FB0C
FB8E
FB5F
FA8F
FA21
FA9E
FB5D
FB6B
FAD7
FA78
FAB1
FAF6
FAC5
FA82
FADD
FBA1
FBCA
FAFD
FA5C
FB81
FEB2
0277
04FF
05B4
0558
04E8
04C1
04C3
04D3
04FD
0534
0544
0515
04DB
04E4
0532
0572
055B
0507
04D3
04E6
04FE
04D3
0489
049C
052A
0570
044C
015E
FDAD
FAED
FA10
FA99
FB3F
FB3B
FACF
FAB4
FB1C
FB8D
FB85
FB20
FAE2
FB08
FB46
FB3F
FB02
FAE5
FAFE
FB0E
FAF3
FAE3
FB04
FB09
FAAD
FA8A
FBE2
FF2D
031A
0591
05C1
04D4
0471
04E7
0543
04E2
044E
0452
04D2
0512
04D0
048A
04A8
04F0
04FF
04F5
0529
0573
0556
04DF
04C8
054D
0550
0356
FF6D
FB84
F99D
F9EC
FAFA
FB70
FB3C
FB0D
FB2B
FB4C
FB32
FB08
FB09
FB29
FB39
FB2E
FB1D
FB08
FAF1
FAFA
FB37
FB5E
FAFF
FA43
FA41
FC19
FFA5
034A
0560
05A5
052E
0502
052A
0527
04E0
04BE
04F1
0518
04D6
046F
0476
04FC
0574
056D
0516
04D4
04B5
049E
04C1
0556
05C7
04BE
0199
FD95
FAE4
FA7C
FB3E
FB79
FAD9
FA54
FA91
FB18
FB38
FB10
FB34
FBA1
FBBA
FB45
FACD
FAD0
FB0C
FB0F
FB0A
FB6D
FBE7
FB96
FA8D
FA71
FCCF
0103
0485
0587
04BC
0423
04A1
0566
0580
0516
04E1
0501
0500
04BD
04A0
04DF
0513
04E6
04AE
04DE
052A
04DA
0405
03C8
04BF
05B4
0497
00EC
FCAC
FA5E
FA8C
FB93
FBBC
FAFF
FA77
FABF
FB53
FB7F
FB42
FB0A
FB07
FB10
FB15
FB31
FB52
FB34
FADD
FAD1
FB55
FBD4
FB81
FAB9
FB1A
FDC8
01D4
04ED
05BB
050B
048B
04D5
0538
051D
04DA
04EF
0531
051F
04C5
04A4
04D1
04D3
047B
0459
04DE
057E
055A
04A1
0476
0522
0529
02F1
FEF9
FB9F
FA87
FAFB
FB39
FABF
FA7F
FB10
FBB2
FB78
FAAD
FA62
FAE2
FB66
FB57
FB1C
FB50
FBB5
FB9C
FB07
FABB
FB10
FB56
FAFB
FACA
FC50
FFD1
0392
0586
0568
04AC
04A1
051C
053A
04C7
046F
04AD
0526
0548
050F
04E6
04E8
04D4
0497
0484
04BF
04E5
04A8
0472
04E4
058F
04DF
01D7
FD96
FA89
F9F7
FAE2
FB85
FB53
FB0C
FB3A
FB79
FB48
FAED
FAF7
FB45
FB40
FADE
FAC5
FB36
FB89
FB33
FAC1
FB11
FBD5
FBC6
FAA9
FA45
FC86
00F4
04D4
060F
053A
0467
048E
04F6
04D3
047C
04B0
0550
0590
0527
04A9
049C
04C8
04BF
049D
04C6
0515
0502
0492
048B
0540
059D
040A
0060
FC77
FA65
FA7B
FB53
FB97
FB4A
FB24
FB55
FB5F
FAFE
FA98
FA9F
FAF6
FB38
FB5A
FB90
FBC3
FB96
FB10
FAD3
FB33
FB87
FB02
FA33
FAE5
FE13
0264
054F
05B9
04D7
046E
04D6
0528
04EB
04AC
04E6
0536
0510
04B6
04CB
0533
0525
0474
0402
0481
054A
0538
0471
0453
055A
05E1
03DA
FF7E
FB65
F9D1
FA75
FB57
FB3D
FAA4
FA7E
FAD7
FB1D
FB1C
FB20
FB46
FB48
FB0B
FAE9
FB21
FB67
FB5A
FB2C
FB5C
FBCD
FBB0
FAB4
F9FE
FB41
FED1
02F6
0583
05E1
053F
0500
055B
05A7
057F
0527
04F2
04D9
04B6
04A7
04D2
0504
04F3
04BA
04C1
04FD
04E2
044D
0410
04EC
0619
058E
0247
FDCA
FACB
FA60
FB2B
FB5C
FABB
FA49
FA7C
FAC4
FAB1
FAA9
FB19
FB8E
FB53
FAA7
FA86
FB2D
FBA9
FB40
FA99
FAC8
FB8D
FB96
FA9C
FA57
FC9B
00EC
04AE
05E1
050C
042A
0459
0519
058D
0593
057F
0564
0521
04D6
04D4
0514
0525
04D5
048A
04BD
0536
054C
04E5
04B8
0532
0577
0406
008F
FCB0
FA87
FAA3
FBA8
FBFC
FB66
FAC6
FAAF
FAD2
FAC1
FA9F
FABE
FB05
FB1B
FB04
FB14
FB47
FB2E
FABC
FA91
FB18
FB9F
FB32
FA57
FAFD
FE2E
0268
0504
0518
042E
0416
04D6
0547
0503
04CC
051F
0570
052A
04B4
04C4
0528
0519
0494
0475
0516
058C
04FB
040E
043C
0580
05CD
035C
FF05
FB83
FA8A
FB47
FBD8
FB7E
FAE7
FAD0
FB10
FB24
FB03
FB0C
FB4E
FB73
FB49
FB16
FB19
FB2D
FB13
FAFB
FB47
FBCE
FBCE
FAF6
FA55
FBA0
FF39
0358
059B
0571
046E
0443
04F1
0551
04E7
046E
0497
04FD
04DB
0451
0437
04CD
0558
0540
04E0
04CC
04D6
0481
041E
047C
0555
04ED
0204
FDC6
FADA
FA7E
FB5C
FB92
FAF4
FAAB
FB2E
FBAD
FB7A
FB12
FB2F
FB94
FB7C
FAF1
FAD3
FB69
FBCF
FB52
FAA1
FADA
FBC1
FBE8
FAEE
FA8A
FCAC
00E2
048D
05B4
04F6
044D
0498
0514
04F9
049D
04B1
0514
0519
04AD
0473
04B7
04EB
0497
0437
0490
0563
059B
04E1
044D
04D2
0584
0451
00A4
FC76
FA46
FA81
FB7C
FBBA
FB57
FB24
FB36
FB0E
FAB6
FACF
FB78
FBEA
FB99
FB0B
FB10
FB78
FB5E
FAA4
FA44
FAD5
FB80
FB2A
FA5B
FB09
FE33
0260
051A
0584
04D7
048C
04D2
0506
04EF
04E5
0506
04FC
04AC
0485
04D1
051D
04D1
0436
0437
0513
05D9
05A2
04DB
04B8
055E
0548
02FA
FF00
FB9F
FA7C
FB0E
FB99
FB4A
FAC1
FACD
FB41
FB6C
FB29
FAF8
FB1B
FB40
FB22
FB13
FB68
FBBF
FB6C
FA94
FA2E
FAB0
FB49
FB16
FABB
FBF8
FF69
035F
0588
056A
0496
0483
0505
052D
04DD
04C4
0516
0530
04B3
0433
0460
04F3
0518
04BB
04A3
0521
056D
04E6
0441
049C
058A
050A
01EC
FD99
FAC0
FA6C
FB3C
FB74
FAFE
FAD2
FB30
FB4F
FACB
FA61
FAD0
FBB0
FBF8
FB73
FAEF
FAFD
FB2F
FAFE
FAC5
FB2B
FBD8
FBB4
FAB2
FA87
FCE1
0122
04B6
05C5
0504
046F
04D8
0564
053B
04C2
04CE
054A
0568
04E9
047C
04AA
0506
04EE
048C
048E
04F5
0507
0488
044B
04EB
0560
03D4
000B
FC1F
FA5C
FACE
FB98
FB64
FAB2
FA9E
FB2C
FB7C
FB37
FAED
FB06
FB1D
FAD5
FA9A
FB03
FBB7
FBCC
FB2B
FACE
FB49
FBC9
FB45
FA66
FB33
FE93
02DA
0574
059F
04D8
04AF
051D
0535
04BF
046D
04A6
04FC
04EC
04AB
04B4
04F0
04E1
0489
047D
04F3
054A
04EA
0453
048D
058D
05AF
0362
FF20
FB42
F9B5
FA48
FB4C
FB8B
FB39
FB14
FB44
FB5D
FB2D
FB06
FB31
FB82
FBA0
FB88
FB6F
FB51
FB09
FAC0
FADE
FB5A
FB78
FACB
FA42
FB94
FF3F
0387
05FC
05E8
04CB
045D
04C7
0511
04CA
0482
04B3
04FF
04DA
0471
045F
04AF
04D3
0499
0486
04EB
0543
0502
04A3
0507
05CE
052B
01FE
FD9B
FAAD
FA5E
FB50
FB9E
FB11
FAC4
FB3C
FBBC
FB94
FB27
FB2D
FB8B
FB8E
FB1B
FAE1
FB3E
FB9F
FB70
FB08
FB14
FB59
FAF8
FA08
FA25
FCB9
0106
0498
05C3
0524
047C
049A
04F1
04E1
049E
04A1
04D7
04D0
0488
0472
04BB
04FC
04D4
0485
0491
04EB
0508
04CA
04CE
0570
05CA
0459
00C5
FCAF
FA42
FA28
FB29
FBC0
FB9C
FB5A
FB56
FB4D
FB16
FAFE
FB3B
FB74
FB40
FADE
FAE8
FB62
FBA6
FB57
FAFC
FB1D
FB50
FADA
FA39
FB1F
FE65
0293
0533
0569
0488
0436
04A4
04F5
04C9
049B
04CA
0504
04ED
04BB
04CA
04FD
0504
04EA
04E8
04F0
04D2
04C2
0511
054A
0433
0133
FD75
FAFD
FA95
FB2C
FB6B
FB2D
FB14
FB4B
FB6C
FB4A
FB26
FB2A
FB28
FB09
FAFF
FB1F
FB23
FAE9
FAD1
FB2A
FB72
FB07
FA99
FBE3
FF75
0377
0581
053A
0460
046D
0519
0558
04FE
04BA
04E1
050B
04ED
04CA
04D0
04C0
0489
049B
0513
0551
04F4
04A8
051D
0571
03CE
FFE2
FBD8
FA25
FACC
FBAF
FB6A
FAB2
FAB2
FB3C
FB66
FB1F
FB0B
FB49
FB51
FB02
FAE1
FB2F
FB72
FB43
FB02
FB22
FB40
FADB
FAC9
FCB8
00C2
0493
05E7
0514
0448
04A7
055C
0551
04BD
047F
04BB
04DE
04B3
04A4
04E0
0504
04E2
04D6
0503
04FA
04A2
04AE
0559
054D
02EF
FEB3
FB1A
FA11
FAF3
FBB5
FB71
FAF8
FB17
FB67
FB41
FADF
FAD6
FB18
FB37
FB31
FB48
FB5E
FB2C
FAF1
FB2A
FB96
FB5A
FA81
FAB4
FD6F
01D0
051E
05C9
04F0
0488
04EC
0524
04C6
0473
04A2
04FE
0518
050C
0510
04F8
049E
0465
04B7
0528
04F3
045D
0483
055F
0518
0234
FDD6
FABD
FA3A
FB16
FB80
FB23
FAD2
FAFC
FB38
FB38
FB35
FB4F
FB3E
FAFB
FB03
FB74
FBA6
FB3C
FAE9
FB57
FBE1
FB71
FA88
FB38
FE94
02E9
056F
0565
0488
0483
0517
0538
04E0
04C3
04F5
04F1
04A8
0499
04D7
04D9
0476
0447
04B0
0514
04C7
0453
04BB
056F
045A
00A5
FC55
FA30
FA9C
FBA5
FBB9
FB2D
FAFF
FB33
FB28
FAD9
FAD9
FB3E
FB73
FB42
FB35
FB8D
FBBB
FB61
FB17
FB5C
FB8D
FAF0
FA6C
FBF6
FFF4
042E
0613
0581
0485
048C
050A
04FB
0491
0499
050B
053B
04FE
04C3
04B5
0491
045D
047C
04E5
04F8
0488
046B
0531
05A0
03BB
FF81
FB88
FA1F
FACB
FB60
FAF5
FA79
FAC9
FB68
FB7A
FB1A
FAFA
FB30
FB40
FB14
FB28
FB83
FB8A
FB1A
FAEE
FB59
FB83
FAE0
FAAD
FCC0
00EB
04AB
05E5
0522
047B
04E0
056E
0544
04C8
04BA
04F4
04EF
04C1
04D4
0504
04EB
04AC
04C1
0511
0508
04AE
04C9
0574
0538
029A
FE55
FB07
FA44
FAFD
FB54
FAF5
FACB
FB27
FB64
FB29
FAF2
FB1F
FB56
FB2D
FAF2
FB1C
FB66
FB3C
FAD8
FB02
FB94
FB78
FAAA
FB00
FDF5
024F
053B
0589
04AC
047C
0507
0537
04CD
0498
04F6
0544
0505
04B2
04C5
04E1
049D
045E
04A1
04FB
04C2
045A
04B0
0565
04A2
0160
FD31
FABC
FABA
FB79
FB69
FAE0
FAE7
FB5E
FB6F
FB10
FAED
FB27
FB38
FAFD
FAFD
FB68
FBA2
FB45
FAED
FB46
FBBB
FB42
FA7D
FB93
FF53
0398
05A1
0535
045C
0476
04F8
04F0
0496
04A5
0506
050F
04BE
04BB
0516
0516
0487
043F
04B1
050D
04A5
0442
04DD
058C
0424
0026
FBE7
FA0D
FAA6
FB96
FB88
FB22
FB4E
FBA4
FB63
FADC
FADC
FB48
FB5A
FB00
FAE7
FB48
FB87
FB45
FB07
FB3F
FB64
FAE1
FAA1
FC6E
006F
045D
05F4
0568
049C
049B
04DE
04C4
048B
04AA
04F5
04FE
04D6
04D9
0504
04FB
04C8
04CE
04F5
04B7
0439
0470
0571
058E
0322
FEE3
FB6D
FA69
FB05
FB75
FB34
FB04
FB4E
FB87
FB4A
FB08
FB24
FB42
FB01
FAC0
FAF3
FB41
FB1E
FADF
FB3F
FBF7
FBDB
FAC6
FA91
FD0E
0174
04DF
0591
04B2
0455
04E3
0548
04F5
0482
0481
04BE
04D9
04E7
050F
051A
04D5
0498
04C4
04FB
04A2
0418
046C
0574
053B
0250
FDF7
FAFB
FA9A
FB7B
FBC5
FB3D
FADA
FB09
FB49
FB39
FB24
FB42
FB3F
FAF8
FAE0
FB36
FB74
FB30
FAF2
FB5D
FBE9
FB88
FA9E
FB28
FE5C
02BB
0574
0585
0483
043D
04B1
04E2
04AC
04AA
04F7
050B
04C6
04A1
04D3
04F6
04CA
04B2
04FF
0536
04CB
0449
04A6
055A
0464
00E0
FCAA
FA6D
FAA3
FB7F
FB85
FB0D
FB0B
FB6A
FB67
FAF4
FACB
FB2E
FB82
FB59
FB1B
FB2D
FB42
FB11
FB06
FB74
FBB7
FB25
FA9F
FC05
FFC5
03D8
05CA
0564
0482
0481
04EC
04DA
047A
0487
04F4
051C
04E0
04B4
04C3
04CA
04BB
04DD
051F
0501
0475
0450
0509
056A
038F
FF78
FB8E
FA07
FA92
FB4E
FB4B
FB16
FB40
FB7E
FB66
FB32
FB3C
FB50
FB1A
FAE0
FB26
FBAB
FBA8
FB1E
FAF6
FB6F
FB85
FABB
FA89
FCD0
0122
04D1
05E9
0528
0492
04DB
0526
04DA
0489
04BE
0506
04D6
048A
04B6
0516
0504
0495
0468
048D
0481
044D
04A4
057E
054E
029A
FE3A
FADF
FA25
FB00
FB84
FB36
FAE7
FB05
FB32
FB36
FB53
FB92
FB8C
FB22
FADD
FB22
FB7D
FB59
FB10
FB61
FBF7
FBA7
FA90
FAC2
FDC6
024E
056B
05D9
04FB
04A1
04F7
051A
04D1
04BB
0503
050E
049A
0448
048F
04F9
04F8
04CC
04E2
04ED
0481
0422
04A8
0584
04C5
016B
FD11
FA65
FA3D
FB0C
FB3F
FAF7
FB09
FB61
FB5B
FB02
FAF7
FB4D
FB76
FB42
FB25
FB5C
FB78
FB2E
FB02
FB6F
FBD6
FB4D
FA7F
FB83
FF28
0379
05CA
05AB
04D7
04AD
04E7
04D0
0494
04C4
0535
0538
04C1
047E
04B3
04D9
04A2
0484
04C2
04D5
046C
0448
0512
05B3
042E
0038
FC15
FA36
FA9B
FB50
FB25
FAC0
FAFB
FB6D
FB4B
FACC
FABB
FB28
FB72
FB62
FB5C
FB85
FB83
FB3E
FB32
FB88
FB8B
FAC8
FA66
FC3B
004D
043B
05CD
054C
04A0
04C4
0528
0526
04FA
050A
052B
0506
04CC
04DC
0505
04C9
044A
0435
0494
04AF
045B
047B
0561
0594
0355
FF20
FB83
FA53
FADD
FB45
FAEF
FAA7
FAEE
FB2C
FAE8
FA9E
FADC
FB44
FB3D
FAFC
FB16
FB74
FB8E
FB6E
FB9F
FC02
FBBB
FABD
FAA8
FD21
0172
04DE
05AD
04E6
0492
0529
05A9
0577
0515
0511
053A
052A
04F2
04D5
04D0
04BD
04C0
04F9
0508
0483
03EC
0438
0520
04C7
01EE
FDD2
FAFC
FA7C
FB23
FB69
FB1D
FAF0
FB0F
FB03
FAAA
FA7D
FAB9
FAFA
FAF8
FAFE
FB38
FB47
FAF9
FAE0
FB69
FBE9
FB7E
FAC0
FB93
FED9
02FB
057D
05A6
04E9
04B8
04F9
04EE
04A6
04B7
0521
055B
053A
0515
0511
04F6
04C1
04C4
0506
0502
0482
043E
04DE
057D
0433
0085
FC6B
FA46
FA5F
FB1F
FB46
FB08
FB0A
FB41
FB3D
FAF9
FAD5
FAEB
FAFC
FAF4
FB09
FB33
FB22
FAE7
FB03
FB7D
FB89
FACF
FA81
FC3F
FFFC
03B1
057A
0569
04ED
04E8
0513
050B
050C
054A
0561
04FA
047E
0484
04E8
050D
04E2
04E7
0530
0526
0497
0455
0508
05A9
043C
0055
FC12
F9F4
FA3F
FB29
FB41
FACC
FAAA
FAEF
FB08
FAD2
FAC1
FB04
FB36
FB12
FAF3
FB2D
FB6A
FB34
FADB
FB17
FBC2
FBBC
FA8C
F9A0
FB0F
FF11
0368
0599
056B
04A5
04B5
054E
0571
0506
04CA
0511
0556
0524
04D4
04E6
052A
0511
04A2
048A
04FC
053F
04C1
0428
048B
0598
0568
02A0
FE4D
FAFF
FA1F
FAD2
FB6E
FB5B
FB1E
FB17
FAFB
FA98
FA5C
FAAF
FB3E
FB66
FB25
FB0C
FB51
FB75
FB1C
FAC3
FB16
FBD2
FBE8
FB02
FA76
FC08
FFD5
03DE
05EF
05B0
04A4
044E
04D5
0564
0572
053E
052A
0523
04EB
049B
0489
04BF
04F1
0501
051C
0546
051D
0482
041E
04A7
057D
04C5
0178
FD08
FA35
FA27
FB5F
FBC1
FB04
FA74
FACD
FB55
FB32
FABE
FADE
FB87
FBCC
FB4C
FAC5
FAE0
FB37
FB17
FAB5
FAD0
FB56
FB5E
FAC6
FB08
FD9A
01D3
0535
060E
051D
044F
0477
04E7
04F2
04D6
0509
0555
0535
04C2
049A
04E8
051E
04D7
0483
04BF
054D
055D
04CF
0484
0501
053F
038A
FFB4
FBB8
F9DD
FA6D
FBAB
FBF6
FB59
FAE6
FB0B
FB39
FAF3
FA8E
FA9C
FB10
FB66
FB6A
FB5B
FB5A
FB2A
FAC9
FAB8
FB44
FBC2
FB5E
FAA3
FB70
FECD
0341
0610
061C
04DE
0461
04EE
054B
04D6
0459
04AF
056E
0595
04FE
0478
048B
04DE
04F5
04ED
050A
050C
049B
041F
0467
0537
04EC
0241
FE1A
FADA
F9EF
FA93
FB21
FB09
FAEA
FB38
FB85
FB54
FAEC
FAE1
FB2B
FB42
FAFD
FAD3
FB12
FB5B
FB40
FB04
FB3B
FBC6
FBD1
FB1C
FADE
FCAC
007F
0458
0623
05B7
04AA
0464
04DA
0527
04ED
04A2
04B0
04E6
04E9
04D0
04F1
053C
0543
04ED
04A8
04BC
04D1
0483
0429
046F
04F8
0433
010F
FCBD
F9DC
F9CA
FB4B
FC26
FBA5
FAD9
FACD
FB40
FB64
FB28
FB1C
FB5C
FB5F
FAEC
FA8A
FAB3
FB1C
FB3E
FB3A
FB86
FBEC
FBB0
FAF9
FB50
FE01
022E
055B
0600
0505
044F
048B
04F1
04DE
04AE
04E1
0531
050A
048E
046E
04DB
0537
050F
04C2
04D5
0502
04B1
0419
0430
0515
0548
0329
FF16
FB62
F9FE
FA95
FB5B
FB43
FAD3
FADF
FB4A
FB64
FB0F
FADC
FB1A
FB63
FB4A
FB09
FB16
FB5C
FB5D
FB14
FB1D
FBAB
FBF8
FB50
FA88
FB8D
FF20
038C
062F
0628
04F5
0472
04E1
0541
0501
04A0
04B3
0507
0517
04EA
04E2
0507
04FF
04B6
0490
04B6
04B8
0446
03F4
0489
0588
052E
0251
FE04
FAB4
F9C3
FA74
FB2E
FB44
FB1F
FB26
FB2D
FB01
FADD
FB0A
FB54
FB52
FB0D
FAF3
FB24
FB47
FB2E
FB39
FBB8
FC26
FBB4
FA9C
FA72
FC97
0084
0418
05A8
056D
04D1
04BE
04FE
0510
04FB
0511
0546
053C
04E6
04AE
04D5
050F
04F4
04A6
0491
04B3
0495
0421
040A
04CB
0582
0471
0107
FCEF
FA90
FA9C
FB90
FBB0
FAE5
FA56
FA9E
FB23
FB29
FAE0
FAE8
FB4B
FB79
FB3E
FB10
FB44
FB7D
FB51
FB0A
FB38
FBA5
FB82
FADC
FB29
FDBE
01E0
0520
05D8
04CD
03FF
0451
0502
0529
04E2
04D6
0519
0530
04F2
04C0
04D5
04E3
04AB
047B
04B6
050C
04E0
0459
0462
053B
058D
03A6
FF9D
FBA5
F9E1
FA5B
FB66
FBB6
FB70
FB47
FB50
FB24
FACA
FABA
FB19
FB6D
FB57
FB22
FB3F
FB7C
FB52
FAD8
FAC7
FB56
FBA6
FAFA
FA2C
FB32
FEC7
0332
05DE
05F6
04E5
045F
04A5
04E8
04CA
04C0
0515
055B
051D
04A4
0487
04CA
04E6
04B0
0499
04E5
0521
04DE
048C
04F6
05C4
054F
0275
FE3C
FB0F
FA4A
FB0C
FB90
FB32
FAAD
FAB4
FB10
FB31
FB12
FB16
FB4D
FB59
FB1B
FAEB
FB0D
FB41
FB2F
FB06
FB29
FB6C
FB28
FA62
FA63
FC87
0079
041E
059F
052D
047A
04B0
0563
058D
0500
0470
0461
0496
04A6
04A7
04E6
054D
0574
053F
0505
04FD
04EC
04AF
04A8
052C
058B
0454
0100
FCFA
FA76
FA3E
FB16
FB62
FAEB
FAA4
FB16
FBB3
FBC7
FB6E
FB38
FB3D
FB17
FAB0
FA76
FAAE
FAFF
FB05
FAFD
FB4A
FB9C
FB3E
FA72
FAD0
FD90
01C9
0509
05D8
0517
049A
04EE
0532
04BF
0421
042D
04C5
0525
0514
0513
0564
058D
052B
04B0
04BA
0510
04EA
0450
0443
052B
05AA
03DB
FFC6
FBC5
FA1F
FAB9
FB9E
FB80
FAE5
FADF
FB6E
FBB3
FB51
FAD4
FAC1
FAE2
FAD5
FAC5
FB0E
FB7E
FB80
FB11
FAE6
FB5A
FBB2
FB2A
FA77
FB6F
FED2
0309
059A
05B8
04C4
0463
04C3
0509
04D9
04B4
04F6
053F
0524
04E2
04EA
0516
04E3
0464
044B
04D3
053F
04E3
044A
048B
056E
0522
0255
FE11
FAE4
FA32
FB02
FB8D
FB46
FAE6
FAF8
FB22
FAF5
FAB3
FAD3
FB32
FB52
FB31
FB49
FBB4
FBDA
FB5C
FACB
FAF3
FB95
FB99
FABA
FA6B
FC69
0080
0462
05F4
0555
0459
045B
0513
057E
0543
04E1
04C6
04DB
04E5
04EB
04FB
04E6
048D
0447
0480
0503
0516
048E
043E
04DB
0593
0489
0109
FCCB
FA5D
FA80
FB92
FBBC
FAF4
FA79
FADE
FB69
FB58
FAF6
FAF7
FB4F
FB5C
FAFF
FAD8
FB38
FB92
FB5C
FAFE
FB2F
FBB1
FB8C
FAC7
FB04
FDAE
01E2
0508
05A4
04C9
0473
0514
0588
0511
0463
0476
0518
0552
04DD
046C
0489
04D7
04D0
04A1
04C8
0518
04F4
0467
0450
0502
0542
0368
FF85
FBB5
FA08
FA75
FB4C
FB55
FAE9
FAE6
FB5A
FB9A
FB5A
FB01
FAF5
FB12
FB16
FB20
FB63
FB9B
FB5A
FAD3
FACA
FB74
FBEB
FB64
FAAF
FBB7
FF38
037D
05FF
05FE
04F8
0492
04DC
04E5
0471
0437
04A1
051B
0503
04A9
04C1
053B
0556
04D8
046B
0495
04DA
0492
041D
0472
0559
0507
022A
FDD8
FAAD
FA07
FAD7
FB48
FAEF
FAB8
FB2A
FBA9
FB82
FB02
FAEF
FB5B
FB99
FB4C
FADD
FACB
FAFB
FB16
FB34
FBA1
FC1F
FBF4
FB19
FADD
FCB9
0087
044B
060F
05B7
04C9
049B
0519
055B
04FF
0489
0490
04FA
0534
04F8
048F
0465
0498
04F8
053F
0532
04C0
0436
0423
04B0
0505
03C1
0078
FC8E
FA24
FA0F
FB1C
FB93
FB0D
FA80
FABD
FB69
FBAA
FB53
FAF4
FAF8
FB2B
FB36
FB21
FB1D
FB2D
FB3F
FB72
FBC9
FBD3
FB2C
FA72
FB33
FE43
026F
055C
05E5
0516
04AC
051A
057C
0534
04B6
04B1
0503
050A
04AE
047B
04BD
050A
04F9
04C0
04C8
04E3
048F
03F7
03FD
04DF
0550
039D
FFBF
FBC8
F9E1
FA30
FB14
FB35
FAC8
FAB9
FB2D
FB71
FB20
FABB
FAE1
FB5F
FB7D
FB0E
FAC1
FB22
FBCB
FBDF
FB42
FAC8
FB17
FBB7
FBB7
FB1F
FB3E
FD4D
00E6
043A
05C0
0580
04B9
0475
04BE
050A
050C
04F0
04F4
050D
0509
04DC
04B1
04A2
04A2
049C
04A7
04DD
051B
0508
048C
0422
045B
04FB
04D0
02C4
FF31
FBE0
FA6C
FAC9
FB8F
FB92
FAF9
FAA3
FAE8
FB49
FB48
FB10
FB10
FB4A
FB56
FB1A
FAF6
FB37
FB90
FB7D
FB0B
FADD
FB4F
FBD4
FB9D
FAD6
FAE0
FCFA
00C2
0444
05BE
0536
0443
0445
0512
058C
052C
0491
048C
0503
052E
04C4
0462
04A3
0535
054B
04CE
047B
04C9
0524
04CB
0415
041E
050C
0552
0344
FF39
FB89
FA2D
FAD8
FBB3
FB94
FAF1
FABD
FB11
FB47
FB12
FADE
FB11
FB68
FB61
FB02
FAD0
FB0E
FB5C
FB4F
FB15
FB30
FBAD
FBE4
FB50
FA7F
FAD7
FD3B
00FB
0446
05B8
057C
04D7
04C3
0523
0546
04F4
04A3
04C2
051C
0535
04F9
04D0
04F3
050F
04C8
0457
044E
04BB
04FB
04A2
0438
0493
0575
0553
02E3
FEC1
FB23
F9CC
FA78
FB76
FB89
FAE9
FA8B
FAD5
FB4E
FB5C
FAF9
FA98
FA89
FABC
FAFE
FB44
FB8E
FBB5
FB93
FB49
FB39
FB83
FBB0
FB3F
FA8F
FAF4
FD74
0169
04C6
05F6
0559
049D
04D6
0582
0596
04FB
048F
04D8
055A
0560
0500
04D5
0501
04FA
0475
03FE
0440
04F8
0537
04B0
043D
04B4
0581
04FF
0247
FE56
FB33
FA0F
FA70
FB0B
FB18
FAC2
FA91
FAB8
FB00
FB26
FB25
FB27
FB45
FB64
FB64
FB50
FB4E
FB5F
FB52
FB15
FAE7
FB09
FB50
FB4B
FB0E
FB90
FDCA
016F
04C8
0637
05BC
04C5
0494
051E
058B
0567
0506
04D2
04BE
048C
0457
046F
04D2
0514
04FA
04CE
04F0
0533
050D
0473
041B
0499
0554
04C5
0214
FE38
FB3B
FA54
FAE9
FB7A
FB43
FABA
FA9A
FAE7
FB18
FAF8
FAE9
FB3B
FBA4
FB9F
FB29
FAC8
FADB
FB26
FB45
FB3E
FB68
FBB9
FBA2
FAE3
FA47
FB2C
FE10
01D8
04A9
058D
051C
049B
04AE
04FC
0500
04C3
04B4
04FD
0543
052B
04D9
04B6
04DE
04FF
04DA
04A8
04C0
0501
04F3
0488
0465
0505
05B9
04F8
01FA
FDE0
FADB
FA27
FB04
FBC6
FB96
FB01
FAE1
FB41
FB82
FB4F
FB01
FB0B
FB49
FB41
FADD
FA9E
FAE7
FB67
FB7E
FB1C
FADD
FB1E
FB5F
FAFA
FA61
FB1D
FE21
0255
055A
05DD
04CD
0416
047D
052D
0531
04BA
049C
04FE
0537
04E0
0479
04AA
053B
0568
04FD
04A7
04E9
0551
0511
044B
0414
04FA
05E5
04F3
018D
FD45
FA7A
FA2C
FB4F
FC20
FBD8
FB11
FAB2
FAE2
FB17
FAF0
FAAC
FAB7
FB0B
FB43
FB33
FB19
FB2C
FB33
FAE5
FA82
FAA2
FB49
FB9D
FB03
FA58
FB6C
FEF1
0346
05D7
05B0
0453
03D5
04A5
0581
0560
04AF
047D
04FE
0567
0527
04AC
04B2
0532
0570
0513
049E
04B3
052D
055D
050A
04C3
04FF
052A
0407
0119
FD6D
FAC0
F9F7
FA80
FB26
FB43
FB0B
FAF3
FB10
FB27
FB1C
FB13
FB2B
FB4E
FB4F
FB2B
FB09
FAF5
FAD9
FAB4
FAC0
FB2A
FBA7
FB9B
FAE4
FA68
FB83
FEA7
02A0
0574
0623
0567
04BB
04CE
0527
051C
04BA
0491
04D1
050F
04F2
04B1
04B7
04F5
0500
04C0
04A7
04FB
054C
04F4
0426
03EA
04C2
059D
04A3
0148
FD2A
FAA1
FA7E
FB7A
FBDA
FB38
FA8B
FAA6
FB3D
FB7C
FB33
FAF6
FB30
FB89
FB6C
FAEF
FABF
FB2F
FBB5
FBA6
FB26
FAF5
FB59
FBA1
FB28
FA94
FB79
FE93
029A
054D
059F
0494
03F5
046C
0539
056E
050C
04B4
04B9
04D4
04BD
049B
04B3
04E5
04CF
0470
043F
0488
04F0
04EB
0496
04AD
0574
05E8
048B
011C
FD2E
FAD2
FA9F
FB64
FBA8
FB2B
FABC
FAEB
FB56
FB60
FB16
FB04
FB58
FB95
FB59
FAFC
FB1C
FBB0
FBFA
FB88
FADE
FACD
FB47
FB5E
FAA3
FA1F
FB7C
FF13
0331
0597
0599
048F
042A
04BE
054E
0510
0465
0433
04AF
0528
0507
048B
0459
049A
04D7
04B8
0482
04A3
04FD
050F
04CA
04C1
0544
0588
0431
00E3
FCFB
FA74
FA13
FAE9
FB8B
FB7B
FB3A
FB45
FB71
FB56
FB06
FAF2
FB44
FB9E
FB9C
FB5E
FB4B
FB77
FB7E
FB28
FAD2
FAF6
FB64
FB5D
FAB0
FA6A
FBFB
FF8C
0378
05BB
05C8
04D8
0463
04B3
050D
04EF
04A7
04AC
04E4
04D3
046D
0433
047C
04EE
04F7
049E
047B
04DD
0548
0521
049A
0485
051B
054A
03AB
002A
FC69
FA54
FA5C
FB47
FBAB
FB43
FACD
FADC
FB39
FB5F
FB42
FB3F
FB77
FB98
FB5F
FB10
FB1D
FB75
FB8A
FB1A
FAA6
FACD
FB62
FB91
FB16
FAFA
FC99
0001
0394
0588
0590
04D9
0492
04D0
04F6
04C8
04A7
04DC
0518
04E9
046C
0434
0480
04DF
04CD
0469
0455
04CF
054B
052F
04B1
04A2
0534
0553
0398
FFF1
FC14
FA00
FA27
FB37
FBAE
FB49
FAD5
FAE7
FB35
FB37
FAFA
FAFD
FB63
FBB6
FB97
FB4B
FB4D
FB8F
FB8E
FB1F
FACB
FB12
FB8E
FB5F
FA82
FA55
FC4A
0032
0417
0608
05D6
04EC
04A2
0509
054F
0505
0491
0480
04C6
04E8
04B4
047D
0495
04D4
04D8
049E
0488
04C3
04F3
04BD
0476
04CF
05AA
05B5
0399
FFA6
FBD8
FA0C
FA4D
FB1A
FB34
FABF
FA92
FAF0
FB58
FB5C
FB35
FB49
FB84
FB82
FB37
FB0B
FB3F
FB81
FB5F
FB02
FB04
FB8A
FBDF
FB4B
FA40
FA45
FC88
0076
0415
05BE
0580
04BB
0497
0509
0559
0533
04F4
04F8
050D
04CD
044E
041D
0475
04DF
04D6
0482
047E
04E8
0521
04B2
0425
046C
0567
0589
0363
FF66
FBBD
FA3A
FABA
FB9C
FBA5
FB09
FAAE
FAE7
FB36
FB25
FAE8
FAFB
FB67
FBB5
FB94
FB41
FB2A
FB53
FB63
FB38
FB27
FB6F
FBA9
FB3C
FA6E
FA9D
FCF8
00F7
047C
05C6
0514
0429
044B
051F
057E
050D
0480
0484
04E3
04FD
04BA
0495
04CA
04F0
04A3
0434
044B
04E7
053E
04CD
0431
046F
0569
0582
0340
FF23
FB6E
FA05
FAB1
FBB0
FBBA
FB15
FAC1
FB0E
FB6C
FB5E
FB16
FB0A
FB40
FB5D
FB45
FB42
FB75
FB94
FB5A
FB0A
FB21
FB8A
FB8F
FAD2
FA1F
FAE0
FDA7
016A
045D
057C
0532
04A1
0482
04C2
04ED
04D4
04AB
04A9
04C2
04C7
04B5
04BD
04E9
0502
04D6
0493
0491
04C9
04C6
0458
0415
04AD
05B2
058E
0323
FF38
FBE9
FA99
FACF
FB29
FB01
FAC2
FAEA
FB47
FB6B
FB56
FB55
FB76
FB7E
FB5D
FB42
FB46
FB44
FB28
FB1F
FB45
FB61
FB3A
FB05
FB20
FB5F
FB39
FACE
FB49
FD9C
0124
040A
0522
04EF
04B0
04DB
04FB
04BE
047B
048D
04C5
04CD
04BB
04D0
04EF
04CE
0487
047C
04B9
04D1
049C
0487
04E2
052E
04CB
042B
0468
0572
0574
02D9
FE84
FB22
FA4B
FB13
FB9B
FB5A
FB22
FB75
FBC0
FB7D
FB18
FB36
FBA5
FBB4
FB4A
FAFD
FB1E
FB57
FB54
FB3C
FB4B
FB52
FB20
FB12
FB89
FC02
FB88
FA69
FA8F
FD61
01BD
04F2
059E
04D9
046E
04BA
04DE
0477
0427
046B
04D2
04CA
0489
049A
04ED
0507
04DE
04D6
04F9
04DA
0460
041F
0471
04C8
0482
0421
04B3
05DD
0597
028D
FE23
FB26
FAB6
FB6C
FB83
FAF3
FACE
FB5F
FBCB
FB85
FB10
FB0E
FB4F
FB4F
FB1E
FB21
FB4B
FB41
FB20
FB5B
FBDB
FBE9
FB4B
FAD6
FB3E
FBCB
FB40
FA09
FA60
FD9E
0234
0538
0591
04B9
0473
04DD
050F
04CE
04B6
0501
051D
04BA
0460
0490
04F3
04EF
04A6
04A8
04F4
0503
04BA
04A0
04E4
04E8
044D
03E4
04A9
05E1
0556
01FC
FD85
FAAA
FA45
FAF8
FB54
FB4C
FB70
FBAA
FB79
FAFC
FADA
FB33
FB6D
FB37
FB14
FB63
FBA2
FB38
FA93
FA9A
FB4C
FBB5
FB67
FB24
FB89
FBE5
FB3F
FA57
FB4E
FEEE
0337
0578
0544
0474
0489
0523
0531
04AE
0469
04AB
04E9
04C9
04A8
04D3
04F9
04CC
04A4
04EE
0555
053D
04C3
04A1
04F3
04F6
0457
03FE
04C3
05A9
0489
00CB
FC88
FA54
FA79
FB35
FB3C
FAED
FB13
FB7A
FB6F
FAFC
FADB
FB3C
FB7A
FB34
FAEF
FB2C
FB8B
FB64
FAE0
FABB
FB16
FB53
FB2A
FB24
FB95
FBCC
FB1C
FA6E
FBB7
FF7D
03BB
05EA
05AF
04CA
04AF
051F
0532
04D3
04A6
04DE
0508
04E1
04BA
04D1
04DF
04A6
047C
04C1
052E
0538
04EE
04DD
050E
04E8
0446
0406
04CF
058E
043E
006A
FC2C
FA07
FA46
FB25
FB35
FABF
FABD
FB44
FB9B
FB68
FB16
FB0F
FB2E
FB2E
FB22
FB31
FB36
FB0C
FAF1
FB28
FB73
FB69
FB35
FB63
FBE1
FBC9
FACA
FA40
FC0B
0021
0428
05DC
0561
049B
04B9
0537
052E
04B1
0474
04A5
04D1
04BF
04B8
04E1
04ED
04B4
0499
04E4
0533
0509
04A4
04A0
04E7
04C1
0415
03EC
04E8
05BD
0442
002A
FBE0
FA00
FA96
FB8F
FB70
FAC0
FAA9
FB3A
FB97
FB63
FB2C
FB64
FBB9
FBA2
FB30
FAD7
FACA
FAE3
FB09
FB35
FB42
FB26
FB31
FBAA
FC1F
FBB0
FA6E
F9F4
FBEC
FFF5
03BB
0568
055B
051B
0540
052C
0486
03FB
043D
04F4
053F
04F3
04AD
04C3
04D4
0491
0452
047B
04CC
04D2
04AF
04D4
0526
0519
04C0
04EB
05C2
05D2
0378
FF30
FB84
FA5F
FB17
FBAE
FB5B
FAFF
FB5B
FBE8
FBCA
FB23
FAC4
FAF6
FB34
FB28
FB21
FB63
FB99
FB6D
FB23
FB22
FB36
FAF5
FAA4
FAE8
FB98
FBA2
FAAF
FA46
FC55
00A0
048B
05E1
051B
044F
048D
051A
0505
0486
045C
049F
04C9
04A6
0495
04D0
0506
04F2
04C7
04CB
04DB
04C9
04C3
04F2
04FC
048B
041E
049C
05C4
05C3
031F
FEBF
FB4C
FA59
FAF8
FB5C
FB15
FAF5
FB5B
FBA7
FB6A
FB20
FB5B
FBBE
FB8E
FAE8
FAB1
FB37
FBB8
FB8A
FB12
FB01
FB39
FB24
FAD4
FAED
FB70
FB7F
FADE
FAEC
FD35
013C
0495
058E
04EA
0483
04E8
0530
04C1
0435
0451
04D6
04F8
0495
0446
046B
04B0
04B7
04A7
04C1
04E6
04E3
04DE
04FF
04FC
0495
044A
04D7
05CC
0563
0270
FE1F
FB0A
FA7D
FB4D
FBA8
FB33
FAD8
FB0D
FB4C
FB2B
FB08
FB54
FBBB
FBA4
FB29
FAF7
FB42
FB81
FB58
FB2C
FB5E
FB97
FB5F
FB02
FB1A
FB6F
FB28
FA59
FAA2
FD6D
01D6
053C
05FD
0503
0446
047F
04F3
04FD
04DE
04FD
0528
04FD
049D
047D
04AF
04D7
04CA
04BC
04CA
04C1
049A
04A8
04F9
0506
0485
042C
04D7
05E9
0564
0228
FDA6
FA9C
FA2F
FB07
FB56
FAEC
FACA
FB48
FBAA
FB60
FACC
FAA0
FAE1
FB1C
FB25
FB2F
FB48
FB43
FB2C
FB4F
FB98
FB8A
FB10
FADA
FB58
FBCE
FB3F
FA3F
FADC
FE3B
02C9
05A6
05B4
048C
043D
04FD
0589
052E
0488
0466
04C7
0528
054B
0546
0521
04D9
049E
04AB
04D2
04B1
045A
0454
04B9
04EF
04A5
0487
0541
0600
04DB
0123
FCA5
FA04
FA04
FB1E
FBA2
FB6D
FB41
FB4F
FB2A
FAC8
FAAB
FB04
FB57
FB34
FADE
FAD2
FB08
FB24
FB2A
FB75
FBE9
FBEC
FB62
FB0C
FB5C
FB9A
FAF3
FA30
FB4C
FEFC
035E
05CA
05A8
04B6
0497
0516
051E
0492
044E
04B2
0527
051D
04D5
04D6
0516
0524
04E6
04B0
04AF
04B4
04A7
04B8
04DF
04C0
045F
046C
0534
05A1
040F
0062
FC8D
FAAA
FAD2
FB68
FB41
FABE
FABC
FB35
FB83
FB76
FB65
FB6B
FB42
FAE4
FAC4
FB1A
FB71
FB49
FAD7
FAB9
FB03
FB3C
FB43
FB7F
FBEF
FBC1
FAA8
FA00
FBB4
FFCA
03E8
05B1
0531
045B
0485
052F
054E
04E0
049B
04B9
04D2
04B6
04B1
04E3
04FC
04C7
0496
04C4
0513
050F
04CF
04CF
050F
04F8
0470
0443
04E6
0542
03AB
0009
FC50
FA7B
FA95
FB25
FB29
FAEE
FB07
FB4D
FB50
FB2D
FB48
FB8D
FB86
FB26
FAE3
FB00
FB31
FB2A
FB20
FB5C
FB9E
FB6C
FAEF
FAD2
FB2C
FB3B
FAB8
FAC6
FCD3
009D
041F
05A3
0566
04DC
04DC
050B
04F1
04C3
04DC
0515
0510
04E0
04D5
04E6
04CD
0496
049D
04E2
04ED
048B
0443
0495
0520
051E
04B3
04D9
05AA
0598
0315
FECC
FB3F
FA25
FAC8
FB55
FB15
FAC9
FB20
FBB2
FBC4
FB59
FAF8
FADA
FAD8
FAF3
FB51
FBC3
FBC7
FB40
FAB1
FA99
FAD8
FB09
FB30
FB85
FBB4
FB22
FA2C
FA78
FD43
019E
050A
05F5
051C
0453
0477
04F7
050A
04B3
046A
046A
049E
04ED
0534
0534
04E3
04A4
04D2
0534
053A
04D8
04A4
04EE
0528
04BB
0426
0475
0581
057C
02E4
FE91
FB0D
F9FA
FAA1
FB44
FB2B
FAF3
FB3B
FBB5
FBC9
FB71
FB21
FB15
FB21
FB1C
FB13
FB15
FB1A
FB20
FB2C
FB2C
FB06
FAE3
FB16
FB98
FBC4
FB22
FA67
FB1E
FDFC
01D4
04A1
0577
0517
04BD
04D8
050E
050E
04EA
04CA
04AD
049B
04B9
04FD
051D
04F5
04C4
04C5
04C9
048E
0453
0496
0533
0554
0494
03D4
043F
0572
0567
02B0
FE58
FAFA
FA1C
FAE3
FB7D
FB2E
FA98
FA77
FABB
FAF8
FB1E
FB60
FBA8
FB9F
FB35
FACE
FAC3
FB03
FB49
FB7A
FBA4
FBB4
FB80
FB17
FAE1
FB23
FB93
FB96
FB08
FAA4
FB7F
FE08
017E
046B
05C2
05A3
0507
04C7
04F3
051D
0507
04D9
04C0
04A1
045E
0431
046E
04F4
0539
04FE
04B4
04DD
054D
0557
04CD
044B
0466
04D3
04E0
048E
0492
050A
04CB
0294
FECA
FB6C
FA12
FA70
FB0D
FB18
FAFA
FB43
FBB2
FBBA
FB6C
FB61
FBB8
FBDB
FB5F
FAB5
FA98
FB0A
FB57
FB1F
FAD9
FB14
FB8D
FB92
FB1B
FAF5
FB97
FC45
FBEC
FACE
FABA
FD27
015D
04ED
0612
054A
0472
049F
0547
055C
04BD
0428
0429
047F
04B2
04B9
04D6
04FD
04DD
0479
044C
04A3
0519
0514
04A3
0473
04D5
0539
04FD
0471
0476
0511
04E5
029F
FEBC
FB5B
FA1B
FA97
FB34
FB19
FAD6
FB28
FBC6
FBD6
FB3B
FACC
FB24
FBCA
FBDC
FB4E
FAE6
FB14
FB5A
FB1F
FAA9
FABC
FB67
FBCE
FB64
FAC9
FAEF
FBAE
FBE7
FB43
FB1D
FD1C
0105
04AA
061C
058D
04AC
0497
04F0
04ED
0491
0478
04C7
04FE
04CF
049E
04DF
0552
054D
04BB
044F
0491
051E
0532
04BE
0470
04AA
04E1
0478
03D7
0403
050A
055E
035E
FF59
FB89
F9E7
FA55
FB2F
FB45
FADF
FACA
FB1F
FB4E
FB19
FAEA
FB1E
FB6F
FB61
FB06
FAE9
FB3D
FB88
FB4E
FAD0
FABF
FB44
FBC5
FBBA
FB6B
FB78
FBD4
FBBD
FB06
FAE0
FCCC
00AE
0473
0603
0557
0445
044D
052A
05AE
056E
0511
0525
0559
051F
0497
045E
04A1
04EA
04E3
04CB
04E4
04E7
0472
03D5
03D4
048C
0518
04BF
0406
0419
0507
0548
035B
FFA1
FC25
FA8D
FAA9
FB20
FB0F
FAB8
FAB3
FB07
FB37
FB0B
FAD7
FAF5
FB43
FB59
FB23
FB03
FB4A
FBC1
FBEB
FBA1
FB41
FB2A
FB49
FB58
FB63
FBAD
FC0C
FBE6
FB1B
FAC0
FC4E
FFE7
03CE
05EA
05CA
04D0
0471
04CD
0518
04F0
04BD
04DD
0510
04EF
04A0
049C
04EB
0510
04C8
0477
0499
0504
0523
04CF
0488
04A8
04D0
0481
0401
0429
0510
056F
03CD
003A
FC83
FA81
FA6C
FB09
FB34
FAE3
FAB3
FAEB
FB3B
FB54
FB44
FB3F
FB43
FB33
FB1B
FB28
FB50
FB52
FB0F
FAD2
FAF9
FB6C
FBAC
FB7E
FB45
FB7B
FBEB
FBCF
FAEE
FA62
FBBE
FF4E
0366
05CE
05DB
04DB
0474
04F2
056D
053E
04C8
04B6
04FD
0505
04A4
045D
0494
04F8
050D
04E0
04DD
0509
04F6
0480
0432
047C
04F2
04D1
042F
0414
04F2
0598
043E
00A2
FC95
FA41
FA29
FB0E
FB89
FB51
FAF5
FAE0
FAF8
FB03
FB0A
FB2C
FB5E
FB79
FB78
FB7A
FB8B
FB87
FB4F
FB03
FAF0
FB2A
FB65
FB56
FB25
FB38
FB85
FB74
FAC2
FA58
FBBC
FF51
0376
05DD
05D6
04CB
0473
04F7
054A
04E4
0471
04AB
053F
0544
0495
0400
0420
0495
04AD
0469
0459
04A9
04E4
04BF
049A
04E4
054E
052B
0483
0442
04F3
05A0
0490
013D
FD29
FA81
FA11
FAD4
FB5E
FB4D
FB35
FB7D
FBCB
FBA7
FB37
FB07
FB45
FB89
FB78
FB40
FB43
FB81
FB97
FB61
FB2E
FB3E
FB57
FB23
FAD2
FAEE
FB7E
FBBC
FB1B
FA6B
FB59
FE99
02C5
0589
05E0
04DC
0437
0478
04D2
0490
040B
0404
047D
04C8
0496
0465
04B9
0541
0546
04B9
0458
049E
0516
0508
048A
045B
04B8
0500
04C3
0486
04F6
0582
0494
0175
FD7B
FADB
FA73
FB3B
FBBB
FB9A
FB6A
FB83
FB9C
FB79
FB52
FB70
FBA4
FB8C
FB22
FAD9
FB00
FB5B
FB71
FB32
FB05
FB34
FB82
FB81
FB31
FB10
FB65
FBC1
FB84
FAEF
FB64
FDFD
01FF
052D
05F0
04E6
03FB
0433
04DD
04E5
0458
0423
04A4
0531
051F
04AC
047B
04A2
04B0
0488
048B
04E5
052B
04F5
0490
0497
04F6
04F2
0446
03C5
0447
0535
04CC
020B
FE0D
FB13
FA59
FB1E
FBC3
FB8C
FAFD
FAD9
FB27
FB6A
FB61
FB3F
FB38
FB39
FB21
FB12
FB3D
FB82
FB87
FB33
FAE7
FAFF
FB4F
FB66
FB3C
FB49
FBB8
FBFC
FB7C
FABB
FB36
FDE1
01DE
0512
0617
056B
04A0
04A2
0505
04F9
046F
0412
0453
04DF
051E
04F8
04D5
04F6
051D
04FD
04B6
04A1
04C1
04C1
048A
0470
04A3
04CA
048A
0441
04A0
056D
0526
028B
FE59
FAEB
F9E2
FAA1
FB5D
FB39
FAD5
FB03
FB99
FBD9
FB8F
FB34
FB2B
FB47
FB37
FB0C
FB07
FB22
FB24
FB10
FB2B
FB83
FBC2
FBA3
FB57
FB4E
FB8E
FB95
FB0C
FA81
FB25
FDA4
014A
046D
05D3
05A7
050A
04D8
04F3
04D2
0466
0430
0472
04CF
04D1
0494
0489
04BD
04C9
0481
0450
04A0
0526
0534
04AE
0438
0450
049E
0495
046D
04D1
0595
054F
02CD
FEB7
FB41
FA0A
FA9A
FB31
FAD7
FA2A
FA3E
FB2A
FC08
FC25
FBBB
FB6B
FB66
FB62
FB36
FB22
FB60
FBB2
FBB1
FB5C
FB16
FB13
FB2B
FB3D
FB7A
FBEC
FC0E
FB56
FA44
FA65
FCCF
00C3
0432
05B6
05B2
0575
0598
05B0
054A
04AA
045B
0472
0492
047E
0465
0476
0489
0465
0435
045A
04D9
052B
04DA
0428
03D7
0446
04F2
051D
04C2
0499
04F0
04D5
02F8
FF61
FBDA
FA3D
FA95
FB4F
FB30
FA97
FA96
FB52
FBE4
FBAF
FB32
FB2B
FB86
FB9C
FB46
FB0B
FB44
FB96
FB8B
FB54
FB75
FBE9
FC13
FBAA
FB35
FB4B
FBA2
FB74
FAD4
FB06
FD31
00E1
043A
05B4
0571
04CC
04C1
051A
0520
04A7
042E
0423
0463
0497
04B7
04E9
0516
04F0
0480
0448
04A4
0528
051C
0481
0421
046F
04D7
0497
0401
042B
053F
05B2
03BE
FF8C
FB68
F98F
FA1E
FB5A
FBB8
FB2C
FAA5
FABF
FB42
FBA5
FBA9
FB75
FB42
FB27
FB2A
FB4D
FB7E
FB8C
FB65
FB3A
FB4F
FB98
FBB4
FB6C
FB16
FB36
FBB4
FBCB
FB21
FAB4
FC20
FFB2
03B6
05FC
05FD
0512
04B7
050F
054C
0507
04A8
0498
04AF
04A2
0492
04BD
04FB
04E8
0498
0497
0513
0577
0520
0453
0400
0488
052B
04FB
0425
03C8
0467
04F6
03C9
0078
FC89
FA1B
F9F7
FB0C
FBBD
FB68
FAAA
FA5C
FAB3
FB4C
FBBC
FBDC
FBB6
FB65
FB19
FB02
FB22
FB46
FB3C
FB08
FAD2
FAAF
FA9E
FAB6
FB18
FBA0
FBDC
FB83
FB03
FB4F
FD16
0011
0322
051F
05A5
0544
04E1
04EC
0522
0512
04B7
0478
049B
04E6
04F3
04B9
0488
0491
04B4
04D5
0507
0540
0535
04D1
0480
04AD
050D
04EA
043C
03F2
04AF
0577
046D
0108
FCFD
FA8E
FA50
FB01
FB43
FAE4
FA80
FA7D
FABC
FB00
FB28
FB23
FAFC
FAFA
FB66
FC09
FC3B
FBB3
FAF0
FAA3
FAE0
FB35
FB5B
FB67
FB61
FB29
FAD6
FADE
FB6B
FBDF
FB84
FAC9
FB36
FDC3
018C
0496
05B5
055F
04C1
0488
04A6
04DF
0515
0536
0529
04FC
04E2
04E7
04DF
04B6
04A6
04DD
0523
0519
04BB
046B
0469
048A
0495
04A6
04EA
052C
0503
0486
045D
04CF
04FE
039D
007A
FD04
FAFA
FAC4
FB59
FB8E
FB31
FAC5
FAA9
FACC
FAF9
FB17
FB14
FAE1
FAA2
FAA3
FAFE
FB64
FB81
FB6D
FB7F
FBB9
FBC4
FB86
FB4D
FB4B
FB3D
FAEF
FAC6
FB35
FBCC
FB8F
FA8B
FA76
FCF6
015F
0502
05F9
0503
0439
048C
0539
0561
052B
0529
0560
0569
053F
053D
0566
054C
04D8
0492
04CE
051B
04E3
0450
03FF
0423
046C
04AF
050F
0571
0554
04AB
044B
04D4
055C
0414
0092
FCB4
FAB1
FACB
FB7D
FB95
FB3D
FB0D
FAFE
FAB5
FA53
FA4E
FAA7
FADB
FAB9
FAA5
FAE0
FB11
FAF2
FAE7
FB5C
FBF3
FBEA
FB3D
FABA
FAD8
FB1B
FAFE
FAE3
FB6B
FC28
FBF4
FAD5
FAAD
FD23
015E
04AC
0567
0482
03FE
049A
057E
05CC
05A2
057D
0563
0521
04E4
050F
0586
05B8
0563
04E3
04A3
0499
0489
0487
04D3
0548
0573
0531
04DC
04B1
047F
0432
0441
04FA
0580
0441
00D3
FCD9
FA86
FA5E
FAFF
FB0B
FA99
FA77
FAC2
FAE3
FAA7
FA8C
FAE2
FB3F
FB25
FAC8
FAB8
FB09
FB45
FB3D
FB3D
FB62
FB54
FAF4
FAC1
FB16
FB74
FB35
FAAF
FACB
FB88
FBBE
FAF5
FAB2
FCEC
014E
051E
0644
0577
04D3
0521
057D
053D
04EB
0523
057B
0540
04AC
049B
0522
0566
04FA
048E
04CB
0540
0523
0496
0464
04BB
04FF
04DA
04B7
04E3
04EC
0476
041F
04B1
0574
0475
00F2
FCBD
FA5D
FA53
FB02
FB00
FA81
FA66
FACC
FB19
FB09
FAF3
FB0B
FB13
FAF0
FAF1
FB38
FB5C
FB13
FACC
FB0F
FB95
FBA1
FB27
FAF0
FB60
FBCE
FB87
FAF6
FB0E
FBB6
FBC1
FAE4
FABD
FD01
011D
0486
0586
04E8
048F
051C
05B2
059B
053F
053F
056B
053B
04CF
04C2
0527
0557
04EC
045B
044C
04AE
04EE
04DB
04C8
04DE
04D9
0496
0471
04A4
04CB
0482
0436
0491
051C
0438
010D
FD06
FA98
FAA1
FBA3
FBC6
FAE6
FA2B
FA3B
FAAC
FAEC
FB01
FB22
FB38
FB26
FB1E
FB59
FB8E
FB56
FAEC
FAFB
FB86
FBC2
FB46
FABD
FAE8
FB71
FB87
FB3F
FB73
FC2D
FC4B
FB4D
FAC4
FCC5
0106
04B4
05A8
04B7
0426
04B5
0548
050B
04A4
04EC
0589
058F
04F0
048B
04CA
0522
0514
04E6
04F6
0504
04B7
046C
04A8
052A
0536
04BC
046D
0490
0489
03F4
039A
045B
055C
047A
00F0
FCB8
FA7C
FAB5
FBA0
FBB0
FB11
FAB6
FAE3
FB26
FB3D
FB4C
FB50
FB0B
FA9C
FA8B
FAFA
FB51
FB18
FAC0
FAF4
FB89
FBB4
FB4E
FB12
FB7A
FBF4
FBC4
FB37
FB3B
FBCF
FBDC
FB00
FAB4
FCCB
00F9
04C2
0617
0560
048F
04BC
054C
0554
04EC
04C9
0510
0535
04E7
0487
0494
0502
0559
0550
0500
04AF
048E
04AD
04E4
04D9
0465
03EC
0404
049B
04EF
049F
0453
04CD
056C
0475
0129
FD14
FA9C
FA77
FB2C
FB2F
FA96
FA60
FACE
FB34
FB28
FB05
FB1D
FB32
FAFC
FAC9
FB0D
FB8B
FB98
FB27
FAEE
FB44
FBA1
FB87
FB53
FB8C
FBE5
FBB9
FB3E
FB4E
FBF1
FC03
FAFF
FA67
FC56
00A3
0499
05EF
0535
0496
0507
05AC
05A2
053A
051C
0533
04FF
0494
0484
04E7
052A
04F9
04B5
04B6
04BA
0475
043A
046C
04BC
049A
042D
042B
04A4
04C8
0433
03C8
0476
0565
047E
010D
FCF7
FAB4
FAA1
FB22
FAF9
FA85
FA9A
FB13
FB2A
FAB8
FA67
FAA8
FB23
FB55
FB41
FB32
FB31
FB24
FB34
FB90
FBF7
FBF8
FBA6
FB85
FBBE
FBCA
FB44
FAB5
FAE9
FBA7
FBD4
FB26
FB0D
FD2D
0127
04B3
05FD
0568
04A9
04B4
0512
051B
04F0
0509
0557
0568
0529
04FC
0514
052D
050D
04E1
04E4
04E3
0483
03E7
039C
03E5
0469
04BF
04DC
04CC
0474
03FF
041F
052D
0610
04E4
0124
FCCB
FA7E
FAC6
FBBC
FB8B
FA71
F9DC
FA52
FB0A
FB3E
FB0C
FAE2
FACB
FAAB
FAB8
FB25
FB95
FB82
FB18
FB0F
FB82
FBB1
FB3C
FAD5
FB31
FBD0
FBBA
FB08
FAD0
FB60
FBA7
FAFF
FAB9
FCC9
00EE
047D
0570
049B
0430
04DA
0579
0540
04D0
04F6
0565
0557
04DF
04C2
052A
0561
0503
04A2
04CE
0527
0507
0495
0476
04B3
04BC
0473
045F
04C0
0503
04BC
0489
0534
0611
053E
01EF
FDC1
FB16
FA94
FAF3
FAF2
FA91
FA67
FA8C
FAAC
FAB3
FAD6
FB13
FB20
FAFF
FB0E
FB62
FB85
FB31
FAD5
FAF3
FB4B
FB3F
FADA
FAD7
FB73
FBF1
FBA6
FB08
FB06
FB7A
FB49
FA3A
F9ED
FC1A
003C
03D5
051C
04BA
0483
052C
05E1
05DA
056C
054C
057D
0576
0514
04B8
049C
0492
047E
0495
04E4
0508
04B7
0459
048F
0534
056E
04E9
0453
045C
04B7
04B6
047D
04C8
0564
04D3
020E
FE2F
FB87
FB19
FBAC
FBA5
FAE4
FA60
FA80
FABB
FAA9
FA99
FAE7
FB59
FB78
FB44
FB1B
FB1D
FB23
FB37
FB90
FBFA
FBE8
FB52
FAF3
FB40
FBA5
FB6F
FB00
FB39
FBEA
FBC5
FA70
F9C0
FBE0
006F
0482
05D7
0519
0474
04CD
054E
0530
04C9
04B6
04DD
04D0
04A2
04B4
04EF
04DF
048C
048D
0500
0530
04A8
0408
0422
04B2
04C1
0427
03D0
044F
04F7
04E6
0472
04A3
054F
04C3
01DB
FDBB
FAC8
FA1E
FAC7
FB49
FB39
FB18
FB38
FB61
FB53
FB2A
FB1B
FB2B
FB46
FB6B
FB8A
FB76
FB36
FB20
FB64
FBB5
FBAA
FB61
FB55
FB99
FBB1
FB5D
FB1B
FB73
FBF4
FBA3
FA97
FA7A
FCD3
0105
04A8
05F3
055D
04A8
04CA
053E
052F
04A4
0442
045F
04BB
04F9
04FC
04CB
047E
0447
045C
04A4
04BA
046E
0419
042B
048E
04C5
04B4
04C1
051D
054C
04E7
0466
048E
050A
044B
0155
FD41
FA61
F9D3
FA93
FB0D
FAED
FAE7
FB4D
FB9F
FB76
FB27
FB2B
FB62
FB53
FB00
FAEA
FB46
FBAE
FBC5
FBAF
FBB2
FBB2
FB75
FB29
FB25
FB5A
FB69
FB40
FB32
FB4C
FB20
FA97
FAB1
FCB2
006D
040B
05D9
05E4
0576
0563
0577
0551
0510
04FF
050B
04F3
04C5
04BF
04D7
04BC
046B
0442
046C
0499
048F
0496
04EB
0531
04EA
045C
044A
04D6
052C
04B8
0429
0481
0551
04BE
01B6
FD8A
FAAC
FA22
FACD
FB27
FAE7
FABC
FAFC
FB3F
FB25
FAF4
FB1D
FB86
FBA9
FB47
FABC
FA8A
FAD1
FB45
FB83
FB64
FB15
FAE6
FAFD
FB37
FB5A
FB4F
FB33
FB23
FB25
FB32
FB48
FB54
FB34
FB12
FBA6
FDB6
0113
0452
05EE
05AE
04C1
045B
0492
04B8
0480
0458
04A0
0510
052D
0504
0503
0537
052A
04AC
044A
049C
055C
05AD
0546
04D6
0500
0565
053C
048F
0443
04C6
0551
04FC
042E
0426
0518
056D
0383
FFBA
FC38
FAAB
FACF
FB43
FB3F
FB0C
FB17
FB40
FB34
FB05
FB09
FB44
FB5F
FB30
FAFA
FB0A
FB4D
FB68
FB28
FAC4
FAA2
FAD9
FB20
FB29
FB09
FB1B
FB78
FBBA
FB7E
FB05
FB09
FBB8
FC32
FB9A
FA8F
FAFD
FDFF
0254
0577
0622
054C
04AA
04C8
0504
04E7
04CC
0514
056E
0553
04DB
049A
04C3
04F9
04ED
04D3
04F5
052B
050C
0493
0430
043F
048F
04B6
049F
048C
049F
04A5
046E
0424
043D
04EE
059C
050A
0264
FE59
FADF
F992
FA46
FB59
FB84
FAFD
FABD
FB0B
FB45
FAFE
FAAA
FAD9
FB4B
FB53
FAE2
FA99
FAD8
FB3C
FB4B
FB35
FB75
FBEB
FBF4
FB6D
FB16
FB8A
FC49
FC59
FBA8
FB2A
FB7F
FC02
FBA3
FA8D
FA5E
FC7A
0069
0420
05E6
05C1
0502
04C5
0511
054F
053B
0522
0543
0560
051C
04A2
0483
04E8
0544
050F
0483
044F
049E
04E2
04AB
0450
0464
04C2
04B0
0408
0391
03F2
04AB
04BD
0424
03FD
04E5
05B8
0497
0114
FCEB
FA56
F9F6
FA9E
FAF2
FAAC
FA61
FA7C
FACF
FB03
FB07
FB02
FB11
FB2F
FB54
FB75
FB6F
FB2F
FAE5
FAEF
FB6B
FBED
FBE9
FB5D
FAE6
FB08
FB93
FBE3
FBBC
FB92
FBD5
FC36
FBEF
FAE0
FA22
FB31
FE67
026F
055A
0635
05A3
04FD
0500
0564
0590
056A
0548
054B
052C
04BF
045B
047A
050A
056B
0539
04C2
0486
0489
0472
0447
047A
051D
058B
0533
047B
0447
04BE
0512
04AC
0418
0441
04E7
048B
021E
FE62
FB46
FA08
FA52
FAF6
FB2A
FAF3
FABC
FAC0
FAE4
FAEE
FAD0
FAB6
FACC
FB02
FB21
FB0C
FAF3
FB0C
FB47
FB65
FB5F
FB63
FB72
FB4E
FAF4
FAC7
FB04
FB55
FB48
FB16
FB5B
FC13
FC58
FBAB
FB1E
FC75
FFFB
03D6
05E5
05E0
052E
0505
0557
058B
0584
0588
059B
0577
0521
0505
0550
0592
0555
04C5
0474
048C
04B2
04A1
0491
04D3
0543
0564
04F6
0455
0415
044F
0480
0432
03AA
03B3
0490
0546
0444
010A
FD05
FA69
FA16
FAE7
FB32
FA93
F9EC
F9F6
FA5E
FA75
FA39
FA3B
FAAD
FB18
FB13
FADD
FAF7
FB55
FB71
FB10
FAA5
FAB9
FB40
FBB7
FBCE
FBB3
FBB5
FBD6
FBE1
FBDB
FBFF
FC49
FC3F
FB95
FAE0
FB69
FDE9
0197
04AA
05E4
0599
050C
0510
0576
05AD
058D
0555
0530
0515
050B
0533
0580
05A0
055A
04F1
04DB
0529
0564
0528
04A2
0451
0458
045E
0417
03B9
03B0
040B
0459
043E
0407
0455
0517
0522
0335
FF7F
FBD3
FA11
FA61
FB48
FB64
FAC7
FA6B
FABB
FB28
FB1D
FAD2
FAC3
FAE6
FACC
FA6B
FA47
FAAB
FB37
FB5A
FB1C
FB00
FB43
FB99
FBAF
FBA6
FBBF
FBDB
FBAC
FB4A
FB33
FB9E
FC0C
FBCD
FAF5
FA9F
FC0B
FF56
0320
0591
05E9
0505
045C
0495
0522
0539
04E1
04B9
04FF
0543
052B
0502
052E
057A
055B
04D3
0489
04E0
0558
0539
0494
0431
047C
0503
052D
0506
04F8
0501
04BC
042D
03F6
0478
04FF
043C
019E
FE15
FB55
FA5C
FABF
FB59
FB6A
FB0F
FAD1
FAEE
FB2C
FB3E
FB2F
FB32
FB3A
FB0B
FAB1
FA97
FAF7
FB74
FB8B
FB3F
FB05
FB16
FB21
FAE0
FA9D
FAC7
FB30
FB3C
FADD
FAD7
FB9A
FC63
FC16
FAF2
FABF
FCF3
00EA
046C
05D9
057D
04CC
04B0
04F1
0504
04D5
04BD
04E7
051F
051E
04E5
04B4
04B7
04DA
04E9
04D9
04CF
04E2
04F8
04F2
04D7
04D0
04E8
0507
0515
051B
0517
04E1
046D
0419
0464
0522
0539
0389
002E
FCA9
FA9C
FA63
FB09
FB66
FB2F
FAE3
FAE7
FB15
FB0C
FACB
FAA6
FAD0
FB14
FB21
FAFB
FAF3
FB35
FB8A
FBA7
FB96
FB8F
FB95
FB74
FB31
FB1E
FB56
FB6E
FAF9
FA48
FA24
FABF
FB4E
FB1A
FAC0
FBC9
FED6
02A6
0546
05F6
0592
0547
055B
055A
04FB
0483
045C
0493
04DD
04FE
04FB
04F6
0502
0511
0507
04DA
04AC
04A2
04B2
04B6
04B0
04C5
04F3
0505
04F1
04FB
0542
0569
050D
0485
04A6
0566
0547
02C1
FE58
FA88
F94A
FA25
FB22
FB32
FAED
FB26
FBA7
FBB1
FB38
FAEB
FB1E
FB53
FB10
FA9F
FA8F
FAD9
FAFD
FAD8
FACD
FB15
FB55
FB25
FAB7
FAA3
FB1A
FB99
FB94
FB2D
FB03
FB4C
FB83
FB17
FA62
FAA2
FCD9
0098
0410
05A1
0551
048F
0490
0528
056C
050A
049D
04BA
052A
0556
052B
0516
053F
0543
04E9
049D
04E5
0586
05BF
0555
04E3
04FC
0554
0532
048F
0433
0497
0524
04F2
0425
03DE
04A3
0554
042F
00DC
FD01
FAA8
FA58
FAF3
FB3C
FB0C
FAF2
FB2A
FB56
FB2D
FAE5
FAD7
FAFD
FB0F
FAFE
FAFF
FB23
FB2E
FAF0
FA9B
FA87
FABE
FAF2
FAEC
FAD4
FAED
FB32
FB65
FB6D
FB7C
FBC4
FC1C
FC13
FB7F
FAF8
FBAB
FE40
01EE
04E0
05CC
0526
047F
04C5
056D
0577
04D4
045F
0493
04EF
04E1
04A2
04BF
051F
0527
04BF
0493
0513
05A8
0579
04AF
0454
04DC
0578
053E
0475
041F
0476
04A1
040D
0364
03B6
04CC
04FA
02DB
FEF1
FB56
F9C7
FA37
FB41
FBAE
FB67
FB1C
FB37
FB6F
FB55
FAFA
FADB
FB1C
FB58
FB3A
FB02
FB22
FB83
FB9D
FB35
FABA
FAA8
FAE1
FAF4
FAE6
FB29
FBBD
FBF6
FB7A
FAF3
FB3B
FC07
FC28
FB47
FAD0
FC7D
0038
03F7
05CF
05C0
052E
0510
052B
04EB
0465
0424
0466
04E0
0532
054B
0547
051D
04B4
0434
0404
0457
04E1
051F
04E9
0496
0490
04D4
0501
04DF
04A7
04A5
04C5
04AD
0461
0461
04F2
055E
0457
0152
FD58
FA4C
F952
F9FA
FAEE
FB45
FB13
FAE1
FAEE
FB13
FB2C
FB4A
FB7F
FB9D
FB6E
FB0C
FAE7
FB3E
FBC1
FBE1
FB80
FB0E
FAF9
FB31
FB61
FB67
FB66
FB65
FB3E
FAFD
FB01
FB73
FBD3
FB80
FACB
FB18
FD75
014B
04B8
064E
062E
057A
0510
04FD
0500
0510
0540
056B
0550
04F2
04A3
0498
04AA
0498
046D
0478
04DC
0543
0539
04C0
0465
0492
04FE
0503
0481
0412
0431
048D
0486
0438
046E
054D
0586
038B
FF92
FBCC
FA40
FACF
FBB8
FBAE
FAF2
FA75
FA8F
FAE4
FB18
FB1F
FAF7
FA9D
FA53
FA8C
FB45
FBCC
FB8B
FAD6
FA84
FAD8
FB42
FB42
FB19
FB51
FBD7
FC0C
FBB1
FB52
FB7E
FBF7
FC0D
FB9D
FB44
FB68
FB95
FB1E
FA54
FA9B
FD05
00FA
047E
05F7
0588
04A4
0474
04E5
0538
0519
04EC
051C
0580
059A
053F
04CB
04A7
04DE
0530
055D
0548
04F7
0498
0473
04A0
04DE
04D7
0494
046A
0485
04A6
0496
0489
04CE
052B
0507
0463
0422
04E3
05C9
0504
01D5
FDA8
FACB
FA3C
FAFB
FB7B
FB40
FADE
FADB
FB0C
FB0E
FADB
FAB6
FABF
FADC
FAF9
FB1A
FB38
FB39
FB20
FB1C
FB46
FB66
FB42
FB00
FB0B
FB76
FBC9
FB93
FB11
FADE
FB21
FB5B
FB31
FB06
FB65
FBFC
FBD3
FABF
FA2B
FBC6
FF7B
0340
0522
0526
04C3
04F6
055E
0545
04CA
04A5
050A
0571
0566
0520
04FE
04F4
04BC
0472
0478
04D4
0510
04E7
04A8
04B9
04F4
04D8
045D
041E
0480
050F
050D
0482
0435
0493
050C
04E6
045F
0470
054C
0593
039C
FF89
FB94
F9F2
FAA9
FBCA
FBBC
FACC
FA51
FAD4
FB8B
FB9B
FB31
FB08
FB49
FB6E
FB38
FB13
FB5D
FBBF
FBB0
FB4B
FB23
FB5D
FB79
FB27
FAD6
FB14
FBA6
FBD5
FB82
FB53
FBAA
FBFA
FBA7
FB0A
FAF6
FB60
FB61
FAC1
FAE1
FD42
0167
04E6
05EA
050A
044B
04AE
056C
056B
04BE
0446
0464
04A2
048D
0457
046A
04BA
04D9
04A9
048A
04C6
0527
0542
0508
04C0
0497
0475
0449
0435
0456
0489
049A
0498
04B6
04DE
04C2
0475
049E
058E
0649
051E
0186
FD22
FA5D
FA19
FB11
FB93
FB49
FB0F
FB6A
FBD5
FBB3
FB39
FB10
FB4E
FB66
FB0B
FAA4
FAB4
FB1B
FB52
FB30
FB13
FB43
FB84
FB7C
FB41
FB30
FB5F
FB84
FB78
FB6B
FB7E
FB77
FB19
FAA8
FAA8
FB13
FB38
FAC5
FAA2
FC3F
FFCC
039F
05B1
059A
04BA
0478
04E1
051B
04CF
0482
04AA
04F9
04ED
04A6
04B3
0522
055C
0507
0498
04AC
051E
053C
04D5
0482
04C1
0537
0533
04B5
0467
04A1
04F3
04E7
04B0
04BB
04E8
04C1
0467
048D
053C
0524
02E6
FEEE
FB6E
FA2E
FAD2
FB9D
FB88
FB0D
FB01
FB5C
FB7F
FB38
FAFC
FB1F
FB5A
FB45
FAF8
FADD
FB11
FB44
FB3C
FB1C
FB18
FB18
FAF4
FACD
FAEF
FB4F
FB87
FB5C
FB23
FB4A
FBB1
FBCA
FB69
FB10
FB2C
FB62
FB0E
FA81
FB25
FDF6
020C
0529
05E7
0500
0446
0492
0537
0542
04C5
0486
04DA
054A
054E
0503
04D6
04E1
04DD
04AD
048F
04BC
050D
0534
051E
04F5
04CF
04A2
0478
0477
04A1
04BC
049F
0471
0471
0487
0471
044C
04A0
057F
05DC
0452
00C0
FCD5
FA9D
FA91
FB5E
FB8B
FB04
FAB9
FB27
FBB0
FB8B
FAD3
FA59
FA90
FB1B
FB61
FB4D
FB30
FB2E
FB1A
FAE4
FABF
FADD
FB1F
FB42
FB42
FB4C
FB6C
FB86
FB97
FBC0
FBED
FBC6
FB37
FAC6
FAFF
FB9B
FBAF
FB01
FACB
FC8D
002D
03C0
056C
0536
0499
04A5
0516
0533
04FC
04F7
0540
055B
0500
04A1
04C4
053C
055F
04F3
047A
047D
04DA
0514
0500
04E4
04E6
04CA
0461
03F2
03E6
043F
04A0
04DE
0521
0565
0540
048B
03FE
047C
05A1
0594
02DD
FE55
FAAE
F9D2
FB12
FC2C
FBCE
FAA5
FA0B
FA5C
FAEC
FB27
FB24
FB2E
FB37
FB18
FAF2
FAFF
FB27
FB22
FAFB
FB19
FB92
FBE2
FB8E
FAE1
FAA0
FB0B
FB8E
FB92
FB41
FB28
FB5D
FB72
FB3F
FB30
FB86
FBBA
FB36
FA8E
FB59
FE70
029E
0592
0624
053E
0496
04D0
054A
054D
04F6
04C8
04E3
04F5
04D4
04B0
04B8
04D2
04D9
04DE
04FD
051B
0506
04D4
04D6
0517
053A
04F5
0487
0464
048F
04A2
047A
047D
04EA
0545
04ED
0429
0413
050E
05C9
045D
0084
FC3B
F9E2
F9FA
FB0E
FB8D
FB43
FAF5
FB14
FB52
FB4C
FB1C
FB10
FB26
FB22
FAF8
FADF
FAEC
FAF2
FAD1
FAB4
FAD2
FB16
FB3E
FB3C
FB44
FB63
FB63
FB27
FAF8
FB28
FB84
FB8A
FB34
FB24
FBBA
FC47
FBC6
FA76
FA2D
FC8A
00F2
04DD
0646
0584
047D
0474
0504
0533
04D7
049A
04E1
054D
0555
04FF
04B9
04BB
04DC
04F2
0509
052E
053D
051A
04E7
04E2
0500
0500
04CA
049B
04A3
04C2
04BD
04A2
04A9
04B9
046E
03D1
039C
0467
0584
053D
0292
FE87
FB59
FA5C
FAEB
FB76
FB45
FADA
FAE2
FB43
FB73
FB46
FB12
FB15
FB23
FAFF
FAC6
FABC
FAE9
FB11
FB18
FB1E
FB3B
FB4B
FB33
FB1A
FB38
FB7B
FB94
FB71
FB5F
FB98
FBDF
FBD6
FB90
FB70
FB80
FB3D
FA73
FA09
FB5F
FEBD
02AA
0531
05AF
051E
04BD
04D2
04E7
04C6
04BB
04F6
052B
0507
04BC
04B9
0501
0522
04E0
0498
04BB
0526
054F
04FB
0487
045B
0466
045D
043C
043F
046D
048C
048A
04A9
04FE
051A
0498
03F2
042B
0557
05F3
0440
0055
FC58
FA69
FA9E
FB58
FB4C
FAB9
FA8B
FAF5
FB54
FB39
FAEE
FAE9
FB1D
FB30
FB11
FB06
FB26
FB31
FB07
FAF0
FB32
FB96
FBAA
FB68
FB40
FB72
FBA8
FB84
FB37
FB3E
FB94
FBA8
FB3F
FAF1
FB4D
FBDE
FBA3
FAA5
FA7E
FCB4
00C5
0463
05C3
054B
04B5
04FD
059B
05AE
053A
04E8
04FE
051F
04FA
04C3
04CA
04F4
04EE
04BC
04A9
04C3
04BF
047E
045B
04AF
0531
0543
04CA
045D
047D
04E4
04F6
04A8
047F
04B2
04D2
048C
0457
04D1
057B
04C6
01CE
FDB4
FAB6
F9FB
FAA4
FB22
FAF1
FAB4
FAEB
FB46
FB48
FB15
FB22
FB68
FB6B
FB07
FAC3
FB16
FBAD
FBCD
FB4C
FAC6
FACA
FB22
FB42
FB0F
FAF0
FB1F
FB5C
FB5E
FB44
FB4D
FB61
FB3C
FB07
FB37
FBC6
FBF4
FB4C
FAB4
FBD1
FF21
031C
0592
05D7
0529
0501
0587
05DA
057B
04DC
0493
049E
04A0
048E
04AB
04F6
0511
04CA
0473
046F
04A4
04B5
049C
04B7
0521
056C
0534
04C2
04BA
0531
0589
0549
04BF
0482
0492
047B
043B
046B
052D
055E
0389
FFB2
FBBD
F9AD
F9BF
FA8A
FAD2
FAA5
FAB5
FB2B
FB86
FB73
FB3B
FB3A
FB57
FB44
FB0F
FB09
FB41
FB6A
FB56
FB39
FB4D
FB66
FB30
FAC1
FA8E
FACD
FB28
FB46
FB46
FB76
FBB8
FB99
FB1C
FADF
FB40
FBA9
FB4C
FA8E
FB0B
FDD4
01EE
0512
05F0
054D
04C7
0500
055B
053B
04E5
04ED
054F
0575
051A
0499
0464
0479
048E
048F
04A4
04CF
04D5
049C
0460
0464
0499
04B9
04AE
04A0
04AE
04C9
04DD
04F3
0506
04F0
04A4
0469
048D
04E2
04DA
045B
0416
049C
0542
0471
0164
FD53
FA72
F9D6
FA9C
FB30
FB01
FAAB
FAC7
FB22
FB35
FAF0
FAC5
FAFA
FB5D
FB91
FB80
FB4E
FB21
FB12
FB32
FB6D
FB84
FB48
FAE7
FACA
FB12
FB6C
FB7C
FB54
FB44
FB59
FB51
FB19
FB00
FB38
FB72
FB4A
FAFE
FB34
FBEF
FC47
FB97
FACA
FBC0
FF25
0354
05D4
05CD
04A2
0421
04A7
053E
052B
04B4
047E
04A2
04C8
04C6
04C8
04E7
04FB
04ED
04E4
04FE
050D
04DC
048F
0487
04CD
04FD
04CB
046F
0454
0485
04AF
04A4
048B
0488
047C
0456
0455
04B5
0524
050B
047A
0445
04D7
052F
03B5
002D
FC5A
FA53
FA6D
FB30
FB3D
FAB3
FA85
FAFE
FB7B
FB6B
FB0A
FAE3
FB08
FB27
FB1F
FB21
FB3D
FB38
FAF8
FAD1
FB16
FB8C
FBA9
FB4F
FAFC
FB1B
FB7C
FB9F
FB6C
FB46
FB6D
FBAD
FBB3
FB7A
FB29
FAD2
FA90
FAB2
FB62
FC18
FBF5
FB07
FACE
FCDE
00E9
04A4
0601
0538
0435
044D
0502
0529
049A
0439
0499
053D
0564
050F
04CE
04D8
04D7
0495
0465
04A9
052E
0560
050F
04A9
04A3
04E6
0505
04D4
048C
047B
04B1
04FF
0529
0502
049F
0458
047F
04EB
0505
048B
0415
0474
0562
054D
02EA
FEE4
FB78
FA46
FAD2
FB64
FB18
FA8B
FAA5
FB4B
FBA3
FB4F
FACF
FABB
FB05
FB3A
FB2F
FB21
FB3A
FB4F
FB32
FAFF
FAE9
FAF3
FAFD
FB06
FB25
FB4E
FB4F
FB21
FAFF
FB19
FB4C
FB59
FB43
FB3D
FB4A
FB36
FB0B
FB25
FBA0
FBE4
FB57
FA7D
FAE8
FD95
018E
04A5
0598
0524
04D6
0538
0598
055B
04DC
04CB
0525
0542
04D0
0443
042D
0481
04CA
04DA
04EB
0527
0558
0542
0504
04E9
04F8
04F0
04B4
0485
04AB
0514
0567
055B
04ED
0455
03EB
0401
0491
051F
0524
04BA
049D
052E
0593
0451
00FD
FD0C
FA96
FA54
FB29
FB93
FB37
FAC8
FACC
FAFF
FAE9
FAA4
FA9C
FAE5
FB22
FB12
FAED
FB01
FB3C
FB4C
FB1D
FAF2
FB04
FB3A
FB53
FB41
FB22
FB0F
FB07
FB06
FB0D
FB12
FB0E
FB18
FB4B
FB85
FB71
FB05
FAC0
FB1D
FBCD
FBE2
FB14
FA87
FBDD
FF53
0338
0584
05BC
051C
04F7
0565
05AB
0567
04F9
04D2
04E6
04E9
04D3
04D4
04F4
04FB
04CC
049C
04AA
04E9
0516
050B
04DA
04A7
0485
0484
04A9
04D6
04E0
04C5
04C5
0502
053D
051A
04B3
0488
04CB
04FE
04A7
0425
0451
052B
0550
034A
FF62
FBA5
F9F6
FA56
FB4A
FB97
FB41
FAEA
FAD1
FAC1
FAA1
FAA1
FADB
FB16
FB1B
FB04
FB02
FB0D
FAFA
FADB
FAF2
FB40
FB70
FB48
FB08
FB12
FB60
FB8B
FB66
FB3C
FB4B
FB5D
FB1B
FAA8
FA7E
FAC0
FB09
FB12
FB2B
FBA4
FC08
FB89
FA67
FA4A
FCAE
0100
04DB
0653
05AD
04AD
048A
0509
055C
054E
053B
054A
0540
04FA
04B8
04BA
04E5
04F4
04E6
04E8
04FA
04E6
04A2
0476
0497
04D8
04EB
04DC
04EF
0523
0520
04BE
045A
0465
04C3
04F2
04C3
0499
04C3
04FC
04E2
04AC
04E6
0562
04EA
027A
FEA3
FB47
F9D3
FA0C
FAAD
FADF
FAC2
FABD
FAD0
FAC5
FAA8
FAC0
FB19
FB6E
FB84
FB6B
FB48
FB16
FACE
FA9F
FAC6
FB30
FB84
FB94
FB87
FB8C
FB85
FB45
FAF0
FAEA
FB43
FB8E
FB69
FAFE
FAC6
FAF0
FB3A
FB6C
FB8E
FB98
FB3E
FA7A
FA25
FB78
FEB4
0283
0512
05BB
0557
050E
052D
054B
0531
051D
0540
055E
0526
04BB
0486
04AE
04F2
050D
0500
04EA
04CD
04A3
0487
0497
04BB
04BC
049C
049D
04DB
0510
04F5
04B2
04AB
04E7
0504
04CE
049B
04C0
04F7
04B8
042B
042D
0507
0589
0406
0056
FC51
FA19
FA10
FADF
FB35
FAFC
FAD7
FAF9
FB01
FAC1
FA91
FAC8
FB39
FB79
FB6B
FB4B
FB37
FB10
FAD0
FAAE
FAD4
FB16
FB3A
FB4A
FB71
FB95
FB6A
FAFB
FAC1
FB03
FB5E
FB43
FACA
FAA3
FB14
FB86
FB65
FB0A
FB3E
FBF0
FC18
FB46
FAC4
FC72
0071
0496
0681
05F3
04A7
042F
0489
04D4
04BA
04A8
04ED
053C
0536
04F1
04C8
04D1
04E0
04E6
04FD
051B
0507
04C2
04A4
04E6
053D
0532
04D0
049E
04D5
0503
04B9
0437
041A
0477
04C0
049D
0473
04B6
051C
04F8
045F
0435
04CD
04F0
0305
FF1F
FB53
F9B0
FA3F
FB54
FB9A
FB33
FAF3
FB14
FB28
FAF6
FACF
FAF9
FB3C
FB3F
FB0E
FAF9
FB18
FB35
FB32
FB33
FB4C
FB4B
FB0F
FAE1
FB1B
FB9F
FBE4
FBA9
FB4A
FB3C
FB6B
FB6C
FB2A
FAFF
FB1F
FB4A
FB46
FB4B
FB9B
FBD2
FB4B
FA56
FA81
FD1B
0173
0524
065D
0588
047C
046A
04FE
0559
0547
0537
0560
057B
054A
04FA
04D1
04C4
049A
0456
0435
0451
0485
04A9
04C4
04D7
04BD
0462
040E
0423
0499
04F9
04F2
04B7
04A9
04CB
04DD
04D4
04EA
051B
0507
048D
043E
04AF
0552
0495
0194
FD6F
FA7A
FA00
FB20
FC01
FBC6
FB03
FA9A
FAAD
FAD0
FAD4
FAF0
FB41
FB8A
FB89
FB4C
FB12
FB01
FB13
FB40
FB7E
FBA9
FB9C
FB6D
FB5F
FB85
FB9C
FB70
FB34
FB38
FB6B
FB67
FB08
FAB7
FAD9
FB37
FB48
FAFF
FAE3
FB35
FB71
FB19
FAD0
FC04
FF3F
032D
05B6
0601
0510
0465
047A
04C0
04B3
047C
0479
04AD
04D4
04D6
04DC
04FB
0516
0512
04FA
04DC
04AE
0472
0452
046B
0490
0481
044E
044F
04A4
04EE
04D0
0477
0464
04AC
04DC
04A9
0474
04B6
0536
0540
04BC
0478
04FB
0560
0402
0076
FC61
FA02
FA06
FB31
FBEB
FBC0
FB3B
FAE3
FAC5
FACE
FB15
FB8D
FBE0
FBC6
FB6B
FB38
FB4E
FB70
FB72
FB6B
FB79
FB83
FB69
FB4C
FB5A
FB74
FB53
FB07
FB07
FB83
FBFD
FBDA
FB43
FAF4
FB3F
FB94
FB58
FAD3
FAC9
FB45
FB78
FB04
FAF6
FCC0
0057
03E3
058D
0548
0485
046F
04E0
051E
04F8
04CD
04D6
04DD
04AC
0468
0445
043A
042A
042A
046B
04CD
04F0
04B3
046C
0476
04B6
04D6
04C7
04C0
04CC
04A6
043F
0404
045D
04FE
052A
04B0
0435
044E
04AF
04AF
045F
0477
0506
04CA
0285
FEC1
FB9B
FA9E
FB36
FBAE
FB39
FA95
FAB2
FB71
FBFF
FBF2
FB9B
FB58
FB25
FAEF
FAE6
FB2C
FB75
FB63
FB16
FB0D
FB6E
FBC6
FBAC
FB55
FB46
FB90
FBC8
FBAD
FB7D
FB79
FB80
FB5C
FB48
FBA2
FC39
FC5C
FBC8
FB1B
FB02
FB45
FB2A
FAD6
FB95
FE52
021F
04E4
0584
04DC
047B
04D5
052C
04EB
0479
0481
04F3
0531
04FF
04BB
04BE
04DF
04D4
04B5
04CD
0503
04EB
0464
03E0
03D4
0422
0452
043F
0428
0432
042C
03FA
03EC
0451
04E8
051B
04C4
046A
0477
04AC
0491
043E
0438
0491
04B9
0467
042B
0497
04FE
03D1
008C
FCB0
FA61
FA34
FAE0
FAFE
FA8C
FA67
FAE4
FB74
FB9C
FB89
FB96
FB9E
FB55
FAED
FAEA
FB64
FBCD
FBBA
FB71
FB72
FBB7
FBC5
FB77
FB3C
FB6D
FBC5
FBC4
FB69
FB2A
FB3C
FB5D
FB4F
FB47
FB85
FBD4
FBCE
FB86
FB82
FBE9
FC2D
FBCF
FB2F
FB13
FB81
FBA1
FB16
FAF5
FCBB
0067
0417
05E1
05A9
04D9
0494
04C6
04D7
04B4
04B9
04E7
04DC
0482
0456
04B2
052F
0522
0486
0403
0414
047A
04B5
04B5
04C0
04DD
04BD
0452
0409
043E
04B2
04E0
04B3
048D
04A3
04B6
048E
045E
046B
0481
043C
03C5
03C7
046F
0500
04C6
042C
0438
04E3
04A8
0233
FE38
FAF9
F9F7
FA9A
FB48
FB4A
FB20
FB52
FBA3
FB9F
FB5D
FB4B
FB73
FB6D
FB19
FAE2
FB20
FB8D
FB9D
FB45
FAFE
FB0F
FB2F
FB05
FAB3
FAAA
FB09
FB7E
FBBE
FBD2
FBCF
FB9F
FB34
FAD8
FAE8
FB50
FB97
FB8E
FB90
FBEA
FC44
FC0A
FB57
FAFC
FB5A
FBBC
FB56
FAB7
FB8B
FEAA
02C3
057F
05DA
04E7
0447
0469
04A1
0476
043B
0456
0496
0495
046D
0493
0517
0579
0564
0528
053D
058B
058C
0510
0481
0456
0488
04C5
04E8
0504
050C
04D4
0473
044D
048D
04D6
04BF
0465
0440
0467
0479
0441
0426
0488
0507
04ED
044D
041D
04D5
0553
03D6
0021
FC18
F9F1
FA11
FB0C
FB7D
FB53
FB42
FB7D
FB8C
FB33
FAD7
FAE6
FB31
FB3C
FAF5
FAC5
FAEF
FB32
FB30
FAF4
FAD3
FAEF
FB16
FB23
FB2B
FB44
FB4C
FB24
FAF6
FB0A
FB5B
FB8F
FB6F
FB2E
FB17
FB29
FB3F
FB65
FBBD
FC13
FBF0
FB4E
FAE4
FB4C
FC0F
FC0D
FB1A
FAB5
FC87
005B
040D
05B2
056B
04D4
04FB
0579
0578
04FB
04A9
04CA
04F5
04D0
049A
04BD
0527
0564
0549
0520
052A
053E
0515
04C3
049D
04C0
04F7
050E
0511
0513
04FC
04B3
0460
0445
0466
0486
048A
0497
04BB
04B6
0454
03E8
03FD
048B
04E8
04B2
047B
0506
05DA
0549
0244
FDE0
FA90
F9B7
FA81
FB20
FADF
FA77
FAAA
FB31
FB4B
FADA
FA7A
FA99
FAEE
FB01
FACD
FAA9
FAB3
FAB5
FA94
FA88
FABF
FB0B
FB20
FB04
FB03
FB45
FB95
FBB1
FB97
FB6C
FB3D
FB0E
FAF9
FB18
FB45
FB40
FB15
FB21
FB84
FBC9
FB74
FACB
FAA0
FB2E
FBA9
FB50
FACA
FBCD
FF17
033B
05E2
0624
0536
04CA
053C
05B1
0588
0515
04F0
050B
04F4
04A4
0494
04FE
0577
0578
050F
04BB
04C3
04EB
04E6
04C0
04B7
04DB
050D
0534
054B
0542
0504
04AD
048B
04B8
04F4
04F2
04CC
04D1
04FE
04F3
048E
0439
045A
04A7
0487
0409
03F8
04A5
04F7
035D
FFC1
FC07
FA3A
FA84
FB56
FB5D
FACE
FAA2
FB19
FB8A
FB6E
FB13
FB04
FB3C
FB41
FAE8
FA8D
FA8C
FAC5
FAE7
FADD
FAD9
FAF0
FB03
FB00
FB06
FB28
FB42
FB30
FB10
FB19
FB3D
FB39
FAF7
FABF
FACD
FB02
FB21
FB3F
FBA1
FC28
FC4B
FBC8
FB26
FB14
FB71
FB7D
FB19
FB64
FD8D
0126
043E
055A
04EE
048F
0504
05A6
059A
050A
04C6
0513
0562
053C
04E3
04D8
0518
0531
04FA
04BD
04BA
04CD
04C2
04B0
04CE
0506
050D
04E3
04E0
052B
056E
0546
04D4
0491
04AB
04DC
04E9
04ED
0507
04FD
0490
0404
03EB
0453
04A3
047A
0453
04C9
0556
047B
017D
FD94
FAEB
FA6B
FB06
FB33
FAA6
FA3D
FA91
FB30
FB61
FB17
FAD3
FAD3
FADA
FAB9
FAA6
FADB
FB23
FB18
FAC1
FA91
FACA
FB29
FB50
FB47
FB54
FB79
FB6B
FB13
FAC6
FAD4
FB19
FB35
FB14
FAFC
FB12
FB30
FB3F
FB6A
FBC5
FBF2
FB8E
FAEA
FAC8
FB49
FB9C
FB2F
FAE3
FC55
FFD6
03A0
058E
0557
048C
0490
052C
0560
04F6
049D
04C2
0502
04EA
04B7
04EA
056D
05A6
0560
051C
054D
05B1
05B1
053C
04C7
049F
0493
0469
0449
0472
04C1
04D3
049C
0475
0498
04CE
04D5
04C8
04DD
04F3
04BA
0455
0456
04E8
055E
0507
0445
0432
0503
0547
035C
FF7C
FBCB
FA27
FA59
FAC6
FA7F
FA0B
FA3C
FAE5
FB34
FAEF
FAB5
FAFB
FB60
FB4A
FACE
FA8F
FACE
FB17
FAFF
FABE
FAC6
FB10
FB2D
FAFB
FAD0
FAEC
FB17
FB0A
FAF1
FB28
FB9B
FBD2
FBA0
FB62
FB64
FB69
FB28
FAE9
FB22
FBA4
FBB1
FB19
FAAB
FB17
FBC3
FB81
FA7F
FAA2
FD65
01C9
0526
05F4
0525
049D
04FD
0577
055E
050F
052A
0589
0595
053A
04FE
0529
055E
052F
04C3
0491
04B6
04DF
04D6
04C3
04D7
04EF
04DA
04B4
04BC
04E1
04C5
0455
0402
0436
04BA
0502
04E9
04D8
0512
0542
0504
0492
0488
04EF
051A
04AC
044D
04C3
0576
049F
015A
FD15
FA57
FA23
FB23
FB7A
FAD5
FA49
FA8A
FB1B
FB3F
FB0D
FB0C
FB3C
FB22
FAAB
FA64
FAAE
FB28
FB3D
FAFF
FAF9
FB54
FB9D
FB89
FB68
FB8D
FBB0
FB5C
FAC4
FA9F
FB1E
FB9A
FB76
FAFC
FAE5
FB43
FB71
FB1B
FAB9
FAD0
FB1F
FB14
FAC9
FAE4
FB74
FBA8
FB0A
FAA2
FC13
FF9C
0375
0587
0580
04CD
04C5
0560
05CB
05A5
054B
051A
04F9
04B8
047E
0498
04F9
0539
0526
0503
051E
0551
053B
04CA
045A
043A
0456
0475
0494
04D0
0508
04E8
0471
0428
047F
0530
0581
0524
048E
044E
046F
04A5
04D0
0503
051F
04F0
04AA
04DD
057F
0562
033C
FF58
FBB6
FA1C
FA60
FAF6
FADA
FA6A
FA6B
FAD9
FB18
FAEB
FAAF
FAAF
FABF
FAB0
FABE
FB2D
FBBB
FBE0
FB86
FB23
FB1A
FB4D
FB6D
FB76
FB92
FBB8
FBA6
FB54
FB10
FB18
FB3B
FB2C
FAF8
FAF4
FB3C
FB8E
FBB0
FBAC
FB97
FB5D
FAEF
FA99
FAC8
FB64
FBB4
FB43
FABF
FB91
FE5A
020A
04B6
0562
04C3
044A
04A0
0544
0578
0537
0505
0525
0552
0543
0512
04F8
04E6
04A5
0448
042A
0469
04AF
04A0
045E
0455
04A1
04EA
04F3
04EB
0508
0524
04FC
04A8
047C
0482
0470
0433
042B
04A1
0537
054F
04DF
047A
0477
0482
045F
0479
052D
05AD
0467
00E0
FCBC
FA55
FA68
FB8A
FBF4
FB54
FAA7
FAAE
FB24
FB62
FB36
FAEF
FAD0
FAD1
FADB
FAEF
FB12
FB28
FB18
FAFA
FB09
FB53
FBA8
FBC6
FBA4
FB6A
FB49
FB4A
FB55
FB4F
FB36
FB18
FB07
FB13
FB48
FB95
FBBF
FB93
FB2A
FAE1
FAEC
FB20
FB35
FB2F
FB45
FB78
FB76
FB2D
FB18
FBA5
FC5B
FC37
FB1E
FA84
FC12
FFBD
0397
05B1
05D7
054B
0521
0553
0555
0507
04BE
04B0
04C7
04E4
0505
051E
0514
04E9
04CC
04E3
0518
0535
0528
050C
04F6
04E5
04D9
04DF
04EE
04DB
0499
045C
0467
04B2
04FD
0518
0505
04DB
04AC
0489
048B
04B9
04F2
0506
04E7
04B5
0496
049F
04D2
0509
04F6
0479
0400
0433
04FE
0529
0360
FFC1
FC08
FA04
F9F8
FABA
FB24
FB1B
FB1D
FB57
FB7D
FB58
FB0B
FAD2
FABE
FAC3
FADE
FB06
FB20
FB1A
FB07
FB09
FB28
FB47
FB53
FB55
FB54
FB46
FB2C
FB24
FB44
FB71
FB7D
FB54
FB08
FAB7
FA8A
FAA2
FAF5
FB45
FB5B
FB48
FB4C
FB80
FBB0
FBAC
FB88
FB70
FB5B
FB35
FB39
FBB1
FC52
FC4D
FB7F
FB24
FCBF
004C
03F3
05CF
05B7
0507
04E3
0531
0549
0506
04CC
04D6
04FB
0509
0502
04F1
04D9
04CB
04DF
050C
0521
0508
04EC
04FE
0526
0524
04F6
04E6
0510
052E
04FB
04A1
0482
04BA
050F
0543
0547
0528
04F7
04CB
04B2
04A2
047F
0448
041F
041E
0430
044A
048F
050A
0551
04EF
0439
0428
04EF
053B
036D
FFA0
FBE0
FA23
FA67
FB1B
FB17
FAA0
FA88
FAEF
FB45
FB35
FAF8
FAE1
FAF1
FAF7
FAD9
FAA7
FA89
FAA3
FAEB
FB27
FB28
FAFE
FAEC
FB07
FB17
FAE8
FAA3
FAA8
FB01
FB48
FB39
FB03
FAF1
FAFF
FB03
FB06
FB34
FB7D
FBA2
FB8B
FB62
FB52
FB52
FB55
FB6E
FB96
FB83
FB18
FACC
FB26
FBC4
FB9C
FA93
FA46
FC6B
00A0
0484
0622
05CA
0534
0556
05AA
0579
04FC
04E0
052E
0556
0513
04BF
04BB
04FB
052F
0532
051A
050E
0522
054A
056A
0569
0549
052A
051F
050C
04CE
0482
046E
0498
04B6
04A6
04A4
04E2
052A
052A
04EF
04CD
04DB
04E2
04B9
0483
046C
046D
0479
04B3
0520
054E
04DB
0441
047B
0577
0591
0349
FF37
FBA8
FA40
FA87
FAF7
FAE0
FAC1
FB0B
FB60
FB42
FADE
FAC0
FAFB
FB29
FB17
FAF1
FAEA
FAF7
FB00
FB07
FB14
FB1B
FB16
FB13
FB20
FB35
FB42
FB51
FB6E
FB73
FB3A
FAE5
FAC3
FADA
FAD9
FAAD
FAB3
FB1C
FB82
FB66
FAF2
FABD
FAFB
FB4A
FB5B
FB60
FB96
FBBD
FB81
FB31
FB5F
FBCF
FB94
FAA3
FA8F
FCDD
00EF
046B
05B1
0551
04E7
0519
0556
051B
04BD
04B9
04EF
04F2
04C6
04C4
0500
0536
0544
0548
054D
0530
04ED
04BB
04C7
04F9
0514
0508
04F9
0504
0519
051C
050A
04E6
04BA
04AA
04D1
04FF
04DF
047F
0456
049F
04F4
04E5
04A3
04A5
04EA
04F6
04AA
0498
0518
058C
0532
0470
0472
0541
051B
027B
FE3F
FAEE
FA05
FAAC
FB2A
FAE8
FA8B
FAA6
FAFD
FB23
FB23
FB3C
FB63
FB6A
FB58
FB43
FB10
FAB0
FA70
FAA0
FB0F
FB3E
FB0D
FAE2
FB0D
FB52
FB4C
FB02
FADC
FB06
FB3A
FB37
FB1D
FB14
FB05
FADB
FABF
FADE
FB11
FB21
FB1F
FB37
FB4D
FB2C
FAF8
FB14
FB7E
FBAA
FB51
FB06
FB65
FBF2
FB95
FA78
FA82
FD3F
01B5
0529
05FD
051B
0478
04D6
0573
057E
051F
04F3
051C
053B
0515
04D0
04AF
04CE
051B
055A
054A
04F5
04B6
04C6
04E8
04CB
0485
047C
04CA
0513
050B
04E4
04FA
0538
0534
04E7
04C1
04F3
051D
04EB
049A
048D
04AC
04AA
049E
04D3
052B
052F
04DE
04D8
0561
05B7
051D
0435
045C
056C
0545
0247
FDAE
FA75
FA07
FB0E
FB7C
FAEF
FA7E
FACA
FB3A
FB23
FACD
FAE2
FB59
FB96
FB59
FAF8
FAC9
FAC9
FAD9
FAF1
FB14
FB33
FB43
FB4C
FB4F
FB3F
FB25
FB22
FB44
FB64
FB51
FB26
FB28
FB5A
FB6D
FB40
FB15
FB1D
FB2E
FB1C
FB0A
FB18
FB15
FAD8
FAAC
FAF6
FB7F
FB99
FB23
FAE5
FB6C
FBF9
FB72
FA5F
FADE
FE18
0278
0543
058C
04C0
0481
04DF
0504
04C4
04BD
0532
0599
057B
0524
0514
0533
0522
04EB
04E8
0520
0544
0533
051A
0514
04FD
04C8
04A7
04BB
04CD
049A
044A
0443
0491
04CB
04B9
04A4
04CF
0509
050B
04F4
0503
051C
04FE
04BE
04A8
04BA
04A4
0461
045F
04CC
051E
04D4
046F
04D2
0593
04E8
01D1
FDB4
FB07
FAA2
FB37
FB42
FAB1
FA5E
FA96
FAD8
FACC
FABC
FAEE
FB1E
FAF9
FAB4
FAB8
FAFC
FB2A
FB2D
FB32
FB3D
FB2F
FB11
FB11
FB2E
FB2A
FAF5
FAD7
FB13
FB77
FBA1
FB8B
FB86
FBA0
FB8B
FB34
FAFE
FB25
FB54
FB32
FAF6
FAFE
FB2C
FB26
FB02
FB38
FBC3
FBFF
FB8E
FB05
FB0C
FB44
FADB
FA4A
FB5B
FEE1
0333
05BC
05C7
04DE
049F
0511
0554
051F
04E9
04F4
04F0
04B1
0499
04F3
0569
0587
0563
0556
0555
051B
04BA
0491
04B4
04D7
04CA
04BA
04D4
04F1
04D6
049F
0497
04BA
04B8
0485
0476
04B0
04DD
04C1
04A3
04D0
0516
0521
050E
052E
055C
052B
049D
0447
0470
049C
045C
0434
04DA
059D
049E
011C
FCDA
FA64
FA62
FB50
FBA0
FB45
FB08
FB33
FB6C
FB77
FB81
FB9A
FB7C
FB10
FAB2
FAA6
FAB3
FA95
FA89
FADE
FB5E
FB8E
FB5E
FB2E
FB30
FB3B
FB2D
FB32
FB6D
FBA9
FB9E
FB65
FB52
FB63
FB44
FAE9
FAB9
FAE2
FB09
FAE7
FAC8
FAFD
FB4A
FB45
FB0F
FB1E
FB62
FB4C
FAC8
FA8D
FB0F
FB95
FB30
FA8A
FB95
FF1B
0351
05AD
05A0
04BD
0484
04F0
0534
0518
0503
052F
055C
055B
0549
053A
04FE
048E
0449
046C
04AE
04AD
0483
0485
04AE
04B6
0493
0483
049B
04A2
0479
045A
0483
04D6
0500
04F8
04FD
051A
050C
04C8
049E
04BA
04D9
04CE
04D3
050B
0515
049F
0419
043A
04E7
0532
04BC
0461
04EF
057F
0426
0078
FC83
FAA1
FAF3
FBB2
FB89
FAC7
FA60
FA90
FAE9
FB28
FB68
FBAF
FBBC
FB71
FB12
FAE8
FAE9
FAEC
FAF6
FB16
FB2C
FB22
FB1F
FB45
FB67
FB50
FB23
FB35
FB86
FBBC
FBA2
FB6D
FB64
FB77
FB61
FB1D
FAEF
FAF5
FB06
FB12
FB39
FB6E
FB67
FB24
FB0D
FB4F
FB72
FB1F
FAD7
FB51
FC31
FC2E
FAEA
FA0C
FBAE
FFBD
03CA
05AF
059C
052F
0538
0545
04F7
04C1
050D
0578
0559
04BC
0459
0496
050C
0530
0506
04ED
04FE
0508
04F6
04E3
04DD
04D3
04C7
04C9
04D7
04DA
04DA
04F5
052A
0547
0522
04CF
0492
0490
04B3
04D4
04EB
0503
0518
051D
0500
04C0
048B
04B3
0520
04DA
02BB
FEF2
FB59
F9DC
FA82
FB90
FB95
FAD7
FA7D
FAD1
FB14
FAD9
FAAB
FB08
FB7A
FB49
FAA1
FA5F
FACC
FB46
FB3D
FAF4
FAFB
FB4D
FB64
FB10
FABE
FAC1
FADF
FAC5
FA94
FA9E
FAD9
FB02
FB17
FB4A
FB87
FB7C
FB1D
FAD5
FAF5
FB47
FB64
FB57
FB86
FBE7
FBD3
FAFB
FA47
FB38
FE4D
0248
053A
0624
0599
04EB
04E1
053E
0563
0522
04D4
04C1
04CA
04BA
04A3
04C1
0510
053C
051C
04FB
052B
057F
057B
0513
04CB
0508
0581
05B1
0587
0558
054D
053F
0513
04F1
04FA
0506
04E5
04B9
04B9
04CA
04A6
045F
045E
04A7
04BD
047C
0487
054B
05CE
045A
008F
FC48
F9EC
FA09
FB1C
FB91
FB4F
FB26
FB5D
FB7E
FB4B
FB25
FB60
FBBB
FBBD
FB68
FB27
FB30
FB40
FB07
FAAA
FA91
FADE
FB41
FB57
FB0C
FA9E
FA5E
FA77
FAD6
FB37
FB5C
FB3F
FB12
FB11
FB47
FB8D
FBB1
FBA8
FB8B
FB66
FB27
FAD9
FAC8
FB2B
FBA8
FB8A
FABC
FA63
FBF8
FF97
0371
0573
0554
04A4
04CD
0596
05E6
0568
04DC
04DB
0519
04FE
049F
048A
04D2
04F3
04A0
0447
0468
04D7
04FD
04AB
0448
0435
046A
04B4
0501
0549
0564
053B
0502
04FE
0515
04EA
0474
042C
0468
04DD
0507
04E2
04DA
0503
04F5
0488
045E
051F
0639
05F5
032B
FEC1
FB0F
F9BD
FA6F
FB81
FBD2
FB82
FB3D
FB3E
FB36
FAEF
FAA1
FA96
FABA
FAC3
FAA3
FA99
FACA
FB07
FB1B
FB1A
FB3B
FB7E
FBA3
FB85
FB47
FB1E
FB06
FAE6
FACD
FADD
FB02
FB05
FAE4
FAE8
FB32
FB7A
FB7B
FB5A
FB70
FBB1
FBB6
FB6E
FB4C
FB8E
FBA8
FAFE
FA2F
FAEB
FE13
0256
054F
05DB
04FF
046D
04B6
053A
0566
055F
057A
0594
055A
04E9
04B2
04D6
0504
04FE
04F0
051D
0565
0572
053A
0515
0540
0588
058F
0549
04F7
04C8
04A9
0482
046A
047B
04A2
04BA
04CF
0504
0540
0535
04CE
046B
046B
04A8
04A5
045A
045D
04F5
053A
03C1
0050
FC86
FA6D
FA7E
FB5C
FB8D
FAF9
FA8B
FAC7
FB3C
FB55
FB20
FAFC
FAED
FAA8
FA3A
FA1D
FA94
FB3D
FB86
FB5E
FB31
FB3A
FB3E
FB02
FAB9
FAC0
FB11
FB4C
FB2F
FAD9
FA8B
FA62
FA6A
FAB3
FB2F
FB92
FB9A
FB72
FB84
FBE0
FC18
FBE6
FBA3
FBC1
FBF6
FB84
FA81
FA59
FC7A
0078
0425
05A5
0530
0476
0498
053B
0580
0543
0510
0537
056C
055F
053D
0557
0599
05A5
055D
050B
04F2
0502
050B
050A
051F
0542
0547
051F
04EA
04CA
04BD
04C3
04EA
0523
052A
04D4
046B
0469
04D6
0524
04E4
046A
045D
04C9
04FE
0495
0430
04A6
0596
054B
0291
FE52
FAEF
F9F2
FAB3
FB70
FB4C
FAD7
FADD
FB3E
FB4F
FAE3
FA81
FA8F
FAD5
FAEA
FACE
FAD0
FB04
FB31
FB37
FB38
FB45
FB33
FAE7
FAA3
FABA
FB13
FB4B
FB47
FB55
FB99
FBC0
FB84
FB3B
FB67
FBE9
FC09
FB81
FAEE
FAFB
FB61
FB55
FAC6
FA8C
FB11
FB82
FB01
FA45
FB37
FEA6
0301
05CC
061B
052E
04AF
04FC
0553
0533
04E6
04E2
051E
0549
0546
0534
0527
0511
04F7
04F8
0512
0518
04ED
04C1
04D0
0503
0501
04A4
043A
0420
044D
046B
0453
043D
045F
0495
0498
0474
0482
04E0
052E
0516
04D0
04D4
0518
0515
04AC
0480
04FA
053A
03B8
0026
FC48
FA4F
FAA1
FBA8
FBDB
FB3D
FABD
FAB2
FA9F
FA38
F9E1
FA09
FA7B
FAC1
FAD2
FB01
FB59
FB80
FB53
FB28
FB38
FB37
FAD0
FA58
FA74
FB30
FBDD
FBEA
FB8F
FB5C
FB69
FB64
FB35
FB28
FB5D
FB78
FB2F
FADA
FAFA
FB70
FBA3
FB69
FB52
FBC5
FC41
FBF6
FB1D
FB29
FD46
00DB
03F7
0535
04F3
0489
04BA
052F
0547
04FB
04C8
04F3
0547
0577
0588
05A0
05AF
058A
0544
0524
0534
0528
04D3
047D
048B
04E9
051E
04F3
04C1
04E8
0540
0554
0510
04CE
04C2
04B5
0482
046E
04B8
050F
04F6
0483
044A
0474
047B
040F
03D9
0499
05A0
0502
01CE
FD84
FAB1
FA57
FB38
FBA9
FB59
FB0B
FB1C
FB19
FAAD
FA3B
FA42
FA99
FAB7
FA8C
FA88
FAD7
FB14
FAE0
FA74
FA54
FA9A
FADF
FAD6
FAAB
FAB3
FAF3
FB2B
FB43
FB60
FB93
FBB3
FBA7
FB91
FB9C
FBAE
FB92
FB5B
FB5A
FB9F
FBC6
FB7A
FB0F
FB2C
FBC7
FBF9
FB31
FA68
FB6D
FED8
0305
05A2
05FB
0559
0533
058F
058D
04F8
0498
04F5
058C
0594
0527
0503
0569
05C4
058F
050F
04E1
0516
0534
0503
04D8
04FF
0541
0540
050C
04FA
0519
051E
04E8
04AD
0499
0489
0454
042B
0457
04AF
04BA
0468
0441
049C
0503
04D3
0448
044C
0508
0525
031E
FF2F
FB77
F9DF
FA45
FB00
FAED
FA70
FA76
FB0A
FB6F
FB3F
FAED
FB09
FB69
FB7F
FB29
FADC
FAEE
FB1E
FAF8
FA8A
FA4C
FA80
FAE9
FB26
FB2D
FB2E
FB38
FB30
FB0F
FAEA
FAD0
FABE
FAC3
FB04
FB76
FBC7
FBBA
FB81
FB7A
FBA6
FBA6
FB65
FB56
FBC1
FC20
FBB4
FADB
FB2D
FDD7
01F8
0535
060C
053A
0498
04FD
05A7
059E
0501
04A9
04F0
0554
054E
0505
04F7
0532
054F
0514
04C5
04C1
0502
0533
0523
04F1
04C8
04AE
049C
049E
04B8
04D1
04D3
04CB
04CA
04BA
047E
0437
043C
04A1
0504
0507
04D2
04D1
0505
04EF
046C
041E
0497
052A
043B
010D
FCED
FA23
F9B3
FA91
FB12
FAB2
FA2E
FA35
FA9B
FACF
FAB4
FAA2
FAC7
FAEF
FADE
FAAD
FA9A
FAB8
FAE6
FB0A
FB22
FB2C
FB1E
FB02
FAFA
FB18
FB48
FB70
FB8F
FBB1
FBC5
FBB4
FB91
FB93
FBCC
FBFE
FBE1
FB84
FB37
FB1E
FB09
FAD6
FABE
FB02
FB59
FB26
FA69
FA44
FC09
FFAE
037D
059D
05C1
052B
0516
0586
05C0
0577
051E
052A
0580
05BF
05C8
05C2
05B6
057C
051B
04DB
04E6
0505
04F9
04D8
04E4
0518
0529
04F7
04BA
04AA
04B5
04B0
04AC
04CD
04EB
04B3
043A
0411
0486
0524
0547
04FA
04D9
051F
0547
04E9
0484
04D7
0583
0502
0257
FE7E
FB98
FACA
FB4D
FBA0
FB2F
FA8D
FA5F
FA96
FAC1
FAB5
FA9D
FA94
FA86
FA74
FA8B
FAD8
FB1B
FB16
FAE5
FADB
FB0B
FB2F
FB10
FAD7
FAD3
FB0F
FB48
FB56
FB51
FB4B
FB1D
FAB2
FA54
FA68
FADB
FB2F
FB2C
FB35
FBA5
FC1A
FBDF
FB04
FA7E
FAE5
FB84
FB48
FA89
FB0B
FDF0
020D
0500
05A8
0505
04AA
04F5
053A
051C
0507
054A
0589
0555
04EC
04DC
0524
053B
04E7
0495
04B4
0514
053B
051F
051D
0558
057D
0552
0511
0501
04F3
049C
042E
0432
04B0
0504
04B9
043B
0445
04CF
0516
04CE
04A9
0545
05D4
04A9
0141
FD39
FAD0
FA9E
FB4B
FB61
FADD
FAB7
FB49
FBE0
FBCC
FB4C
FB15
FB4B
FB6A
FB22
FACB
FAD5
FB2C
FB62
FB51
FB35
FB30
FB1E
FAEB
FAD1
FB00
FB48
FB59
FB42
FB5C
FBA8
FBBC
FB60
FAFD
FB06
FB4C
FB48
FB02
FB19
FBB6
FC11
FB81
FAD8
FBD9
FF20
0311
056C
059C
04F7
04DE
0548
0558
04D1
0454
045E
04A5
04AB
047E
047E
04B5
04CC
049E
0476
0493
04C9
04C9
049E
0490
04B7
04DD
04E4
04F0
0511
050D
04B2
0448
044E
04CB
0538
0530
04F2
04EF
0515
04F9
04A9
04BD
0559
056B
0398
FFEF
FC43
FA79
FAB8
FB93
FBC6
FB59
FB03
FB02
FB03
FAD5
FAC0
FAFA
FB42
FB3F
FB03
FAF1
FB27
FB5F
FB67
FB67
FB8F
FBB6
FB9C
FB54
FB37
FB58
FB70
FB4C
FB24
FB3D
FB77
FB76
FB33
FB06
FB14
FB18
FAEA
FAE6
FB5F
FBE2
FB9E
FABB
FAB9
FCF0
00CC
041C
0543
04BB
042D
0476
050F
052F
04D9
0498
0495
0487
0452
0444
0495
04FD
0520
050C
050E
052D
0523
04DE
04A9
04BD
04E8
04DF
04BA
04C5
04F9
04F5
04A1
0469
04A1
04F3
04D6
0468
0456
04D5
053F
0506
04A9
0509
05D0
054E
025B
FE10
FAE9
FA40
FB22
FBBE
FB66
FAD1
FAB7
FAF1
FB07
FB02
FB36
FB90
FBA3
FB54
FB10
FB2B
FB67
FB60
FB27
FB21
FB5B
FB76
FB3F
FB05
FB12
FB30
FB06
FABE
FAD9
FB5E
FBA8
FB4F
FAD4
FAFA
FBA1
FBEE
FB85
FB15
FB3F
FB84
FB07
FA39
FADC
FDF4
022E
050A
0574
04A2
0451
04D1
0549
053F
0528
056D
05AE
0567
04CE
048B
04C2
04F0
04C7
04A9
04FA
0568
055D
04E5
04AD
0506
0571
055E
04F7
04CE
04F6
04F9
04A4
046C
04AD
0513
051A
04E7
0501
055F
054C
0491
0415
04A5
0567
045F
00D9
FCAC
FA6F
FABE
FBE0
FC05
FB2B
FA84
FA9F
FAEF
FAF0
FAEB
FB4C
FBC7
FBC3
FB49
FB02
FB31
FB55
FAF0
FA5B
FA4A
FAC6
FB22
FAEE
FA89
FA87
FAE1
FB26
FB33
FB49
FB7D
FB84
FB3E
FB01
FB1B
FB42
FB03
FA96
FAA7
FB36
FB5A
FA9C
FA2F
FBE9
FFF2
0419
05F8
056C
0464
046D
0532
0584
0524
04DC
0520
0574
0541
04C6
04A4
04EA
050D
04CA
0487
04AE
0507
051A
04E6
04CC
04ED
04FD
04D2
04B2
04DF
051E
050C
04CA
04D6
0546
0592
055C
04FD
04F9
0526
04FB
0494
04B6
0579
0580
0344
FF22
FB6A
FA0D
FAB2
FB7E
FB5C
FADA
FAD8
FB36
FB33
FAB5
FA65
FAAA
FB0F
FB03
FAAB
FA97
FAE3
FB2B
FB38
FB4B
FB8F
FBB6
FB6D
FAF6
FAD5
FB0E
FB1E
FACC
FA8F
FAD6
FB4B
FB44
FAC5
FA82
FADA
FB49
FB3E
FAF4
FB08
FB5F
FB40
FAB9
FB2A
FDC5
01C2
04DB
05A2
04DD
0450
04AB
053C
0559
0543
056B
0598
054B
04B8
049D
052E
05B2
057E
04DD
0497
04D7
050A
04DE
04BE
0517
0595
0592
0515
04C7
04FD
0542
0516
04B3
04A5
04EF
050B
04D3
04BF
0510
0543
04D6
0440
0467
0518
04B9
021A
FE26
FB28
FA5E
FAE3
FB23
FABA
FA6A
FAA1
FAED
FADB
FAC0
FB15
FB91
FB74
FAB4
FA32
FA89
FB40
FB72
FB0C
FAC4
FB00
FB4C
FB24
FABF
FAB4
FB0E
FB40
FB06
FAC8
FAF0
FB46
FB4F
FB10
FAF9
FB26
FB3B
FB10
FB07
FB5D
FB8B
FB01
FA66
FB63
FEAD
02CD
0565
05A1
04CB
0488
050B
0573
0559
053E
0585
05BA
0555
04A9
0486
0510
0587
0554
04CC
0499
04C6
04D3
0497
0482
04DE
054B
0544
04DB
0497
04A3
04A7
0470
044D
0493
0505
052B
0507
04FF
0522
0502
0485
0455
04E3
0546
03E1
0060
FC8A
FA96
FAD8
FBAD
FB97
FACD
FA6A
FAB8
FAF7
FA9E
FA1F
FA2A
FAAC
FB05
FB00
FB08
FB64
FBBE
FBA7
FB41
FB07
FB23
FB4B
FB56
FB73
FBC2
FBFC
FBCD
FB55
FAFC
FAE8
FADD
FAC7
FAE6
FB4B
FB8D
FB51
FAF6
FB24
FBC1
FBE2
FB30
FADC
FC92
0061
0446
062A
05E9
0515
04F4
055A
0579
0528
04EA
04FF
0513
04DA
0492
049D
04EB
051D
0512
04FF
0500
04F6
04D1
04BF
04D8
04E3
04A3
0451
045C
04C2
04F7
04AA
0446
045E
04D5
0506
04BD
0481
04BB
0503
04C6
044E
0479
053B
0512
029B
FE74
FAF0
F9C2
FA72
FB40
FB34
FAC0
FAA4
FAE4
FB07
FAF3
FAEC
FB0A
FB0E
FADF
FAC0
FADF
FB03
FAE5
FAB7
FAE3
FB5B
FB8F
FB31
FAB3
FAB3
FB24
FB71
FB58
FB3D
FB7C
FBD2
FBC5
FB63
FB32
FB64
FB97
FB7E
FB60
FB8D
FBA9
FB29
FA80
FB2E
FE18
022A
0524
05DB
0539
04DA
053B
05A3
0584
053B
054C
0585
0555
04BF
0467
04A5
050A
050C
04C6
04B5
04EE
0505
04CB
04A2
04E5
054D
0549
04CF
0475
04A1
0500
050D
04C1
0487
0490
04AC
04B1
04B4
04BC
0493
0435
0424
04BE
054B
0449
011D
FD1A
FA66
F9DA
FA6E
FABC
FA89
FA84
FAF0
FB3C
FB00
FAAF
FAE5
FB73
FB90
FB00
FA72
FA95
FB38
FB9A
FB6A
FB08
FAE2
FAE9
FADE
FAC6
FAD5
FB0A
FB32
FB40
FB60
FB9E
FBCA
FBC5
FBB1
FBB0
FB9A
FB4D
FB15
FB63
FBF9
FBFD
FB2F
FAC6
FC68
002B
0413
05F6
0592
047E
0434
04B2
051D
051B
050B
052E
0542
050B
04D3
04FF
0569
0586
0528
04BD
04B6
04F7
0514
04EE
04C7
04CF
04E3
04D7
04B3
049B
0490
0486
048B
04AF
04D0
04B9
047D
046F
04A3
04B3
0455
03F3
0442
0518
0524
0332
FF9F
FC3C
FA96
FA9C
FB1B
FB31
FAEE
FABE
FAB1
FA99
FA7E
FA9E
FAFC
FB47
FB42
FB17
FB15
FB43
FB68
FB60
FB41
FB1D
FAED
FABA
FAB4
FAFC
FB63
FB9C
FB9C
FB9B
FBAD
FBA3
FB63
FB33
FB5C
FBAF
FBAF
FB57
FB39
FBA7
FC07
FB88
FA8D
FAC6
FD6C
01A0
050B
062B
0599
04EE
04DF
04E8
0490
0440
0495
0558
05BA
056B
04FB
04FB
053C
0533
04D2
048C
0499
04A8
0471
043A
046A
04DB
04FF
04A8
044B
0456
04A0
04B8
0499
0497
04C4
04C8
0484
045B
0498
04DB
0496
040E
041D
04CB
04AA
024B
FE32
FABB
F9B8
FAA9
FBA0
FB8A
FB01
FAF5
FB58
FB6C
FAFB
FA93
FAA8
FAF8
FB0C
FAEB
FAF0
FB34
FB73
FB89
FB95
FBA7
FB8B
FB34
FAFF
FB4A
FBDB
FC18
FBD6
FB86
FB76
FB59
FADB
FA68
FABB
FBAE
FC1A
FB60
FAA2
FBCA
FF48
0350
05A6
05D1
0522
04DF
050D
050C
04C6
04B1
04FA
053E
0531
050D
0521
053A
04F4
0471
0449
04B1
051B
04F2
0465
0429
047B
04D3
04B0
0445
0423
045D
0481
0459
043B
0473
04BB
04A6
0470
04BE
0578
055C
033F
FF96
FC4D
FAE1
FB00
FB44
FAEF
FA7F
FA9A
FAFF
FAF5
FA63
F9FB
FA44
FAE8
FB36
FB0C
FAE2
FB04
FB37
FB34
FB24
FB57
FBB3
FBCB
FB83
FB48
FB78
FBDA
FBF6
FBBD
FB8C
FB84
FB61
FB04
FAD8
FB37
FBAA
FB5F
FA83
FAA1
FD18
014C
04EA
0626
0568
047F
0495
0546
05A3
0570
0528
0524
053F
0540
0531
052C
0518
04DA
049B
0496
04B1
049C
0453
0434
0477
04CC
04C5
0476
045E
04A3
04CE
0487
042B
0454
04E5
051D
04B3
045E
04D4
0578
04A9
01A3
FDAB
FAE8
FA48
FAD8
FB26
FAD4
FA88
FAB7
FB11
FB13
FAC6
FA96
FAB0
FADC
FAEE
FB01
FB2F
FB4F
FB39
FB17
FB3B
FB9D
FBD3
FB97
FB2C
FB02
FB27
FB53
FB68
FB94
FBD6
FBC7
FB2B
FA87
FAA7
FB72
FBD0
FB18
FA5D
FB9B
FF5E
03BE
0621
05DC
049E
044E
0509
0599
054C
04B9
04AF
0516
0545
0510
04E6
0501
0509
04B5
0459
0475
04E5
0507
04A1
0436
0448
04A8
04D4
04C0
04D1
0519
0522
04B7
0459
0490
0507
04F3
045A
042C
04D2
050B
0324
FF32
FB6E
F9F3
FA8F
FB5C
FB22
FA78
FA80
FB32
FB94
FB2E
FAA2
FAAE
FB2B
FB6C
FB3E
FB0F
FB2B
FB57
FB41
FB06
FAF6
FB19
FB39
FB44
FB5A
FB67
FB24
FA9A
FA5D
FADF
FBB0
FBEB
FB63
FAF3
FB50
FBF7
FBD2
FAF9
FB14
FD94
01C8
0549
0663
05A1
04D4
04F7
057C
057D
04F7
0497
04AE
04DB
04C5
049A
04BD
051C
054D
0522
04E3
04DC
04F4
04EA
04C5
04C5
04F9
0523
0513
04EB
04D9
04CA
0497
0462
0471
04A6
048A
040E
03DD
0483
053E
0456
010A
FCCD
FA16
F9F2
FB19
FBA4
FB1C
FA88
FABE
FB5D
FB91
FB3C
FAEF
FAFA
FB10
FAEA
FAC4
FAE6
FB18
FAED
FA76
FA47
FAAE
FB49
FB8F
FB77
FB52
FB37
FAFD
FABA
FADA
FB6D
FBDD
FBAA
FB33
FB40
FBCB
FBE4
FB1F
FAAF
FC53
0021
040E
05EE
05A0
04C7
04B2
0524
0536
04C7
0484
04CA
052E
052B
04DE
04BD
04E2
0506
0500
04FD
0512
050C
04D0
04AC
04F1
0566
0571
04F0
046F
046F
04AD
0496
0433
042F
04CC
0559
0516
0468
046D
0549
0575
034C
FF2D
FB6C
FA00
FA9B
FB68
FB3F
FAA2
FA89
FAF8
FB26
FAC4
FA68
FAA4
FB2F
FB5C
FB0C
FACB
FAF7
FB46
FB4A
FB17
FB10
FB46
FB62
FB3F
FB23
FB4A
FB7A
FB5A
FB0E
FB03
FB40
FB4A
FAF1
FABA
FB12
FB74
FB05
FA1A
FA78
FD73
0206
0580
063F
0533
0473
04D6
0572
0551
04BA
0492
0504
056C
055F
0532
053D
0541
04D6
0437
040D
0480
04F6
04DF
046E
043C
0478
04C7
04E4
04E8
04F2
04DA
0497
047F
04DD
0556
0545
04BA
049D
0561
05F9
04AD
0124
FD12
FAA1
FA55
FAEB
FB10
FAB0
FA7B
FAB5
FAF2
FADE
FAB2
FACC
FB1F
FB53
FB4D
FB3D
FB3C
FB25
FAE5
FABD
FAF2
FB6B
FBC3
FBCA
FBA5
FB7C
FB48
FB0B
FB04
FB5D
FBC0
FB9B
FAEA
FA6C
FAB7
FB57
FB44
FA6C
FA3E
FC4C
005A
0446
0609
059A
049D
0478
0516
0590
0574
051E
04FF
050F
050F
04F7
04E9
04DA
04A9
0476
048F
04F5
053A
0508
049E
047F
04BF
04EF
04CB
0494
049F
04C5
04AC
046F
048B
050B
053F
04BC
042B
0486
057D
054B
02A0
FE6B
FB1E
FA2F
FAD1
FB47
FAF1
FA87
FAB0
FB1A
FB21
FAC9
FA98
FABD
FAE6
FAE5
FAFE
FB59
FB99
FB5A
FADC
FAC0
FB28
FB88
FB6F
FB21
FB14
FB36
FB1A
FACE
FAE4
FB80
FBE7
FB77
FAB9
FAC5
FBAB
FC1D
FB33
FA09
FAD1
FE47
029E
0556
05BA
0513
04CC
0500
050C
04CC
04BB
0511
0562
054A
0503
0504
0548
055E
051C
04D9
04DF
04FA
04DB
04A0
04AE
0503
0523
04D1
047E
04B1
0536
0552
04D0
045F
049F
052A
0520
0481
0454
051F
05B2
0434
006A
FC55
FA3E
FA6B
FB38
FB3D
FAB0
FA88
FAF6
FB44
FB03
FAA8
FAC3
FB2C
FB50
FB18
FAFE
FB3A
FB63
FB19
FAA7
FA9F
FB05
FB4E
FB32
FB0C
FB35
FB70
FB52
FAFF
FB01
FB5D
FB67
FACC
FA47
FAB7
FBB5
FBE8
FAEF
FA6E
FC5D
008B
047C
05FF
055B
0491
04D8
0596
05B4
0527
04BF
04DA
0504
04D4
0487
048B
04C7
04D1
049F
048E
04C6
04FA
04E9
04C1
04CA
04E7
04CD
049A
04C5
055C
05B8
0553
0493
0457
04C9
0529
04F3
04B3
052D
05EE
0551
0257
FE16
FAD7
F9DC
FA59
FABE
FA83
FA55
FAC7
FB73
FB98
FB23
FAC3
FAEF
FB5B
FB7B
FB45
FB26
FB55
FB90
FB87
FB52
FB30
FB29
FB13
FAEF
FAF0
FB21
FB3D
FB1F
FB04
FB31
FB70
FB4D
FADC
FABE
FB2B
FB6A
FAD1
FA1F
FB25
FEA9
0315
05D8
0600
04FD
04AB
0547
05B3
0547
049B
0480
04D4
04E7
0495
046C
04C1
0521
0506
0494
045E
0495
04DD
04F2
04F8
050C
04F2
0482
0428
046E
051A
054A
04A9
0408
0450
0538
0596
0505
047C
04CD
0518
0399
FFF9
FC25
FA50
FAA6
FB75
FB69
FAD4
FABA
FB41
FBAC
FB87
FB35
FB2B
FB43
FB1F
FAD2
FABF
FAEF
FB02
FAD5
FAC0
FB11
FB89
FBB6
FB8F
FB69
FB63
FB3C
FAE8
FAD0
FB3D
FBB9
FB93
FAEB
FAB3
FB69
FC36
FBE7
FAAC
FA58
FC87
00B3
0485
0614
0585
0478
042E
0495
04EF
04E4
04B9
04BB
04D5
04D3
04BC
04C6
04F8
051E
0515
04F2
04D5
04BE
04A6
04A2
04C9
0500
050C
04E1
04B3
049F
0481
0440
041F
046E
04F4
050E
049D
0458
04DC
0579
0495
0189
FDAC
FB1B
FA97
FB09
FB24
FADC
FAF1
FB85
FBDE
FB7F
FAE3
FAC6
FB1C
FB3E
FAF7
FACC
FB24
FB98
FB8C
FB14
FADD
FB2D
FB85
FB60
FAF4
FADA
FB2D
FB70
FB57
FB31
FB59
FB9E
FB93
FB51
FB5D
FBBF
FBC3
FB03
FA71
FBAE
FF23
0330
059D
05C4
04EA
0498
0507
0564
0527
04B1
0497
04D4
04EF
04C6
04AD
04E2
0522
050B
04AC
0482
04D2
054E
0573
0523
04BC
049A
04B3
04C9
04D0
04E8
050B
0504
04CD
04C3
0525
055B
0434
012A
FD54
FAA5
FA14
FACA
FB42
FAF7
FA97
FAC3
FB24
FB11
FAA1
FA8F
FB24
FBBA
FBA6
FB20
FAE9
FB33
FB6D
FB23
FAAA
FAA3
FB17
FB76
FB5F
FB11
FAF5
FB01
FAE5
FAA3
FA9B
FAF0
FB34
FAFB
FAA1
FB3F
FDA0
013C
046D
05D3
0585
04C9
04B4
0536
058F
056F
0545
057A
05BD
057A
04C5
045A
049D
0510
0515
04CD
04DA
0552
0594
0534
04AB
04AF
0528
0555
04F0
0496
04D0
0534
050D
048F
04B1
05A0
05F8
0419
0027
FC36
FA53
FA9C
FB83
FBAB
FB15
FA98
FAA3
FAE3
FAE3
FAA7
FA89
FAB3
FAF8
FB26
FB40
FB55
FB49
FB01
FAAF
FABC
FB37
FB9B
FB5F
FAAF
FA4C
FAA0
FB33
FB54
FB0F
FB0C
FB73
FB83
FAAD
F9E2
FAF8
FE91
02F8
0598
0592
0465
0408
04CE
058C
0568
04DC
04CE
053C
0565
04F3
047C
04A0
0527
055C
0509
04B3
04C9
0514
051C
04E1
04CF
050C
0540
0523
04ED
04F6
0521
0507
04A5
048B
0511
059A
04EB
026D
FEEF
FC0E
FAD9
FB06
FB77
FB5F
FAE1
FA9B
FACD
FB11
FAF9
FAAB
FAAA
FB0C
FB50
FB1A
FAB7
FAAD
FAF7
FB10
FACA
FA9B
FAE7
FB4F
FB31
FAAB
FA83
FAFC
FB62
FB1F
FAAF
FAEF
FBA4
FBAA
FABD
FA6D
FC7E
0095
0440
0586
04D8
0422
0472
052D
055C
04FA
04AD
04C9
0504
050D
0506
0535
0588
05A7
0563
04F1
04AA
04B1
04E8
0518
0529
052E
053B
0541
0520
04EE
04DF
04EF
04D3
0472
043B
0496
04FC
0413
011D
FD30
FA76
FA08
FAE7
FB52
FAC6
FA34
FA7C
FB42
FB91
FB23
FAA0
FAA5
FB0B
FB47
FB2C
FAFD
FAEE
FAEA
FADC
FADD
FAFF
FB22
FB22
FB12
FB24
FB4E
FB48
FB03
FADF
FB39
FBCD
FBD9
FB1D
FA86
FB89
FEA1
0291
0559
05FB
053C
04A5
04EC
057E
0583
04F9
04A0
04EB
056C
0570
04F3
04A2
04EA
056B
057A
050C
04BB
04EB
053E
0524
04B0
047E
04C9
0516
04E5
0473
0459
04A6
04D1
04A2
049E
0511
0508
030B
FF0E
FB19
F96C
FA34
FB8C
FBBC
FAE5
FA51
FAA1
FB3A
FB54
FAFB
FAC6
FAED
FB25
FB2E
FB26
FB34
FB36
FB00
FAAE
FA92
FACC
FB1B
FB32
FB13
FB03
FB28
FB5F
FB78
FB7E
FB96
FBA5
FB5C
FAC7
FABD
FC5E
FFCE
0396
05C3
05CA
04F5
04CD
056A
05B0
0505
042D
043A
0517
05AD
055E
04B4
047F
04BF
04E5
04C2
04B5
04EA
0508
04C5
0474
049D
052F
0587
0546
04D4
04BB
04E1
04C3
0456
0444
04ED
0584
048D
0171
FD6A
FA9A
FA1C
FB0D
FBA9
FB28
FA51
FA3C
FAF5
FB8A
FB5A
FACC
FAAF
FB21
FB89
FB74
FB1E
FAF5
FB01
FB06
FB01
FB29
FB75
FB8A
FB40
FAEA
FAEB
FB2C
FB48
FB2E
FB41
FBAA
FBE5
FB65
FAA2
FB02
FD74
013F
0475
05B6
0552
04B5
04D6
056C
05A4
0547
04DC
04D4
04FC
04E9
04A8
04A9
0508
054E
0511
0495
0477
04DA
053C
0530
04E9
04CC
04CA
0493
043E
044A
04D6
053A
04DA
0423
042E
052A
05AC
03FC
001C
FC0B
F9E6
F9FF
FAEB
FB3B
FAC7
FA5B
FA86
FB01
FB40
FB20
FAF0
FAF3
FB22
FB60
FB9C
FBBD
FB99
FB2D
FAD1
FAE7
FB59
FBA4
FB72
FB10
FB03
FB51
FB7E
FB4A
FB1E
FB6C
FBE2
FBB3
FAC5
FA43
FB9F
FF08
02F8
0582
05F6
053D
04BA
04FA
0578
057E
04FF
048F
04A0
04FB
0522
04F9
04D9
04F8
0516
04E7
0489
0456
045A
0450
0428
043B
04BB
053A
0525
0498
044A
0486
04C1
048A
0456
04DB
05A6
051A
0237
FE0B
FADC
F9F2
FA8B
FB17
FAF8
FAB5
FADC
FB3F
FB62
FB2D
FAF5
FAF5
FB10
FB1A
FB1C
FB3F
FB79
FB93
FB76
FB58
FB74
FBB3
FBC0
FB7F
FB3B
FB42
FB77
FB70
FB1D
FB00
FB72
FBED
FB92
FA8A
FA63
FC94
00AE
047F
0629
05C9
04F0
04C3
0516
0535
0500
04DA
04EC
04EC
04B3
048B
04C5
0534
0557
0501
0491
0472
049A
04A7
0475
044D
0475
04BE
04C3
047C
0451
0486
04C9
049F
042E
043C
050B
0587
041B
008D
FC97
FA5C
FA57
FB29
FB54
FAB9
FA48
FA93
FB34
FB82
FB64
FB36
FB2D
FB2C
FB1E
FB23
FB48
FB61
FB47
FB22
FB39
FB89
FBB3
FB6F
FAFC
FAD8
FB2D
FB96
FBA8
FB84
FB98
FBE3
FBCA
FAF1
FA2D
FB14
FE52
0294
058E
062B
0561
04D0
04F3
0519
04C8
047E
04DA
058F
05BC
0525
0482
047F
04DC
04E8
0487
0442
046B
04AC
049C
046B
048E
04FD
052C
04CF
045D
0474
04F5
051E
04A4
043A
04AD
0594
0558
02CC
FEA7
FB16
F9BF
FA52
FB35
FB4C
FADB
FAB3
FB01
FB3D
FB05
FA9D
FA7D
FAB4
FAF0
FB04
FB13
FB3E
FB67
FB6A
FB5F
FB71
FB8D
FB77
FB27
FAEA
FAFA
FB2E
FB35
FB0A
FB0A
FB6B
FBC3
FB78
FAAB
FA92
FC6E
0019
03D2
05BD
059B
04D1
04C2
0565
05BB
0554
04D2
04E7
055A
056F
0503
04AE
04DA
052B
051D
04C6
04A9
04DF
04F1
049B
044E
048C
051C
054E
04F7
04B4
04FD
056E
054A
0498
043F
04D3
0578
0481
0147
FD23
FA52
F9DF
FAD1
FB70
FB13
FA7A
FA81
FAF0
FAF5
FA6A
FA15
FA87
FB47
FB77
FB02
FAA3
FADC
FB58
FB8B
FB78
FB80
FB99
FB59
FAC6
FA8E
FB14
FBC4
FBC6
FB33
FAF2
FB5E
FBAC
FB14
FA40
FAED
FDF7
021E
0523
05DF
051B
045B
045C
04C8
050B
050B
050E
0534
0557
0554
0549
055B
0564
0524
04A8
045A
047A
04CB
04DE
04AE
049C
04D0
04ED
0496
041E
042E
04CE
0536
04DA
044C
047E
054C
053A
0307
FF3B
FBCE
FA46
FA79
FB27
FB64
FB35
FB07
FB0A
FB23
FB31
FB36
FB3C
FB3F
FB37
FB23
FB10
FB10
FB2A
FB4D
FB5B
FB48
FB2B
FB2A
FB4B
FB75
FB8E
FB8A
FB66
FB2B
FB0D
FB45
FBB6
FBD8
FB63
FB00
FC01
FF00
02E7
05AF
0641
055F
0496
049A
04EE
04F4
04CB
04E8
053D
054A
04ED
04A5
04D1
051C
04F5
046B
042A
0486
0500
04F6
0489
0463
04B8
0501
04C8
045D
0452
04A4
04CD
04A4
04A9
0521
0556
0426
0157
FDFC
FB77
FA58
FA4A
FABC
FB3C
FB77
FB4C
FAF5
FADE
FB1F
FB5E
FB3C
FAD6
FA9F
FACF
FB31
FB76
FB8A
FB84
FB73
FB60
FB51
FB3C
FB11
FAF7
FB2C
FB98
FBC4
FB72
FB13
FB27
FB65
FB02
FA22
FA61
FD24
0190
0501
05DA
0518
04B7
053C
0599
0523
0487
049E
0525
0542
04E0
04B8
050B
0538
04D4
0462
0482
04E8
04E3
047D
045C
04B0
04E8
04AC
0472
04B6
051F
0510
04C8
0504
057A
0495
0170
FD5E
FAB7
FA4E
FAE3
FB08
FAB7
FABD
FB3E
FB92
FB5B
FB0B
FB21
FB6E
FB7C
FB46
FB1A
FB11
FB0F
FB1E
FB5E
FB99
FB79
FB14
FAF7
FB5B
FBBC
FB94
FB36
FB52
FBBD
FB80
FA7C
FA44
FC8B
00DF
04C4
063A
059A
04BB
04B7
0521
053C
050B
04FA
050B
04ED
049D
0471
0484
0496
0485
0486
04BB
04E1
04BB
0486
04A1
04E1
04BE
043A
0404
0474
04F1
04D7
0482
04B8
051E
0422
00EF
FCEB
FA79
FA65
FB41
FB66
FACF
FA7C
FAC3
FB0D
FAF8
FAD7
FAFC
FB2A
FB16
FB02
FB4A
FBAF
FB9F
FB2B
FB0C
FB80
FBE0
FBA7
FB41
FB46
FB73
FB29
FAA2
FABD
FB83
FBD1
FB1F
FAE3
FD17
016D
0532
064F
0581
04E3
0529
055C
04DE
046B
04C4
056D
0572
04E2
04A8
0513
0563
050C
0493
04A2
04FC
04F4
0497
047C
04BE
04E1
04BD
04C7
0530
0554
04BA
0411
0459
050F
0442
00FC
FCD3
FA47
FA0A
FAAF
FAD6
FAA2
FAD7
FB67
FB8E
FB15
FAA3
FAC0
FB20
FB3B
FB0C
FAE7
FADF
FADD
FAFA
FB4F
FB8D
FB4F
FAC9
FAA8
FB1B
FB76
FB2E
FAC3
FB0D
FBCD
FBD5
FAF9
FAEC
FD62
01AE
0522
05F2
04F2
0433
0486
0516
0516
04DD
0515
0593
05A4
052A
04C0
04CE
0516
0536
0530
0531
0525
04E5
04A0
04AC
04EF
04F8
04BA
04AC
04FB
0525
04CD
0488
050D
05B7
04B5
0133
FCD0
FA24
F9FE
FAD3
FAFC
FA91
FA9F
FB4B
FBA8
FB3D
FAAF
FABE
FB32
FB54
FB03
FAC2
FACF
FAE0
FACE
FAE7
FB45
FB77
FB3A
FB0C
FB68
FBDC
FB94
FAB0
FA3E
FAAD
FB13
FAAE
FA8D
FC90
00BC
04A5
0613
0574
04D9
053E
05C2
057B
04D8
04C8
053C
055F
04F0
049A
04E0
055A
056B
0523
04E7
04C3
0488
045A
0480
04D1
04E2
04BB
04D4
053E
0563
04F3
04A7
053A
05E2
04BB
0126
FCF9
FAA0
FA8C
FB31
FB36
FACD
FABA
FAF9
FAF0
FA8C
FA69
FACF
FB41
FB3F
FAFB
FAE2
FAF1
FAE9
FAEB
FB45
FBC1
FBCD
FB56
FB07
FB4E
FBAA
FB66
FAC6
FAB4
FB44
FB66
FA95
FA2C
FC15
0044
0457
060E
0592
04C1
04BF
0508
04CD
0460
0496
0564
05D3
0559
048E
0459
04D4
0559
056C
0525
04D1
0495
0486
04B5
04FF
0515
04E8
04C5
04D3
04C6
0473
0457
04F7
05A8
04C3
017E
FD4B
FA9C
FA55
FB20
FB60
FB03
FAF2
FB67
FBB4
FB73
FB19
FB21
FB4E
FB2E
FAE4
FAED
FB3D
FB51
FB12
FB04
FB4E
FB55
FAC0
FA42
FAA5
FB89
FBDC
FB72
FB36
FB97
FBB8
FAEC
FA6D
FC51
00A4
04BE
0620
052C
0439
0482
0526
050C
047B
0469
04EC
0535
04E1
047A
048A
04DA
04F5
04E5
04F1
0507
04ED
04C0
04C7
04EA
04DB
04AD
04C4
0510
04FE
0469
042B
04FC
05E9
04E8
0149
FCE9
FA58
FA38
FB10
FB60
FB17
FAE1
FAF3
FAFB
FAED
FB19
FB82
FBB9
FB87
FB4B
FB51
FB53
FAFE
FAA5
FAD9
FB76
FBBB
FB5B
FAED
FB01
FB3F
FB05
FA8D
FAB2
FB7A
FBCB
FB12
FAA4
FC72
007E
0467
05F2
0555
0491
04D9
0583
0578
04D4
0487
04D9
051D
04D2
0458
0453
04C4
051F
050B
04BB
048A
049D
04E5
0537
054C
04F5
0479
0460
04B6
04E3
0493
046A
051F
0605
0535
01BA
FD21
FA29
F9E6
FAED
FB62
FB07
FACD
FB21
FB7C
FB78
FB64
FB97
FBCB
FB99
FB32
FB0F
FB24
FAFB
FA9E
FAA6
FB39
FBA2
FB5F
FAFC
FB3D
FBDC
FBF3
FB6A
FB1C
FB62
FB5D
FA7B
FA12
FC33
00CA
050A
0665
054B
0432
0473
0537
053F
04A7
045C
049C
04C6
047A
0427
044C
04CA
0530
0552
0531
04C1
0431
0406
047A
0500
04EC
046E
045B
04E2
0534
04BF
0435
0492
0553
0498
017A
FD7D
FB00
FAAF
FB35
FB3B
FAD0
FAB5
FB0D
FB4F
FB3A
FB26
FB53
FB82
FB73
FB5A
FB7F
FBBC
FBBC
FB8F
FB8B
FBAD
FB98
FB46
FB30
FB96
FBF0
FBA4
FB0A
FB0B
FBAF
FBD9
FAF3
FA55
FC08
002A
0455
0610
056D
0486
04CD
05A3
05C2
051D
04B2
04F8
054A
04FA
0443
03DA
03F8
0440
0466
0476
0480
046D
0456
0479
04CA
04D8
047C
042E
0456
0499
046F
042C
04A4
059D
0554
026D
FDFA
FAB8
FA15
FADB
FB17
FA81
FA32
FAA2
FB11
FAE5
FAA3
FB0F
FBF1
FC5F
FC0A
FB8E
FB6C
FB79
FB70
FB76
FBA2
FB9D
FB3D
FB0C
FB83
FC1F
FBF9
FB2B
FAD5
FB68
FBD1
FB20
FA68
FBE2
FFF0
0426
05F2
0569
04AA
04F8
059D
0586
04DE
0488
04B7
04D3
0488
0434
0431
044E
0459
0483
04E9
051D
04C7
044A
0448
04A1
04A7
0441
0427
04BE
054C
04FB
0446
0462
0536
04E1
01FB
FDAC
FA9B
FA0D
FAD2
FB2E
FAE3
FAD6
FB5B
FBC0
FB88
FB2E
FB5D
FBE4
FC0F
FBB5
FB55
FB46
FB51
FB38
FB26
FB54
FB91
FB8B
FB59
FB4E
FB5D
FB2A
FAD0
FAED
FB9B
FBEE
FB3E
FA96
FBF3
FFCF
041A
063D
05D6
04C0
0495
050C
050F
0485
043F
0488
04C6
0489
0433
044D
04A4
04AD
0462
0441
046E
0482
0454
0453
04C0
052A
051D
04DC
04E4
0506
04C3
045D
04AF
058F
053A
0241
FDB9
FA80
FA11
FB16
FB7D
FB03
FAD6
FB66
FBD4
FB7F
FB08
FB43
FBEA
FC0E
FB8F
FB3B
FB80
FBD5
FBB7
FB71
FB72
FB79
FB27
FACC
FAF7
FB68
FB5D
FAD4
FAAF
FB46
FB9D
FAE5
FA40
FBD3
FFE5
0408
05C2
053C
0487
04C4
053F
0516
049C
0497
04E9
04D9
044E
03F9
0434
0476
0443
03FC
043B
04D4
051F
04F8
04D2
04EA
04FB
04E3
04E3
0512
0502
047A
042F
04F4
061A
058E
022B
FD71
FA34
F9BD
FADA
FBA8
FB90
FB3C
FB39
FB5D
FB64
FB72
FBB8
FBF9
FBE3
FB91
FB5C
FB53
FB3A
FB08
FAFE
FB33
FB5D
FB46
FB28
FB51
FB92
FB73
FAFD
FAC1
FAED
FAF7
FA92
FAA9
FC98
0053
03F8
05AA
057B
0501
0533
057C
0505
0424
03DC
045E
04D3
0499
041C
041B
049E
0505
0504
04F5
0523
0557
053D
04EE
04BB
04B5
04BE
04D6
0500
0505
04BB
0470
0498
04E8
0438
01BC
FE31
FB54
FA27
FA2F
FA79
FABB
FB25
FB90
FB99
FB51
FB2F
FB59
FB6B
FB24
FAE6
FB26
FBA4
FBBB
FB4D
FAEE
FAF6
FB07
FAC6
FA80
FAAC
FB1D
FB57
FB5E
FB98
FBE1
FB85
FA89
FA68
FCB6
00FF
04CF
0622
0568
0496
04CC
0573
0592
051A
04B7
04C0
04E4
04C6
0484
047D
04CB
0521
0533
0507
04D8
04D3
04EF
04FD
04E4
04C0
04BB
04D1
04DC
04DC
04DE
0493
0342
0093
FD45
FAC8
F9F3
FA52
FAC6
FABD
FA83
FA8C
FAC9
FAE6
FAD5
FAD1
FAFA
FB31
FB5D
FB83
FB9A
FB83
FB32
FADA
FAB9
FAD0
FAED
FAFD
FB23
FB6B
FB85
FB13
FA66
FA93
FC92
001D
0399
0561
0544
0498
04B3
0584
05F0
0574
04CD
04E9
0599
05E5
0567
04C6
04B1
04EB
04C7
044B
0433
04CB
056D
0570
050E
04E8
04F9
04BA
043C
0458
055B
0601
047D
009D
FC65
FA2F
FA6F
FB9B
FC08
FB72
FAB2
FA7D
FAB8
FADF
FABA
FA87
FA9A
FAF1
FB4C
FB7C
FB86
FB7E
FB65
FB3A
FB14
FB0D
FB1E
FB2F
FB46
FB84
FBC7
FB95
FAC7
FA44
FB82
FEF2
0318
05AB
05C1
0485
03CA
042D
04E5
0527
0510
0525
0565
055F
04FB
04B1
04D0
0500
04CD
0462
0452
04BC
050B
04D8
048B
04C3
053D
050D
0408
0368
043D
0599
0513
018D
FCDD
FA13
FA4B
FBCA
FC51
FB8B
FAC6
FAD6
FB2F
FB10
FAC0
FAFA
FBAD
FBFD
FB81
FACE
FAAB
FB21
FB9B
FBB8
FB8F
FB49
FAEB
FA9E
FAD5
FBB8
FC9F
FC92
FB78
FA8C
FB68
FE83
028A
055B
05D6
04CA
0402
0465
0549
058E
050D
0492
04A3
04DB
04B5
046D
0493
04FD
04EB
044F
0415
04C5
058C
054F
0450
03D7
0451
04AC
040F
035B
03F5
0556
050B
01B5
FD13
FA45
FA62
FBAE
FC13
FB5F
FAC9
FAF6
FB5A
FB47
FAE9
FAD2
FB15
FB4A
FB42
FB3F
FB6B
FB8B
FB5A
FAFA
FAD6
FB1C
FB83
FBAB
FB9E
FBC3
FC36
FC68
FBCB
FAE8
FB58
FE27
0260
0598
063D
051B
043B
0490
053C
0529
0495
047D
0517
058A
053C
04AB
04A1
050D
0532
04CC
046E
0492
04DF
04C6
046A
0468
04C6
04C7
0418
038C
0411
051C
04C7
01E6
FDA1
FA81
F9DC
FABC
FB4F
FAFB
FA95
FAD8
FB64
FB73
FB07
FACF
FB17
FB5F
FB2B
FAC1
FAC1
FB2F
FB6F
FB3B
FB09
FB52
FBC8
FBC5
FB54
FB31
FBAF
FC1E
FBBD
FB10
FBB0
FE7E
0260
0527
05B4
04E8
046D
04EB
05A8
05BE
053A
04DC
0503
0549
0531
04DC
04C7
0507
052C
04F9
04BC
04C1
04CE
0482
040D
040E
0496
04E3
0469
03CC
0414
04EF
0490
01C3
FDAF
FAD9
FA7F
FB83
FC05
FB74
FAAA
FA6B
FA86
FA7C
FA60
FA97
FB0A
FB37
FAF5
FABC
FAF6
FB6D
FB8F
FB3E
FAF4
FB21
FB97
FBC9
FB98
FB7E
FBD2
FC24
FBC9
FB10
FB6B
FDFA
01FB
0525
05DC
04D1
0402
0469
0532
054D
04EB
04FE
05AC
0616
05AB
04F8
04CB
050E
050A
0499
0461
04C0
052A
0502
0494
0496
04E9
04B4
03C7
0337
0403
056B
054E
0273
FE10
FAB9
F9E9
FADA
FBC0
FBAC
FB16
FADC
FB22
FB57
FB10
FA95
FA73
FABB
FB01
FB0F
FB23
FB75
FBBA
FB88
FB04
FACE
FB23
FB7F
FB64
FB21
FB61
FBFA
FBFE
FB36
FB04
FD07
00FE
04B2
062B
0596
04AC
0491
04EB
04F0
04A6
04A7
050F
0551
0513
04B4
04B6
04FB
0500
04A3
045D
048E
04F1
04F9
04A3
046F
0499
04B4
045A
03FA
0459
0549
054F
0316
FF21
FB97
FA36
FAB7
FB75
FB5C
FACB
FAA5
FB11
FB75
FB6A
FB29
FB10
FB24
FB32
FB36
FB53
FB80
FB7F
FB3D
FAFF
FB0B
FB43
FB4D
FB26
FB37
FBBC
FC3C
FBF9
FAFF
FA9A
FC48
000E
040C
0615
05C4
04A1
044F
04E8
055F
0519
0494
047F
04C0
04C9
048B
047F
04C6
04E1
0486
0438
048A
0531
055A
04DD
0476
04AF
0510
04DA
0448
0452
0521
055C
038A
FFE5
FC4F
FA78
FA6F
FB0D
FB60
FB53
FB40
FB42
FB32
FB08
FAF8
FB26
FB6B
FB8B
FB80
FB75
FB79
FB6B
FB2F
FAF3
FB03
FB52
FB70
FB1D
FAC1
FAF1
FB85
FB9C
FAE0
FA73
FC00
FFB8
03B7
05BC
0562
0443
0406
04BD
0556
0538
04D2
04C0
04F1
04F2
04B5
049D
04D6
050C
04E5
0495
0497
04F8
0535
04EF
047E
0478
04DE
051F
04F6
04D9
0532
055C
0404
00BD
FCE7
FA89
FA55
FB2E
FBA7
FB73
FB30
FB3A
FB48
FB1A
FAEE
FB0F
FB49
FB3D
FAFE
FAFA
FB3F
FB50
FAED
FA91
FAD3
FB76
FBA7
FB20
FA99
FAD1
FB77
FB83
FAB1
FA36
FBA7
FF2D
0322
057E
05A6
04B4
0428
0477
04F6
04F5
04A0
049D
0511
0570
054D
04EE
04D6
0507
0515
04E4
04D9
052B
0570
052C
04A2
048A
0505
055C
051E
04D9
0531
0586
0447
00E3
FCDE
FA73
FA5C
FB5A
FBDB
FB8D
FB22
FB0D
FB18
FB07
FB03
FB31
FB4D
FB0B
FAA1
FA94
FAFE
FB5F
FB49
FAFE
FB0E
FB79
FB9E
FB24
FA8F
FAA2
FB3E
FB6F
FABE
FA34
FB81
FF05
0315
0576
0589
04AA
0473
0515
058E
0538
0491
046C
04D7
0527
04F8
04A8
04BD
0526
0564
053D
04F5
04D0
04B7
0489
0478
04C9
0542
054A
04BF
045A
04C5
056A
04A5
0195
FD68
FA76
F9F3
FAE9
FB8C
FB35
FAA4
FAA6
FB0D
FB33
FAFD
FAE4
FB1A
FB3F
FB0E
FAD9
FB03
FB5D
FB62
FB0D
FAE5
FB2E
FB72
FB33
FAB7
FAB5
FB3A
FB70
FADE
FA6A
FB9D
FED7
02A6
0519
0588
04E7
0489
04E2
0570
059F
056B
052C
0512
0500
04D4
04A2
0497
04BA
04E9
0507
0513
0508
04D6
0494
0498
0510
0595
057B
04C4
0456
04DE
0594
04B5
0179
FD47
FA87
FA3F
FB41
FBC3
FB43
FA93
FA74
FABF
FAF2
FAF8
FB17
FB5D
FB82
FB65
FB39
FB27
FB0E
FACE
FAAB
FAFD
FB91
FBB7
FB24
FA75
FA83
FB3D
FBA1
FB13
FA74
FB70
FE94
026A
04D6
0528
048A
046A
04F7
0565
0544
0506
0527
056B
0545
04C4
0481
04BF
0504
04E0
0496
04AA
0507
0513
04A6
045D
04B7
053F
0519
044E
03F8
04CB
05D1
0528
0214
FDF9
FB15
FA6F
FB25
FBB0
FB70
FAEC
FAC6
FAEE
FAEA
FAA9
FA96
FAEE
FB55
FB5A
FB1A
FB18
FB74
FBB3
FB71
FB04
FB06
FB6F
FB99
FB47
FB09
FB57
FBA9
FB29
FA3A
FA98
FD68
019A
04C7
05A5
051C
04CA
051C
0558
050F
04C6
0502
056D
0553
04BC
0469
04BF
0533
0514
0481
0433
047C
04E7
04EE
04AD
0498
04CB
04EB
04D1
04D7
0548
05A7
04E1
025D
FECD
FBBF
FA5E
FA92
FB41
FB68
FAE5
FA58
FA4D
FAB3
FB19
FB39
FB32
FB33
FB32
FB17
FAFF
FB1E
FB68
FB91
FB7D
FB67
FB7B
FB86
FB4C
FAFF
FAFC
FB23
FAE8
FA60
FAD3
FD7C
01BB
052F
0607
04E4
03EA
044A
0546
059D
0530
04D7
04FE
053A
0521
04F5
0513
0542
050F
048C
043E
045E
049A
049A
046C
044F
0459
048E
0504
0570
04DE
026F
FEA2
FB5C
FA28
FABA
FB86
FB8D
FB1E
FAEE
FB0B
FB0C
FAD6
FAB9
FADB
FAFE
FAF6
FAF3
FB25
FB65
FB7E
FB80
FB88
FB7C
FB51
FB55
FBC3
FC25
FBC3
FAE7
FB23
FDBA
01CF
04F5
05B5
04EC
0461
04AA
0503
04DF
04AE
04FD
0581
058D
0515
04AF
04B2
04D8
04D7
04CD
04D6
04BB
046C
044F
04A9
0500
04B5
041B
042F
04F3
04CA
0234
FDF3
FA9E
F9E0
FADA
FB9C
FB79
FB37
FB6D
FBA5
FB54
FACC
FABB
FB1C
FB46
FAF0
FA94
FAB0
FB23
FB85
FBB8
FBC3
FB8D
FB26
FAFF
FB58
FBA4
FB36
FA93
FB68
FEA3
02E0
0592
05B3
04A6
043E
04B1
0501
04C3
0491
04D8
0527
04F4
048B
049A
0525
0583
055A
0500
04CC
0497
0446
0436
04A4
0513
04F1
0491
04BC
052E
0458
013F
FD25
FA7E
FA48
FB34
FB90
FB36
FB0A
FB4C
FB5D
FAF6
FAAB
FAF5
FB6C
FB67
FB01
FADF
FB2C
FB6A
FB56
FB4B
FB86
FBA8
FB68
FB2E
FB5C
FB72
FAC7
FA12
FB2A
FECA
0326
05A3
05A6
04EA
04FF
0583
0554
048E
044F
04ED
0577
052C
0489
0471
04D7
04F2
0488
043B
0474
04D0
04D3
04AA
04AC
04B4
0490
04AB
0567
05ED
0493
00E4
FCB2
FA63
FA6C
FB27
FB16
FA7A
FA5C
FADB
FB3F
FB36
FB2D
FB67
FB92
FB68
FB37
FB5B
FB9B
FB85
FB3B
FB3D
FB7B
FB5F
FAE5
FADB
FB8C
FBF3
FB29
FA3B
FB6E
FF5B
03C1
05D9
0567
048E
04E2
05B9
05BB
04FB
049F
0506
055D
04FE
045A
042E
0478
04AC
049E
0497
04AD
04A6
0490
04C6
0532
052C
0496
045D
0523
05C2
0433
0020
FBCF
F9D5
FA60
FB6D
FB67
FAAC
FA5B
FAA0
FAD8
FAC9
FAD5
FB20
FB4D
FB30
FB1F
FB5A
FB93
FB77
FB46
FB6F
FBBC
FB93
FB0E
FAF8
FB74
FB7D
FA87
F9F4
FBE1
0050
04A0
0644
0572
0475
04BE
0593
05B7
053E
0513
0568
058E
0526
04AE
04AB
04F3
050A
04D7
0495
045E
042D
0432
0492
04E8
04A7
0423
0474
05BF
063B
03F0
FF46
FB0E
F994
FA5B
FB2A
FAD4
FA2A
FA47
FAFA
FB57
FB26
FAED
FAF7
FB09
FB01
FB21
FB7E
FBB8
FB87
FB3D
FB4D
FB8C
FB81
FB3F
FB57
FBB7
FB84
FA8A
FA49
FC83
00E5
04EE
0673
05C0
04CF
04D6
055D
057F
0534
04F6
04DF
04B8
0499
04CC
052C
0539
04D2
046A
0462
048B
0493
0499
04D8
0509
04BA
043F
047E
0560
053A
0297
FE4B
FAEB
FA14
FAE3
FB6A
FB00
FA89
FABD
FB30
FB37
FAFC
FB0F
FB6C
FB8B
FB43
FAFD
FB0A
FB43
FB6D
FB90
FBA8
FB73
FAEE
FAB7
FB4E
FC12
FBD0
FAA8
FA96
FD4D
01E2
0579
063D
051A
043F
049C
055E
058B
052C
04D5
04B7
04AD
04B9
04EC
050F
04DC
0486
0478
04B1
04BE
0481
0473
04D5
051F
04BC
0429
0475
0574
054B
0286
FE20
FABA
F9DD
FAA7
FB4A
FB1A
FABE
FACF
FB16
FB2E
FB24
FB27
FB1C
FAEC
FAD8
FB21
FB80
FB86
FB4C
FB4D
FB92
FB96
FB2A
FAED
FB59
FBBD
FB1A
F9FB
FA82
FDE9
02A1
05B9
05FB
04E6
0483
0521
059B
0546
04B5
04A2
04F7
052E
052C
052E
0538
051C
04E5
04C0
049E
0453
041B
0465
050C
0537
0489
03F2
0493
05CD
0565
021C
FD81
FA76
FA1F
FB16
FB7A
FAF6
FA76
FA82
FAC0
FAD4
FAE6
FB19
FB27
FAE2
FAB1
FAFD
FB80
FBAB
FB7C
FB68
FB80
FB53
FACC
FA97
FB1B
FB99
FB22
FA58
FB38
FEA1
02E0
0564
0585
04CF
04C9
0555
058A
0542
051A
0541
0539
04CA
047C
04BC
0524
0526
04DF
04C0
04BC
047C
043A
0493
056B
05B8
04F5
042C
04A4
05AE
04F6
0166
FCDC
FA34
FA28
FB0B
FB44
FAF0
FAED
FB3F
FB3C
FACF
FAA2
FAFB
FB49
FB19
FAD5
FB03
FB66
FB6D
FB33
FB3A
FB79
FB64
FAFD
FB07
FBBD
FC06
FAF4
F9AB
FAB1
FEDA
03CD
066E
061E
04D9
0479
04EB
0523
04E3
04BA
04EB
0516
0506
0508
053B
0536
04C9
0474
04AA
0506
04DF
0463
045A
04D0
04E2
0434
03D0
04AF
05CA
04C8
00ED
FC70
FA25
FA6D
FB56
FB4E
FAB9
FAAD
FB2E
FB61
FB08
FACA
FB15
FB6A
FB39
FAC8
FABD
FB23
FB70
FB60
FB2B
FB04
FAE5
FAE7
FB53
FBF9
FC06
FB23
FA7D
FBE9
FFAE
03CA
05E9
05B7
04C1
046B
04B5
04F7
0503
051A
0541
0537
0500
04E9
04F6
04CF
0472
0460
04D1
052D
04DC
0449
045A
050D
0560
04D9
0461
04DD
0560
03E2
FFF2
FBC6
F9E4
FA6C
FB66
FB65
FADC
FAD0
FB39
FB4A
FACF
FA6B
FA8E
FAE9
FB1B
FB42
FB87
FBA4
FB64
FB29
FB5D
FBA7
FB5C
FAB1
FAA2
FB6D
FBEC
FB36
FA6F
FBE2
FFFF
045E
0647
05A1
0484
0478
050C
0538
04F1
04E3
0535
0563
0535
050C
051A
0503
049A
0455
0493
04E9
04C6
0467
0476
04E5
04F2
0479
0468
053F
05AE
03C9
FF9F
FBA3
FA10
FA9F
FB6A
FB64
FB0D
FB01
FB04
FAB4
FA65
FA9F
FB31
FB71
FB44
FB39
FB7C
FB85
FB13
FAC5
FB25
FBAB
FB81
FAE8
FADF
FB83
FBAF
FAD7
FA71
FC7F
00CD
04BE
061E
0564
0492
04A8
0509
0508
04E3
0506
0539
0508
0499
0475
04A7
04B8
0489
0488
04E2
051A
04E1
04AF
04FB
054C
04E3
0424
044A
056D
05A9
0323
FE91
FAD2
F9D3
FAB2
FB59
FB13
FABF
FB00
FB5F
FB4A
FB09
FB30
FBA0
FBC0
FB77
FB42
FB54
FB4D
FB01
FAE0
FB2F
FB6F
FB22
FAC0
FB1E
FBF1
FBF3
FAE2
FA8A
FCE8
016F
0538
0626
050D
043A
04A1
054A
053A
04BF
04A5
04ED
0500
04B3
047A
0499
04C6
04C9
04D6
0510
0521
04CE
0477
048A
04B9
0472
03F6
043B
0541
0561
02FC
FEC4
FB55
FA65
FB17
FB7C
FB06
FAA6
FAFA
FB6E
FB49
FACB
FAAE
FB08
FB49
FB2F
FB12
FB2F
FB44
FB2A
FB31
FB7B
FB95
FB2D
FAD4
FB42
FC02
FBD6
FAB1
FA7D
FD0C
0190
051E
05E2
04EE
0474
050A
0587
051B
046A
0464
04E9
052A
04DE
0485
048E
04D2
0506
0525
0531
0509
04C1
04C1
051A
0536
04AD
0421
0482
0566
04FB
0215
FDF4
FB20
FAAF
FB5A
FB68
FABC
FA65
FAD3
FB63
FB80
FB65
FB78
FB94
FB5D
FAF9
FAE0
FB17
FB26
FAE1
FABB
FAFD
FB40
FB17
FAD6
FB0A
FB77
FB4E
FAB3
FB2A
FDF6
0231
055B
05F0
04E0
0432
04A3
0541
051A
047C
0454
04D1
0542
051E
04AF
048B
04C1
04E9
04D6
04D6
051F
0559
050C
0462
0429
04CC
057F
04BF
01E0
FDFD
FB1E
FA61
FB16
FBBB
FB8C
FB03
FAE1
FB36
FB77
FB5B
FB26
FB2D
FB4A
FB2A
FAE1
FADE
FB44
FBA5
FB91
FB33
FB18
FB56
FB53
FAB4
FA42
FB72
FEBF
02C7
0561
059F
048C
03E1
0442
04F5
0520
04CE
04A1
04DE
052F
0542
0539
054E
0553
04F2
0451
040A
0467
04E8
04E0
046D
0467
052B
05C3
04A5
0165
FD6A
FAC2
FA50
FB34
FBE6
FBBB
FB2F
FAF8
FB28
FB47
FB0D
FAB7
FA99
FAB6
FAE0
FB14
FB72
FBD9
FBE7
FB7C
FB14
FB3C
FBBC
FBB8
FAD6
FA1C
FB26
FE64
0268
0524
05C4
0528
04A7
04B3
04D5
04AC
047D
04B7
0540
0589
054D
04DE
04B3
04CD
04CD
048D
045D
0483
04BF
049E
043D
0453
052B
05CE
04AC
0151
FD37
FA92
FA42
FB2E
FBB1
FB4C
FACA
FAEA
FB77
FBB7
FB6F
FB0F
FAFC
FB14
FB09
FAED
FB11
FB69
FB87
FB38
FAEF
FB30
FBBF
FBC1
FAF4
FA70
FBC6
FF3A
032B
0582
05A5
04C5
045F
04BC
051B
04EE
047F
045D
048F
04B2
04A9
04BF
0516
0547
04F0
045F
0452
04F2
057D
0530
045B
0415
04C8
0552
040E
00B2
FCDA
FA8E
FA5A
FB1B
FB75
FB30
FAF9
FB33
FB7B
FB5D
FB0D
FB19
FB87
FBC4
FB7B
FB19
FB37
FBAB
FBB6
FB19
FA8E
FAD8
FB9F
FBC5
FAF9
FA80
FC03
FF9A
0374
0590
0591
04BF
047A
04E9
0549
0517
04AA
0496
04E3
0512
04D6
0476
0461
0493
04A7
0477
045D
04A2
04F5
04CB
044A
044C
0527
05C0
0462
00BB
FC94
FA3D
FA52
FB66
FBC8
FB38
FAAE
FAD8
FB62
FB9A
FB58
FB00
FAE4
FAF4
FB0E
FB37
FB76
FB99
FB73
FB36
FB50
FBD8
FC3A
FBCB
FABB
FA49
FBC7
FF39
0309
0551
058A
04D1
048D
04FB
054E
04F4
0461
045A
04E2
0542
0516
04C9
04D9
0514
04F2
0481
0460
04C0
04ED
044E
037B
03B6
0521
060D
048B
00A4
FC86
FA69
FA91
FB7D
FBC1
FB46
FADC
FAF8
FB4A
FB57
FB1D
FAF6
FB0E
FB3A
FB48
FB49
FB64
FB85
FB72
FB33
FB31
FBAA
FC2C
FBED
FAE9
FA5F
FBD3
FF67
0369
05BE
05C1
04A0
03F4
043D
04D6
0513
04F8
04E3
04EE
04E5
04C2
04C0
04F2
0502
04A8
0432
0438
04CC
0534
04D2
040F
03FB
04D6
0553
03C6
0016
FC2D
FA35
FA87
FB9D
FBE2
FB40
FAB6
FAD8
FB3C
FB41
FAF7
FAE3
FB26
FB52
FB22
FAEC
FB1F
FB8D
FB9D
FB30
FADC
FB22
FB9F
FB8B
FAF2
FB0E
FD0F
009E
03F4
057C
053E
0488
046C
04D9
0520
04FE
04D6
0500
0544
0530
04CD
049B
04E3
0548
0542
04D3
0484
04A6
04E3
04C9
048D
04C5
055E
0528
02FA
FF2C
FBA4
FA19
FA7F
FB57
FB6E
FAF5
FACD
FB2F
FB77
FB25
FA98
FA88
FAFF
FB52
FB0A
FA8C
FA8B
FB12
FB81
FB73
FB44
FB75
FBC4
FB73
FA89
FA60
FC6C
0074
0467
063E
05E4
04F1
04C4
0535
0551
04D7
0478
04BE
0544
0553
04EF
04C9
052F
0593
0557
04B5
0473
04C3
04FC
049E
042B
0486
057C
058A
0360
FF7F
FBE9
FA3E
FA5C
FAEF
FB01
FABA
FABA
FB14
FB4C
FB1B
FAD4
FAEA
FB3F
FB4B
FADB
FA6F
FA9B
FB41
FBA9
FB70
FB04
FAFD
FB37
FB0A
FA84
FADC
FD39
0119
0471
05A4
0515
0472
04BA
055D
0563
04D4
048A
04E7
0557
0534
04B9
04A2
0517
0572
0527
048B
0459
04B8
0514
0507
04EC
0549
05C5
052E
02AD
FEE6
FB9A
FA25
FA6B
FB38
FB8A
FB4C
FAFD
FAE9
FAF0
FAEC
FAF6
FB28
FB54
FB39
FAF7
FAFC
FB68
FBBD
FB7A
FADF
FABA
FB54
FBDE
FB66
FA4C
FA47
FCAC
00CC
046A
05DC
0576
04C6
04C3
0514
0508
04AD
04A4
051A
0579
0534
0491
044C
0497
04E9
04CB
0484
04A0
0505
0504
045F
03DF
0460
0576
0574
0320
FF30
FBC1
FA58
FAA9
FB4D
FB5C
FB10
FB05
FB49
FB68
FB21
FAC9
FACD
FB23
FB60
FB4A
FB1C
FB28
FB5E
FB6C
FB45
FB4A
FBAD
FBF8
FB8D
FABC
FAF1
FD53
0141
0496
05AB
04E5
040A
0435
04E6
0517
04AF
046C
04B7
051D
051C
04E9
0510
0582
0594
04FB
044C
0438
049A
04B5
0453
041D
04A0
0545
04A8
0218
FE7D
FBA5
FAA3
FB0C
FBA8
FBB5
FB63
FB39
FB5B
FB71
FB41
FB03
FB07
FB2F
FB14
FAAA
FA74
FAD6
FB7A
FBB2
FB68
FB3D
FB9B
FBF7
FB84
FA99
FAD5
FD6B
018D
04EA
05E2
04F2
03E6
03EF
04B2
052A
04F3
048D
0488
04D8
050D
04FA
04DF
04F2
050F
04F8
04BD
04AA
04CA
04BD
0456
0415
0497
0571
051E
027E
FE5A
FAF1
F9E2
FAC0
FBD2
FBFD
FB8B
FB43
FB48
FB3B
FB01
FAEE
FB27
FB52
FB22
FAD8
FAF8
FB7D
FBC8
FB76
FAF7
FB0C
FBB7
FC10
FB70
FA8C
FB0C
FDD0
01D0
04E4
05C3
0511
0467
048D
04FC
04F7
049D
0490
04F5
0534
04E8
0473
0479
04E6
050A
049D
042D
0456
04D2
04DA
0457
0422
04D6
05AB
04F7
01F6
FDD9
FACB
F9F9
FAAD
FB52
FB23
FA9F
FA93
FB0F
FB73
FB5C
FB20
FB36
FB88
FB96
FB4C
FB2A
FB84
FBEF
FBD1
FB4B
FB1B
FB7A
FBA1
FAE0
F9FB
FAC4
FE15
0290
05C1
0675
058E
04B8
04B4
0511
0534
0519
0511
0520
04FC
0496
0449
045F
04A9
04B4
0460
0415
0437
049C
04BB
047C
0477
0525
05D7
0507
01F6
FDC2
FA92
F99C
FA39
FAF3
FB16
FAFA
FB0E
FB26
FAF6
FAB6
FAE5
FB78
FBCF
FB86
FB03
FAFA
FB82
FBF9
FBE0
FB7E
FB73
FBCC
FBDB
FB2C
FA6F
FB19
FDE9
01EC
051F
0635
05A4
04EB
04ED
0552
055A
04F5
04AE
04CF
0506
04F7
04CA
04D9
0509
04DE
0446
03E0
0432
04D7
04F4
0469
041A
04BE
0595
04E7
01DE
FDAE
FA99
F9D1
FA8C
FB30
FB0D
FAB1
FACD
FB3E
FB60
FB0E
FACD
FB00
FB56
FB50
FB0D
FB2B
FBC9
FC30
FBC0
FAE6
FAAA
FB43
FBB7
FB2D
FA64
FB2E
FE66
02B2
05B8
0661
0598
04F1
04F7
0517
04CF
0475
049F
0538
058B
0536
04A9
0486
04CA
04E1
0491
044E
0488
04F5
04EE
0474
0458
050D
05AC
049A
0155
FD47
FA84
F9E3
FA84
FB0C
FB00
FAD3
FAF9
FB50
FB63
FB18
FACA
FAD0
FB14
FB40
FB30
FB1C
FB3A
FB65
FB4E
FB06
FB02
FB6E
FBB4
FB3F
FAB2
FBAD
FEF9
0329
05C3
05C5
0495
0434
04F8
05A5
055C
04AD
0485
04DC
050B
04EE
04F4
0538
0542
04E2
04A5
04F7
054F
04E2
0403
03E3
04B0
04C7
028C
FE9E
FB6B
FA82
FB13
FB5A
FAD0
FA5C
FAA7
FB37
FB54
FB1C
FB27
FB7C
FB8A
FB22
FABF
FACC
FB09
FB18
FB22
FB7E
FBDE
FB87
FA9E
FA9E
FCE4
00DF
0453
058F
050C
0484
04DF
0580
0581
04F8
04A2
04C4
04EC
04C6
049B
04C8
0511
04FF
04A3
048C
04DA
04FF
04A1
044E
04B6
0546
045C
0133
FD2B
FA8E
FA33
FAE3
FB1D
FAC6
FAB6
FB2C
FB7B
FB34
FAD4
FAFB
FB69
FB74
FB1C
FB0F
FB87
FBD2
FB68
FADA
FB09
FBB3
FBB2
FADF
FADF
FD55
0198
050D
05F1
051C
0499
0520
05A8
0547
0481
0463
04F9
055C
050E
048F
047C
04B8
04D0
04C4
04DB
04F4
04A3
041B
0437
0522
0577
038B
FF95
FBDF
FA6C
FAE7
FB6D
FAFF
FA60
FA93
FB4C
FB80
FAFB
FA9A
FAEF
FB7A
FB7F
FB24
FB11
FB5A
FB6C
FB25
FB1D
FB9D
FBE3
FB32
FA67
FB76
FF0C
034E
05A1
0570
047A
047B
054F
05BC
055A
04F1
0511
0546
04F2
045E
044A
04C7
0522
04F5
04AA
04AA
04AC
0449
03F1
0471
056F
0534
0285
FE63
FB3F
FA75
FB21
FB8C
FB29
FAB0
FAB2
FADA
FAB4
FA83
FACC
FB72
FBCA
FB8D
FB2D
FB16
FB21
FB03
FAF2
FB59
FBF8
FBF8
FB31
FAE1
FC8D
0025
03C0
0578
053C
0488
0490
0529
057B
0544
04FD
04FC
04FE
04B8
0465
047A
04E7
052F
0518
04EF
04F0
04DC
047E
0446
04B9
0547
0457
011B
FCFC
FA72
FA6C
FB71
FB9C
FAC6
FA39
FAA6
FB4F
FB52
FAEB
FAE6
FB47
FB5D
FAFA
FAC8
FB27
FB81
FB44
FAE7
FB32
FBD0
FB9A
FA90
FA8D
FD3B
01B3
0520
05D1
04DE
0463
04F1
0577
0535
04BE
04D2
053A
0542
04EB
04D7
0533
0561
04F7
0471
0473
04C2
04B1
045B
04A2
05A6
05F2
03DB
FFAB
FBB5
FA0D
FA90
FB74
FB7A
FAF7
FACB
FB0E
FB2B
FAF2
FACF
FB03
FB37
FB12
FAD4
FAED
FB3D
FB3E
FAEC
FAEA
FB74
FBB8
FAFE
FA2C
FB43
FEF1
0353
05C3
059F
049D
0478
0513
0548
04CA
0472
04CE
0552
054D
04EB
04CA
04F6
04FB
04CD
04E0
0542
0546
0493
03FB
0481
05A1
055F
027D
FE29
FAEE
FA1B
FAC7
FB54
FB31
FAEB
FAFB
FB2D
FB27
FB04
FB12
FB45
FB47
FB02
FAC8
FAD3
FAF4
FAF0
FAF0
FB3E
FBAD
FBA0
FAF8
FAB9
FC4B
FFD5
03B4
05E2
05E5
0502
04A1
04EB
052D
050B
04D9
04E4
04F4
04CA
04A0
04CF
0524
0523
04D1
04BA
0501
050A
0482
0421
04AE
056F
047D
0116
FCEE
FA91
FA9B
FB64
FB4B
FA8F
FA61
FAFB
FB77
FB4C
FAFF
FB20
FB5E
FB25
FAAC
FAAF
FB37
FB78
FB12
FABE
FB2C
FBC9
FB7A
FA8E
FAEB
FDD2
020A
04FA
0572
04B0
048A
0541
05BE
0567
04E0
04E4
052D
0505
047F
045E
04E0
0559
0531
04C5
04CA
0523
0511
0482
045F
0516
0567
038C
FF94
FBC1
FA31
FAB2
FB6A
FB3A
FAB1
FAAB
FAF9
FAE0
FA6E
FA6D
FB16
FBA3
FB71
FAEE
FAE3
FB3E
FB4B
FAF0
FAE3
FB70
FBBF
FB11
FA4D
FB67
FEFE
0343
05BA
05C5
04DD
048A
04E2
0524
0514
0519
0559
0568
0507
049D
04A6
04F6
0503
04C7
04C5
0523
054D
04D7
0451
0498
0556
04E2
0217
FDF0
FAC8
F9FF
FAC8
FB76
FB5D
FB12
FB21
FB45
FB18
FAD4
FAF4
FB5B
FB70
FB0A
FAB5
FAE0
FB2E
FB16
FAC7
FAEF
FB85
FBAB
FB0E
FAE5
FCCD
00A3
0445
05B7
0527
0460
048C
052F
054C
04DD
04A2
04E3
0521
04F0
04A2
04BA
051E
0548
050F
04CF
04C0
04A1
044E
043B
04CD
054D
0438
00FD
FD0B
FA9F
FA84
FB75
FBC2
FB27
FA99
FABF
FB30
FB44
FB0D
FB0A
FB43
FB48
FAF8
FAC4
FAF9
FB3F
FB33
FB18
FB68
FBDE
FBA5
FACE
FAEA
FD6B
01A2
050E
05F6
051A
0470
04C0
0535
0500
048D
04A2
0515
0519
0491
044B
04C5
0562
0555
04D0
049E
04DA
04D5
0459
0438
04F4
0565
03B2
FFBB
FBC0
FA16
FAAE
FB8A
FB55
FAAE
FAC0
FB6F
FBAD
FB29
FABE
FB1C
FBBB
FBAC
FAFD
FA91
FAD4
FB3F
FB51
FB4B
FB8F
FBB5
FB29
FA8F
FB93
FEEC
0306
0575
057C
0493
045E
04EB
0535
04DF
048C
04B7
04FA
04D7
0490
04AE
0510
0518
04B7
048F
04EB
0528
04AF
040E
0453
0548
0526
028F
FE70
FB3E
FA68
FB1A
FBA2
FB64
FB05
FB17
FB52
FB3B
FAF6
FAFC
FB4D
FB77
FB50
FB34
FB5C
FB71
FB1E
FABC
FAEF
FB94
FBB7
FAFD
FA9A
FC43
000C
03EA
05B6
0554
0474
046A
04EC
050E
04BB
04A3
0504
0542
04E3
0455
044F
04C2
0509
04EA
04DA
0513
051C
04A5
044F
04D1
0582
0490
012B
FCEC
FA5D
FA55
FB5B
FBAF
FB30
FADE
FB22
FB66
FB3D
FB0C
FB4D
FBAB
FB84
FAEF
FAAA
FAFF
FB59
FB39
FB05
FB54
FBC8
FB73
FA83
FAAF
FD62
01B5
0511
05DD
0500
0470
04DE
0563
052E
04A3
0488
04D0
04CE
0469
0445
04B8
0533
051C
04B6
04A7
04E5
04CE
045F
0477
055F
05BA
03BF
FF9E
FBBC
FA35
FAB3
FB4D
FB03
FA8E
FACF
FB65
FB6E
FAFB
FAED
FB83
FBEA
FB81
FAD7
FACF
FB48
FB64
FAF9
FAD5
FB61
FBBF
FB14
FA3F
FB49
FEE6
0337
05A9
05A5
04CF
04BA
0541
0562
04EF
04A4
04DE
050E
04B1
0437
0457
04F5
053E
04E7
0494
04CB
0516
04C6
0437
046A
054F
0533
029E
FE62
FB09
FA2D
FAF3
FB73
FB07
FA8E
FAC7
FB47
FB52
FB01
FAFD
FB63
FB9F
FB5F
FB0C
FB15
FB43
FB2E
FB05
FB49
FBCD
FBB5
FADA
FA92
FC76
0058
0419
05C7
056F
04A5
0490
04F5
0511
04CB
04A5
04D6
050A
04F4
04C2
04C2
04E0
04DB
04BD
04CB
04FC
04EE
0486
0458
04D9
0556
0441
00F5
FCE0
FA5E
FA58
FB81
FC00
FB6E
FACB
FAE0
FB4D
FB5A
FB0D
FAF8
FB3B
FB63
FB38
FB1D
FB53
FB79
FB2C
FACA
FAF7
FB81
FB89
FB04
FB63
FDFB
0206
0511
0597
0495
040C
0497
052C
04F6
0479
048E
0509
0517
049E
0464
04CF
0539
04FA
0480
04A3
0541
0552
048F
0411
04AB
0539
03A8
FFAE
FB9E
F9F0
FA97
FB82
FB57
FAC1
FAE5
FB95
FBC7
FB53
FB17
FB7E
FBCA
FB50
FA98
FA8A
FB06
FB2B
FAD8
FAE0
FB8C
FBD9
FB05
FA4A
FBD2
FFD7
03E6
0596
0515
0461
0494
050E
0501
04B0
04B2
04E4
04C0
0464
046A
04DE
0524
0510
052E
059A
0591
04B6
0410
0499
0557
0419
0052
FC2D
FA35
FA8A
FB44
FB2B
FADD
FB2B
FBA4
FB7C
FAF6
FAE4
FB45
FB68
FB25
FB07
FB3A
FB3C
FAD1
FA9B
FB11
FB81
FB17
FAA7
FC26
FFF7
03EC
05B3
056D
04F1
052C
056A
0501
046F
046E
04CF
04EC
04BD
04C2
04FC
04EF
04A9
04D3
056B
057D
04BA
0449
04F9
0570
0382
FF3F
FB57
FA1D
FAFF
FBB4
FB3B
FA9A
FACC
FB5B
FB76
FB44
FB53
FB7A
FB47
FAF8
FB19
FB71
FB50
FAC9
FAB0
FB35
FB64
FAC6
FABE
FD21
017C
0512
05EF
0503
0476
04E8
0559
0522
04BA
04A1
04AA
048D
0480
04B9
04E7
04B5
0483
04D6
054B
050D
045F
0481
0581
055A
0263
FDD4
FAAB
FA44
FB37
FB96
FB27
FAE1
FB13
FB26
FAEC
FB01
FB8C
FBCA
FB51
FADE
FB24
FB9E
FB7A
FB06
FB1E
FB93
FB5E
FA95
FB10
FE2C
029C
0587
05BA
04BB
0472
04F1
0530
04EC
04C2
04E9
04FD
04DC
04CF
04E6
04CB
0476
0465
04C4
04F0
0479
041F
04D4
05C9
04C2
00F9
FC95
FA58
FA92
FB5F
FB5D
FAF2
FAF0
FB35
FB2B
FAEB
FB01
FB56
FB4B
FADB
FAC4
FB41
FB9B
FB64
FB43
FBB1
FBE7
FB16
FA46
FBA1
FF99
03EB
05F7
0590
04A6
0498
04FD
0502
04D3
04EC
0515
04E3
04A0
04D6
0540
052F
04B3
0487
04CF
04CC
0436
0403
04EE
05B1
040D
FFCD
FB93
F9EF
FA9D
FB75
FB55
FAE6
FAED
FB26
FB10
FADF
FB03
FB4F
FB3F
FAEC
FAEB
FB43
FB60
FB32
FB63
FC02
FC01
FAED
FA5D
FC63
00C6
04CF
063B
057A
0496
049B
04F0
04EF
04E2
0523
054B
04F0
0483
049A
04F5
04F2
04AA
04AF
04F6
04D9
0454
044A
0507
0520
02D8
FE97
FAEB
F9C1
FA75
FB30
FB38
FB1D
FB3E
FB4A
FB15
FAFC
FB32
FB5C
FB32
FB04
FB32
FB6F
FB3B
FADD
FB10
FB9F
FB7A
FAA7
FAFC
FDFA
0277
059C
0610
051D
04A7
04F8
051F
04C8
0497
04DF
0507
04A9
044B
047C
04E9
04FC
04D7
04EA
0506
04BB
0462
04C8
058F
04E4
0197
FD0B
FA10
F9DC
FAF9
FB7C
FB2D
FAF4
FB18
FB1C
FAE8
FAF6
FB5F
FB98
FB56
FB05
FB16
FB43
FB1E
FAF2
FB46
FBB8
FB5F
FA96
FB4A
FEA4
031A
05E5
0607
04FC
0489
04D5
0504
04CF
04BB
0507
053B
0503
04B2
04AB
04D1
04E8
0507
0527
04E4
043E
0407
04C8
0579
043C
00A2
FC8D
FA4C
FA46
FB03
FB45
FB29
FB39
FB52
FB24
FAED
FB05
FB2F
FB07
FAC9
FAF4
FB5A
FB56
FAEE
FAEF
FB9A
FBF1
FB34
FA92
FC27
0025
041B
05BB
0556
04D4
0505
052F
04CD
0476
04BD
0531
0521
04C1
04C8
052A
0526
04A3
0469
04BF
04DE
045E
042B
04FB
0587
03B3
FF77
FB6B
F9F3
FAAF
FB73
FB24
FA97
FAB9
FB2A
FB2E
FAF7
FB17
FB66
FB5A
FB0A
FAFF
FB3B
FB3F
FB08
FB25
FBA0
FBA0
FAD6
FAAD
FCF7
0157
0519
062A
053E
0478
04B5
052D
0530
0504
0513
052B
04FB
04B9
04BF
04E7
04D5
04AA
04CE
0511
04D8
0454
047E
055E
0537
0281
FE26
FACC
F9F2
FAA5
FB2E
FB16
FAFB
FB1E
FB19
FAD9
FADF
FB46
FB66
FAF2
FA99
FAE8
FB57
FB31
FADA
FB28
FBCC
FB9B
FAA5
FAE5
FDEC
027C
0593
05D5
04D1
0493
052E
0570
0505
04AC
04C6
04E2
04B5
04A3
04F5
0551
0551
0529
0535
0530
04AF
0430
0497
0563
0496
012C
FCDA
FA51
FA46
FB25
FB65
FB11
FAE8
FB05
FB05
FAF2
FB2D
FB86
FB63
FADA
FAB6
FB27
FB5A
FAE8
FAA9
FB42
FBCF
FB33
FA4F
FB78
FF62
03C8
05D9
056A
049D
04D3
054F
0515
049C
04BE
0529
04FF
0472
0471
050D
055A
04F3
0496
04D2
050D
04A0
0439
04D9
05A4
0446
0021
FBC0
FA08
FADD
FBCE
FB72
FAAD
FAB6
FB44
FB5B
FAF6
FAE0
FB45
FB77
FB27
FAE5
FB13
FB3A
FB0A
FB08
FB85
FBBB
FB08
FA8D
FC46
005A
0463
05F7
053D
044D
0471
0508
0517
04C8
04C6
0506
050E
04E6
04E7
04FD
04DD
04AF
04D6
0520
04F2
0464
0467
053D
056E
0337
FF08
FB6F
FA48
FAD6
FB49
FB15
FAF8
FB46
FB78
FB3D
FB02
FB1F
FB3D
FB04
FACE
FB18
FB8C
FB70
FAEB
FAE4
FB6A
FB68
FA96
FA9E
FD33
0187
04E1
05B2
050D
04C9
0535
0552
04C2
044D
047D
04D2
04C0
049C
04DC
0528
04F4
0482
047A
04C8
04D2
04A1
04EB
0594
0512
0225
FDD7
FAC0
FA2E
FAEF
FB36
FACE
FAA7
FB10
FB6A
FB5B
FB42
FB6A
FB8C
FB5D
FB18
FB1E
FB52
FB5E
FB55
FB7D
FB87
FAEB
FA39
FB24
FE7A
02B4
0567
05C9
051F
04D3
04FC
04FC
04BC
04AE
04E0
04E1
048D
0454
047A
04B0
04B5
04C2
04F6
04EB
0479
0453
050A
05B1
0472
00D5
FCB5
FA64
FA47
FAE0
FAFE
FAEC
FB42
FBAD
FB87
FB04
FAE3
FB45
FB97
FB8A
FB67
FB68
FB5D
FB2F
FB38
FB97
FBA4
FAEA
FA69
FBF2
FFC5
03C4
05B0
0588
0507
0533
0577
0510
045C
043B
04C4
0536
0516
04B2
047C
0478
0486
04A7
04B5
0465
03F8
043E
0548
059C
0390
FF79
FBB1
FA2F
FA9B
FB26
FADF
FA70
FAAF
FB5A
FBAD
FB75
FB17
FAE0
FAE0
FB26
FB8E
FBAC
FB5E
FB34
FBB8
FC68
FC1F
FAE0
FA83
FCD0
011C
04AD
05B8
0511
049D
04F6
055C
0548
0505
04E6
04CD
04A9
04B9
0509
0524
04BC
044D
046E
04BE
046A
03B1
03D2
04F0
051E
0294
FE39
FAE3
FA2B
FAFE
FB73
FB18
FAC8
FAF5
FB20
FAF5
FAE3
FB3B
FB8B
FB67
FB29
FB46
FB80
FB68
FB47
FB9D
FC08
FBAB
FAD3
FB43
FE2B
0251
0526
059B
0500
04E6
0549
0554
0503
04F6
053B
053A
04C3
045C
0460
048B
0493
04A2
04D7
04C5
042D
03D5
049A
05A6
04C2
011E
FCC8
FA7B
FA92
FB33
FB03
FA84
FAA6
FB2E
FB43
FADE
FAC2
FB2B
FB81
FB75
FB79
FBB9
FBA4
FB07
FAC5
FB80
FC45
FBCA
FABC
FB78
FF0F
0383
05E1
0596
04A5
04C0
056D
0571
04E0
04AD
050B
0544
0502
04B3
04A3
0490
044E
0434
0483
04D7
04BB
0483
04BB
04D6
0366
000A
FC6E
FA91
FA9D
FB29
FB2E
FAE3
FAD4
FAF8
FAFB
FAE2
FAEA
FB0A
FB0D
FB0E
FB58
FBC0
FBD0
FB8F
FB8E
FBCF
FB8C
FAA3
FA83
FCBD
00D1
0461
05B4
0557
04EC
0512
052F
04EF
04D3
0527
055D
04FB
0480
0498
0500
04FA
048D
0468
04A6
048E
03E6
03AD
049D
057A
0407
FFE1
FB76
F96E
F9E4
FADB
FAF3
FA9D
FAB4
FB18
FB26
FAE8
FAF9
FB76
FBC0
FB75
FB0E
FB1E
FB77
FB8E
FB6C
FB94
FBF3
FBC9
FAE1
FA6F
FC0C
FFC9
03C4
05E8
05E0
0515
04E3
054F
058E
054B
04F0
04DB
04DD
04AB
0470
048A
04E3
04F9
04A6
0463
0497
04E4
04BF
0468
049E
0528
047D
0180
FD45
FA49
F9D7
FACD
FB45
FAD3
FA84
FAFC
FB94
FB83
FB10
FAFD
FB50
FB6E
FB36
FB2E
FB8C
FBBF
FB5B
FAEA
FB28
FBBA
FB87
FA96
FAA5
FD3A
0189
0504
0610
0570
04E3
050B
0536
04D7
0461
0480
050C
0548
04F2
0485
0476
04A0
04AA
049B
04B3
04DE
04CB
048F
04BB
0571
05A6
03E9
001F
FC1A
F9FB
FA21
FB16
FB6A
FB1A
FAFC
FB50
FB88
FB4D
FB0B
FB37
FB87
FB69
FAFE
FAF1
FB5F
FB97
FB34
FAD3
FB1F
FBA0
FB56
FA8B
FB0E
FE1F
0286
0591
05EF
04D6
043D
049E
0510
04EE
0498
0491
04BD
04C3
04B6
04DE
0513
04F0
048F
0489
0503
0545
04B9
0402
0447
0566
058B
0326
FEEB
FB61
FA51
FB22
FBDE
FB88
FAD4
FACD
FB66
FBBF
FB75
FB08
FB05
FB4A
FB5E
FB37
FB2A
FB4F
FB5E
FB45
FB56
FBA7
FBA2
FAE4
FA63
FBD2
FF88
0391
0589
0525
043F
0467
0535
0555
049C
0424
048D
051F
0501
0484
0482
04F9
051A
04A1
043F
047A
04CE
049A
044A
04C4
059F
0507
01E5
FDA0
FAD5
FA8F
FB7C
FBD1
FB47
FACD
FAEF
FB48
FB59
FB40
FB43
FB40
FB02
FAD3
FB25
FBC3
FBEE
FB6B
FAF4
FB34
FBB5
FB71
FA7E
FA7B
FCD8
00F7
0483
05C1
0522
045A
0467
04DD
04FE
04C6
04AE
04DA
0500
04FA
04FA
0518
0506
0498
043A
0465
04D9
04DB
0468
046D
0561
060F
048B
0093
FC44
FA16
FA61
FB6D
FBB0
FB4B
FB25
FB67
FB73
FB09
FAAA
FABE
FAFA
FAF2
FAD2
FB0B
FB82
FB9A
FB32
FAEA
FB2B
FB63
FAD9
FA21
FAF1
FE28
0275
056A
05E4
04E9
0437
0472
04F1
0505
04CE
04CA
050D
0545
0542
0522
0502
04D4
04A1
049D
04D9
0503
04D6
04A0
04F4
059B
0544
02CA
FEC8
FB65
FA4A
FB0A
FBDB
FBA5
FAE9
FAA7
FB01
FB4C
FB2A
FAEB
FAE4
FAF1
FAE2
FAEB
FB43
FB9B
FB75
FAFA
FAE4
FB5F
FB9B
FB05
FA96
FC0F
FFB8
039A
056F
050E
043E
0464
0522
055E
04F4
04AC
04E2
0511
04CB
0479
04A5
0510
050B
0498
046E
04CD
0507
0491
0414
048C
057C
04F3
01C9
FD66
FA86
FA61
FB9A
FC29
FB91
FAD7
FACA
FB19
FB2E
FB1B
FB49
FBA4
FBB4
FB69
FB32
FB46
FB4D
FB09
FAEA
FB60
FBED
FB93
FA77
FA57
FCC3
0113
04C4
05FE
0544
046B
046B
04C3
04C5
0497
04B4
04FF
04F1
0480
043E
0478
04C1
04A9
046D
048E
04E9
04E1
0477
0482
0563
05E4
043E
004F
FC33
FA2C
FA69
FB3F
FB5F
FB0F
FB2A
FBA6
FBC4
FB55
FB0C
FB5F
FBCA
FB9F
FB23
FB29
FBC7
FC1A
FB96
FADC
FACA
FB20
FAF1
FA64
FB14
FE29
0279
0570
05CD
04C6
0445
04B3
0511
04C4
045A
0476
04C9
04AC
043C
042E
04A7
04F2
04A1
0439
0461
04CF
04C9
0473
04B9
05AC
05AE
032A
FECC
FB34
FA3A
FB21
FBDC
FB90
FB0A
FB1E
FB75
FB66
FB1E
FB4A
FBE0
FC13
FB94
FB15
FB37
FB8C
FB52
FAC5
FAE0
FBB7
FC0F
FB27
FA51
FBC1
FFB6
03D2
05A0
0529
0461
0484
04FA
04D4
045E
047D
051A
0533
0467
03A3
03CB
047E
04C2
0485
0495
052F
057C
04DF
0424
046E
0549
04B9
019A
FD56
FA8D
FA4C
FB49
FBC0
FB5A
FAF3
FB0D
FB4B
FB43
FB2E
FB6D
FBDC
FC03
FBD2
FBA7
FBA0
FB6B
FAE8
FA98
FAF4
FB98
FB9E
FAFD
FB0E
FD2A
00F3
0465
05CC
055F
04A5
04A3
0513
053E
050A
04D8
04CA
04A1
0451
0433
0473
04AF
0486
043F
046C
04F5
051E
04AE
046B
04F1
055B
03EC
0048
FC55
FA60
FAAF
FB85
FB6F
FAC2
FA93
FB03
FB47
FB0E
FAF0
FB5B
FBC8
FB8E
FB04
FB13
FBC9
FC2F
FBAE
FB01
FB12
FB88
FB4D
FA84
FAF5
FDEE
0246
0551
05BF
04D0
0473
04FF
0557
04DF
0455
048B
0527
053A
04A9
0441
047B
04D6
04BF
0471
047C
04C2
04AF
0456
048C
0575
0597
0351
FF13
FB5B
FA21
FADD
FB90
FB46
FACD
FB0C
FBA8
FBBA
FB3F
FB0A
FB69
FBBD
FB8A
FB37
FB4E
FB86
FB46
FAC7
FAE7
FBAF
FBF5
FB0C
FA3A
FB9A
FF78
039F
05AC
0579
04B0
0484
04AE
0492
045F
0495
04FC
04E4
044B
03FE
0468
04E8
04C5
0450
0467
050C
0542
0495
03F4
046E
0564
04D6
01C7
FDA6
FAF1
FAA1
FB7F
FBE7
FB89
FB2C
FB46
FB7F
FB77
FB5D
FB82
FBBF
FBB2
FB6E
FB67
FBAD
FBB8
FB3D
FAD0
FB1F
FBD6
FBE2
FB21
FB11
FD3E
0129
0478
0569
0497
03EB
044A
04E9
04DC
0463
0454
04BE
04ED
0487
040B
03FF
043A
044E
0454
04A6
0510
04EE
0446
040E
04C6
0547
03BE
FFFB
FC14
FA49
FABA
FBA4
FBA9
FB21
FB10
FB90
FBDB
FB95
FB41
FB61
FBBA
FBCE
FBAD
FBBE
FBEC
FBB2
FB09
FABC
FB49
FBF5
FBAF
FAD4
FB48
FE44
0290
058B
05F4
04F9
0473
04C8
050A
04B2
044D
046D
04BD
049C
0435
0435
04A7
04CF
045F
040A
0472
0515
0504
046F
047C
055C
0562
02DA
FE79
FAF4
FA14
FAEF
FB73
FAFC
FA96
FB05
FBAB
FBA4
FB1E
FAF7
FB57
FB90
FB4E
FB23
FB89
FC04
FBD4
FB2F
FAF5
FB49
FB40
FA73
FA2C
FC28
0047
043A
05DD
0563
04AA
04D7
0556
0530
048D
0451
04B7
050C
04CC
045E
0462
04BF
04E0
04A9
0495
04D1
04DE
047B
0454
051F
060F
0522
0176
FCC4
F9E4
F9E0
FB22
FB92
FAEC
FA6C
FACA
FB5D
FB55
FAF0
FAF5
FB7A
FBDC
FBCB
FBA7
FBB8
FBA8
FB2F
FAC7
FB16
FBBD
FBA1
FAAA
FA88
FCF0
015A
052B
0667
0592
04B0
04D7
0563
0561
04E5
04AF
04EB
050F
04BF
0453
0440
0469
046B
043C
0432
0467
0497
04AA
04ED
0566
0539
034D
FFBC
FC32
FA66
FA72
FAFB
FAE9
FA7B
FA80
FB08
FB5D
FB20
FACB
FAF0
FB64
FB96
FB79
FB7C
FBC0
FBD3
FB75
FB1C
FB3C
FB76
FB28
FAC9
FBDE
FF20
031F
0583
0594
04D1
04DF
059B
05CB
051A
0483
04C2
0550
0549
04CB
04A7
0500
050F
0472
03EB
0440
04F8
04F6
0435
03F1
04BC
052E
034D
FF1E
FB02
F944
F9DA
FAE9
FB16
FAAB
FA8C
FADD
FB12
FAED
FAC6
FAEB
FB2C
FB3A
FB2B
FB45
FB78
FB6D
FB1F
FB08
FB7C
FC0C
FBE8
FAF5
FA43
FB39
FE34
0213
0519
0640
05D8
04FC
049B
04D7
053B
0553
051D
04E7
04E9
050A
050D
04E2
04AC
0495
049A
049F
049B
049D
04B1
04DB
051F
0574
0583
049B
0232
FEA2
FB48
F994
F9CF
FAE3
FB77
FB2C
FAB8
FACA
FB34
FB4B
FAE7
FA9B
FAE7
FB81
FBC3
FB8B
FB59
FB7C
FB99
FB3F
FAAA
FA78
FAB5
FAC3
FA86
FB16
FDAA
01C3
0528
061A
0527
045B
04CE
05A4
0596
04C2
0460
04FA
05B6
0599
04D9
046D
04AE
04FD
04D3
0483
049D
04FC
04FF
0495
0485
0546
05FF
0524
0224
FE37
FB49
FA51
FAB9
FB41
FB40
FAF6
FAEE
FB3A
FB76
FB51
FAF4
FAC4
FADE
FAFB
FAE9
FAE0
FB33
FBB6
FBDF
FB7D
FB0F
FB14
FB47
FB04
FA7C
FAFE
FD9A
019E
04EE
0610
057B
04B9
04A4
04D7
04BE
047D
048B
04E0
04FF
04CB
04BC
0528
0597
0554
0476
03E5
0445
0519
055B
04CF
0455
04BD
057E
04FA
0235
FE25
FAFB
FA1C
FAEB
FBAF
FB70
FABA
FA96
FB23
FB9B
FB72
FB07
FAFB
FB48
FB5F
FB11
FAD7
FB13
FB73
FB68
FB12
FB1B
FBA1
FBD0
FB01
FA09
FABC
FDF2
024C
055C
05ED
04F3
0439
048D
0550
0593
052E
04AD
0486
04AE
04E2
0509
0525
051A
04C4
044C
0426
048E
0518
051E
049E
0464
04FD
05A6
04BD
018E
FD6D
FAA4
FA39
FB1B
FB94
FB2B
FABC
FAFC
FB82
FB87
FB07
FAB5
FAE4
FB1F
FAF7
FAC5
FB21
FBDC
FC12
FB63
FA99
FAB9
FB97
FBFA
FB3D
FA6F
FB5F
FE99
029C
0546
05C9
051C
04A2
04C6
04F1
04A9
0445
046C
052A
05C9
05AD
0503
047A
0473
04AD
04CD
04D5
04F2
0509
04D0
0468
046F
051C
058E
0462
0138
FD65
FAD4
FA47
FAE6
FB65
FB57
FB2C
FB42
FB64
FB38
FADF
FAC3
FB05
FB46
FB31
FAEF
FAE8
FB27
FB47
FB0B
FACD
FB0A
FB9B
FBBA
FB0A
FA73
FB7B
FEA1
028E
052F
05AC
04F9
0489
04C8
0517
04FD
04CA
04F2
0541
0526
04A2
0468
04E6
0597
05AA
051F
04BD
04F3
0534
04CD
040C
03FC
04EE
05A1
0469
0109
FD2D
FADE
FAAB
FB78
FBD7
FB5E
FAB0
FA82
FADB
FB44
FB66
FB4B
FB20
FAF4
FACB
FAC2
FAF6
FB3B
FB2E
FABC
FA65
FAB9
FB8A
FBF6
FB82
FB02
FBF6
FEDE
0275
04D3
0546
04C4
0493
04EF
052E
04E7
047D
047C
04D4
050D
04F8
04E0
04FE
0517
04E0
048B
049A
051F
0580
0529
0465
041F
04B9
054A
0456
015B
FD8D
FADF
FA43
FB05
FBB9
FBAD
FB3D
FB07
FB16
FB14
FAF1
FAF9
FB46
FB77
FB3A
FADE
FAFB
FB8C
FBD9
FB68
FAC5
FAD8
FB96
FBEC
FB35
FA75
FB7F
FED5
02D1
0533
0556
047E
042C
0497
04FC
04EA
04C2
04EE
0537
0526
04CC
04B0
0501
0538
04D8
043F
0440
04FD
0587
050A
03FC
03BA
04BE
05A8
0480
00EA
FCC6
FA6A
FA6D
FB71
FBDD
FB72
FB03
FB1F
FB70
FB65
FB04
FAC7
FAD8
FAE9
FAC2
FAA7
FAEA
FB56
FB67
FB14
FAF8
FB82
FC2F
FC06
FB00
FA7B
FC04
FF97
036D
0594
05A7
04CF
0453
0475
04AF
04AC
04A5
04E1
053A
0556
052E
0512
052D
0544
0514
04C6
04BD
04FF
050A
0481
03D6
03E4
04C6
0548
03E7
0077
FC93
FA43
FA29
FB32
FBE7
FBD7
FB87
FB69
FB4C
FAE5
FA77
FA89
FB13
FB6C
FB24
FAA5
FAA1
FB17
FB54
FB05
FAC4
FB42
FC1E
FC32
FB33
FA8A
FC02
FFB6
03AE
05C6
05A2
04A2
042D
046C
04B8
04B9
04B5
04F4
0547
0558
0526
04FC
04FB
04F4
04C5
049D
04C1
0512
0513
048F
0405
042D
04F5
052F
038E
001C
FC7F
FA97
FAC3
FBB9
FC00
FB69
FAD8
FAEA
FB38
FB16
FA95
FA69
FAE0
FB70
FB78
FB15
FAE5
FB18
FB42
FB1E
FB0B
FB7C
FC13
FBF7
FB15
FAB8
FC58
FFE4
0398
0598
0596
04BB
043E
0459
0494
04AA
04D0
0533
058B
0574
04F9
0491
048E
04C2
04D1
04BA
04CD
0518
052B
04B1
0416
042A
04F0
0525
035C
FFB3
FC05
FA3A
FA83
FB6E
FBA5
FB2B
FAD6
FB02
FB42
FB25
FAE4
FAEF
FB3D
FB5E
FB2E
FB10
FB51
FB9E
FB70
FAE1
FAA5
FB1C
FBAE
FB7F
FAB9
FABE
FCD2
009C
043C
05F5
05AA
04AD
0443
048D
04E5
04E7
04DB
051B
0574
0561
04CD
0441
043D
04A3
04F1
04F3
04EC
050D
051A
04D0
047D
04B3
054B
0518
02FC
FF53
FBE7
FA54
FA94
FB53
FB78
FB1C
FAF6
FB3E
FB79
FB40
FACF
FAA8
FAE8
FB33
FB45
FB41
FB58
FB65
FB26
FAC6
FAD0
FB6D
FBF8
FBA7
FABA
FAA6
FCB5
008C
043C
05F7
05A0
049B
043D
04A2
0506
04F1
04B1
04C2
051B
0542
0500
04A3
048F
04C1
04E6
04E0
04DC
04ED
04CC
044D
03E6
044A
054B
0582
0383
FF91
FBBD
FA0A
FA85
FB85
FBA3
FB13
FAE0
FB58
FBBB
FB6D
FAD7
FAC4
FB37
FB72
FB1A
FAC3
FB13
FBBA
FBDC
FB52
FAFB
FB7B
FC30
FBF1
FACE
FA7B
FC8A
0080
0418
0587
0516
0470
049E
052A
0524
0480
0414
0469
050D
0533
04C5
046C
049B
04FF
0505
04AF
0489
04C3
04D9
0463
03E2
043D
054B
0573
0342
FF38
FB99
FA37
FAC7
FB90
FB7F
FB06
FB0D
FB8F
FBC6
FB5E
FAE3
FAF2
FB63
FB9A
FB72
FB5A
FB94
FBBC
FB65
FADC
FAE0
FB8D
FBFA
FB57
FA3E
FA73
FD18
0147
04B5
05D8
052C
045C
046A
04ED
050A
04A5
0460
0499
04ED
04DA
048B
048D
04EC
0506
0479
03D5
03F8
04D3
055F
04F3
0447
0486
058D
0599
0329
FEE3
FB32
F9E7
FA9D
FB85
FB7F
FAF8
FAE3
FB64
FBCD
FBAB
FB51
FB41
FB71
FB75
FB36
FB19
FB5C
FBA8
FB86
FB19
FB00
FB68
FBA6
FB15
FA43
FAC0
FD82
019E
04F0
060B
055C
046B
0437
048F
04CA
04B6
04A5
04CD
04F3
04CF
0482
046F
04B5
04FE
04EF
04A1
0480
04B6
04EA
04C7
0487
04B2
0527
04CE
0293
FED1
FB5B
F9E2
FA62
FB67
FBB5
FB61
FB2A
FB4E
FB66
FB2F
FAF8
FB15
FB51
FB46
FB09
FB0E
FB63
FB7C
FB05
FA86
FAC2
FB98
FC05
FB6E
FA9A
FB16
FD99
0143
045D
05CB
05A8
04E4
0461
046F
04C7
04FD
04ED
04BD
0495
0473
0465
04A1
0533
05B6
05AB
0527
04CB
04F0
0519
04AF
0410
0431
0508
0505
02BD
FEDA
FBA8
FAA6
FB1E
FB64
FAF0
FA92
FAE3
FB5F
FB55
FAFF
FB10
FB92
FBD2
FB6F
FADE
FAB5
FAE8
FB04
FAE8
FAD9
FAFF
FB2E
FB46
FB53
FB38
FAC5
FA64
FB42
FE1C
01FF
04DF
0587
04B4
0405
0440
04ED
055A
0565
0536
04DA
0472
045A
04B4
0516
050D
04D1
04EB
0552
0567
04F1
048D
04D0
0551
0546
04D1
04DA
055D
04D7
0213
FE0C
FB26
FA91
FB43
FB9E
FB51
FB1E
FB52
FB65
FB13
FAE5
FB3D
FB9D
FB61
FAD0
FAA9
FB01
FB32
FAED
FAAB
FAD5
FB1C
FB10
FAF4
FB43
FBA2
FB41
FA73
FAF8
FDEF
0210
04E1
0564
04D5
04BA
051F
0527
04AD
046B
04BB
0514
04FD
04C9
04E4
0512
04EC
04B0
04DF
054B
054D
04E6
04DA
056E
05BC
0504
0416
045B
0578
0519
01CF
FD40
FA79
FA89
FBB7
FC04
FB57
FAD7
FAFA
FB32
FB1E
FB19
FB55
FB63
FAFA
FAA1
FADF
FB55
FB4B
FAD5
FAA8
FAE8
FAF7
FA99
FA82
FB2E
FBCC
FB53
FA7E
FB78
FF0D
0335
0543
04E5
0413
0448
0500
0520
04BB
04AE
0512
0522
04A1
0455
04C5
0554
0543
04E3
0503
058F
05AE
0522
04AE
04E0
0530
04F7
049A
04E1
0546
0416
00B6
FCDB
FACA
FADB
FB89
FB9A
FB48
FB3C
FB5C
FB35
FAE7
FAF7
FB5B
FB75
FB1A
FAD8
FAF7
FAF6
FA7E
FA2D
FAB1
FB88
FB92
FAD3
FA95
FB75
FC3F
FBA2
FA8C
FB7C
FF41
0395
05A5
0539
045E
0485
0519
050F
0494
048A
0508
0545
04ED
049A
04CE
052C
052D
04FD
050D
0540
052A
04E4
04E4
0511
04C9
040A
03CE
04A5
0553
03E6
0039
FC7F
FADA
FB1D
FB8D
FB41
FACE
FADC
FB20
FB10
FADE
FB09
FB63
FB48
FAC1
FA93
FB0A
FB68
FB09
FA79
FAA0
FB55
FB9E
FB34
FAEC
FB53
FBB7
FB56
FB01
FC75
FFF8
0397
0546
0519
04B1
04F8
0560
0542
04EB
04EF
052A
0508
0495
047C
04F3
0566
0559
0518
050A
0500
04A4
044F
0490
0525
0529
047F
043B
04FE
0583
03C7
FFBB
FBCE
FA52
FAFD
FBB9
FB5A
FA99
FA88
FB09
FB4B
FB0F
FAD3
FADE
FAEA
FAC9
FAC1
FB04
FB43
FB35
FB16
FB35
FB55
FB1B
FACA
FAFD
FB83
FB63
FA6D
FA2F
FC71
00C7
0494
05CC
0505
0451
04A7
0545
0552
0502
04F1
0511
04FA
04C9
04FA
0575
057A
04CC
0432
046F
0531
0599
0579
054D
053E
04ED
0463
0461
051E
054B
033A
FF2C
FB80
FA33
FAD4
FB7C
FB38
FAB1
FAB6
FB13
FB2E
FB0A
FB16
FB54
FB52
FAFD
FAD2
FB10
FB4F
FB31
FAF7
FAF2
FAE6
FA86
FA40
FAC4
FBBD
FBEE
FB06
FAAB
FCCB
0103
04AE
05D2
0524
04AD
0520
0586
051E
0476
046D
04E4
0510
04BB
046D
0482
04B3
04C6
04F2
0555
0583
052D
04C1
04CC
0514
04F0
0479
048B
0537
0503
027D
FE57
FB09
FA25
FAD3
FB52
FB27
FB12
FB6A
FB9D
FB47
FAF1
FB2B
FBA2
FB98
FB17
FADD
FB28
FB5C
FB14
FACC
FB05
FB65
FB52
FB0B
FB3B
FBB3
FB80
FAA7
FAE4
FDC2
0244
0586
05DE
048A
03D5
0462
0516
0511
04B4
04A4
04C7
04AD
046F
0482
04DE
0503
04C9
0498
04AF
04C1
049D
049D
04F9
0532
04CB
044F
04A8
0579
04F2
01F0
FDC3
FAFB
FAA0
FB5E
FB90
FB27
FB04
FB4B
FB58
FB06
FAF2
FB64
FBBA
FB66
FADD
FAFB
FBA8
FBF4
FB85
FB0C
FB1C
FB47
FB07
FABD
FB13
FBA5
FB75
FAB7
FB38
FE36
0274
0549
058C
049A
0446
04BC
04FF
04B6
047D
04B1
04E2
04AB
0467
0498
050B
0523
04C8
047D
048D
04B2
04B9
04DC
0528
0525
049E
044F
04EE
05AC
04A6
0122
FCDC
FA5F
FA61
FB5F
FBBF
FB76
FB53
FB88
FB9B
FB69
FB53
FB70
FB5E
FAF5
FAB0
FAF4
FB66
FB68
FB10
FB09
FB7B
FBC6
FB8C
FB47
FB65
FB6E
FADC
FA76
FBDB
FF65
0344
0544
0521
0475
0482
04F1
04ED
0486
0460
048A
0488
044D
0467
0504
057E
053B
049B
0468
04B1
04C5
0464
0426
0479
04DA
04B5
0470
04C4
0538
042F
00ED
FCEC
FA81
FA6D
FB53
FB9C
FB2A
FAD9
FB10
FB64
FB7A
FB76
FB88
FB8C
FB55
FB0C
FAFE
FB35
FB7A
FBA7
FBB2
FB7F
FB11
FAD5
FB41
FBFE
FC00
FAF9
FA47
FBBF
FF75
035E
0559
0540
0498
048E
04F8
0536
053C
0550
0559
050B
0496
047B
04C6
04EB
0498
0435
0440
0492
04A9
048D
04B7
0526
0536
04B6
0473
04FE
0552
03AD
FFDE
FC01
FA5E
FB00
FBF4
FBC8
FAEB
FA8A
FADC
FB27
FB03
FAC7
FAC5
FADA
FAD8
FAF1
FB54
FBB4
FBA3
FB3E
FB0C
FB39
FB61
FB4C
FB44
FB78
FB78
FAFE
FADE
FC75
FFE4
037A
054F
0534
0494
049A
0512
0536
04F0
04C7
04FB
0545
0561
0562
0560
0541
04FB
04C2
04C1
04CF
04BF
04BB
04F5
051C
04AF
03F7
03FA
04ED
0557
0379
FF92
FBFA
FAA9
FB3C
FBC7
FB47
FA71
FA46
FAB6
FB10
FB25
FB43
FB6C
FB4B
FAE2
FAA8
FAD5
FB0C
FAFA
FAE4
FB26
FB72
FB37
FAAE
FAC0
FB90
FC12
FB9A
FB52
FD0E
00CF
0453
058D
04DD
0441
04BA
0570
0556
04B3
047C
04DD
0530
0517
04E5
04E7
04F8
04EF
04FA
0537
0552
04FC
048C
0495
04EA
04C9
0424
03F3
04A8
04FA
0325
FF4C
FBAF
FA47
FAC2
FB54
FB13
FAA7
FAD9
FB5E
FB7C
FB2D
FAF7
FB05
FB0F
FAF9
FAFB
FB1B
FB0D
FAC3
FAA7
FAF5
FB49
FB38
FB1E
FB91
FC2C
FBD2
FA93
FA66
FD0A
0194
051A
05D8
04E4
0469
0501
058F
0547
04C2
04CB
0524
0519
04B8
04A6
0503
054F
0541
052D
0543
052F
04BA
045F
04A4
051F
04F8
045B
046D
055E
0572
02E3
FE6C
FAD0
F9E3
FABF
FB52
FAEB
FA81
FAD2
FB5F
FB67
FB11
FAF8
FB20
FB18
FAD0
FAB0
FAD6
FAE8
FAC1
FAB7
FB00
FB3C
FB19
FAFA
FB6A
FBF1
FB8A
FA70
FA98
FD82
020D
055D
05ED
04E9
045A
04C0
0526
04F4
04B0
04E2
052D
0505
04A9
04B6
0523
0552
0510
04D9
04FF
0531
0517
04F4
0521
054E
04EC
0448
0460
053A
0531
02B4
FE72
FAEE
F9E4
FAB6
FB95
FB9F
FB45
FB1B
FB0F
FAEA
FAE8
FB45
FBAF
FBA5
FB30
FAD2
FACC
FAED
FB03
FB1F
FB42
FB31
FAE6
FACF
FB34
FB93
FB39
FA9A
FB4A
FE25
01F6
048D
050B
047D
0448
04A7
04FD
0510
052C
0555
0516
045F
03EB
0449
04FE
0522
04AC
0472
04EC
0591
05A5
0534
04C8
0487
0444
0438
04DF
05C4
053E
0239
FDEB
FAF3
FA98
FB91
FBD2
FAF4
FA40
FAA6
FB88
FBC7
FB4B
FAE7
FB13
FB70
FB89
FB77
FB84
FB9A
FB71
FB16
FAE6
FB01
FB17
FAF4
FAD9
FB11
FB60
FB3A
FAA5
FA81
FBCB
FE9F
01FE
048C
058C
0548
04B1
0487
04CD
04FE
04C7
0474
0482
04E7
051C
04DA
048A
04A9
050E
0524
04C2
046E
049D
050D
052A
04DF
0499
0492
048D
0471
048F
04E0
0468
0216
FE5A
FB38
FA4B
FB19
FBD1
FB84
FAEF
FB13
FBB7
FBDE
FB4E
FACA
FAE0
FB27
FB07
FABE
FAF5
FBA1
FBEA
FB6B
FADA
FB11
FBD3
FC21
FBA8
FB26
FB40
FB83
FB29
FA91
FB3F
FE12
01F4
04C2
056A
04BC
0436
0470
04E8
0509
04DF
04CD
04EF
0509
04F8
04E1
04EB
04FA
04DC
0499
0464
0452
043F
0419
0418
0474
04F5
0511
04A9
0461
04DF
05A2
051C
024D
FE2F
FB11
FA60
FB53
FC06
FB9B
FAE2
FAE2
FB73
FBA2
FB1B
FA91
FAB4
FB44
FB89
FB58
FB2D
FB50
FB74
FB54
FB3B
FB86
FBE2
FBA3
FAD7
FA72
FB0E
FBE7
FBC3
FAC7
FAC6
FD42
0173
04DE
05DC
0511
044D
046E
04DB
04D0
0474
046F
04DE
0536
0523
04F3
0503
051F
04DF
0463
044C
04D5
0564
054A
04A7
0446
0483
04DF
04CC
0495
04E2
0579
04FE
026C
FE87
FB68
FA75
FB20
FBC9
FB91
FAF4
FAC9
FB24
FB77
FB6B
FB33
FB13
FAF9
FAC7
FAAD
FAF0
FB6D
FBA5
FB66
FB16
FB27
FB70
FB68
FAFC
FAC3
FB2B
FBB8
FB94
FAE0
FB02
FD36
00FF
0458
05AB
053F
0499
04B3
052C
0537
04C3
0474
04A9
050C
0523
04FB
04ED
0503
04F2
04AC
0493
04DF
0532
050A
048E
0470
04E9
0551
0504
0465
046D
0521
050E
02CE
FEDF
FB6E
FA2D
FABB
FB6C
FB49
FAD6
FAE8
FB6D
FBA2
FB3A
FABE
FABB
FB11
FB43
FB35
FB34
FB5F
FB63
FB05
FA9A
FAA6
FB22
FB82
FB75
FB4E
FB6B
FB82
FB06
FA42
FA96
FD27
0154
04F7
0658
05B0
04A2
0464
04C9
0506
04E2
04C9
04FD
052B
04FB
04A2
0498
04DE
0508
04E8
04D9
0527
057A
0541
0493
0433
048B
050D
04FA
0485
049D
0563
0572
033C
FF13
FB34
F9A2
FA39
FB33
FB48
FACE
FABE
FB39
FB8E
FB57
FB02
FB13
FB5C
FB55
FAF9
FAD0
FB1C
FB67
FB30
FAB9
FAB3
FB3E
FBA6
FB5F
FAD4
FAD5
FB64
FBA1
FB2E
FB16
FCD6
0077
0425
05EE
05AB
04D6
04BC
053F
057E
0527
04BB
04B1
04E0
04E9
04D6
04EE
0525
051A
04BA
0478
04B0
0519
0523
04D0
04BD
052A
0577
04F9
0419
03FA
04D7
0537
035B
FF67
FB8F
F9EF
FA84
FB88
FB9B
FAFF
FAB8
FB05
FB42
FAFF
FAA2
FAB4
FB12
FB2A
FAE5
FAC7
FB25
FB9A
FB90
FB1D
FAE2
FB22
FB61
FB27
FABC
FACD
FB5C
FBA8
FB53
FB3D
FCC5
0016
03A4
059D
05A0
04D7
047D
04B4
04E1
04BB
049F
04E5
0557
0586
0562
0535
0521
04F4
049D
046E
04B4
052B
053A
04C4
045F
0491
0507
050A
048A
0451
04D2
0522
03C0
0065
FCA9
FA8B
FA78
FB2B
FB50
FAE0
FAA9
FAFD
FB57
FB38
FAD8
FAB4
FACE
FAC6
FA8E
FA93
FB0D
FB8E
FB8A
FB23
FB00
FB5A
FBA4
FB59
FAD6
FAE5
FB8A
FBD5
FB2F
FA87
FB98
FEE9
02F4
058A
05E5
0521
04BC
0513
056D
053D
04C6
049F
04E3
052E
053E
0539
0551
056B
0546
04E2
0486
045D
044F
0444
045F
04BD
051C
0510
04A9
048A
050D
056C
0442
011D
FD4E
FACC
FA52
FAD9
FB03
FAA0
FA81
FB18
FBC4
FBBB
FB12
FA92
FA9C
FACB
FAB2
FA8F
FAD5
FB5C
FB89
FB34
FAFA
FB5A
FBE5
FBCE
FB17
FAA5
FB01
FB87
FB57
FAD5
FB96
FE7F
0275
0550
05FF
0557
04CD
04E6
0524
0518
04F6
0509
052A
050C
04CC
04D6
0538
0576
052E
04A6
0471
04B0
04F2
04E2
04BC
04DA
0512
04E9
0462
0438
04E2
0595
04B6
0195
FD7B
FAA2
FA1F
FB01
FB90
FB24
FA7F
FA81
FB06
FB45
FAF5
FAA4
FAD3
FB44
FB61
FB16
FAE0
FB0D
FB56
FB62
FB4E
FB65
FB7D
FB2D
FA9B
FA8C
FB4D
FBFE
FB9B
FAA1
FB01
FDF4
024A
0572
061A
054B
04CB
0512
054E
04F2
047B
048C
04F3
050D
04CB
04BC
0519
055E
0514
048E
0475
04CB
04EC
048F
044A
04B5
0575
0599
04EA
045E
04D6
05AF
0525
0239
FDFB
FAA8
F997
FA3B
FB10
FB3A
FB04
FB09
FB5A
FB96
FB90
FB7A
FB75
FB51
FAEB
FA90
FAAD
FB2E
FB81
FB4B
FAEA
FAE7
FB30
FB2E
FABC
FA70
FAC5
FB3D
FB06
FA60
FAD5
FD95
01D1
053E
0650
059B
04D6
04E7
0549
0532
04AC
045B
0482
04CB
04E2
04E1
04FA
050A
04DA
0495
04AB
0520
056B
052E
04CF
04F6
0589
05AC
04F9
0440
0489
0572
0532
028B
FE6B
FB29
FA2B
FABC
FB41
FB12
FAC2
FAEB
FB4F
FB60
FB18
FAEB
FB0E
FB32
FB12
FAE4
FB02
FB51
FB61
FB0B
FAB2
FAB6
FAF1
FAF4
FAB8
FAB3
FB2A
FBA6
FB77
FAD5
FB13
FD5A
0130
049C
05F2
055C
046D
045B
04EE
053B
04F2
04A4
04CB
0524
052C
04E2
04BE
04F3
052A
050E
04C5
04AD
04D2
04EE
04EA
04F9
0532
0546
04FB
04AC
04E4
055F
04DC
0266
FE9E
FB73
FA53
FADE
FB90
FB7A
FAFD
FAE0
FB31
FB66
FB4A
FB3A
FB66
FB69
FAEB
FA58
FA74
FB41
FBD6
FB83
FAC7
FA9E
FB26
FB7E
FB1B
FA92
FAB2
FB3D
FB45
FABB
FAF9
FD44
0117
0466
05A4
052F
048E
04AA
0518
0507
046A
03F9
0444
0506
057F
0551
04DA
04AD
04E5
0526
052A
050F
0503
04FA
04E5
04E8
0523
0556
051E
04A8
04AC
054F
055F
035C
FF67
FB9A
F9F8
FA75
FB60
FB88
FB3A
FB40
FB92
FB98
FB3D
FB12
FB59
FB8D
FB38
FAB7
FABA
FB34
FB66
FAF7
FA77
FA91
FB14
FB3F
FAD1
FA6A
FAA8
FB34
FB2E
FA88
FA90
FCA0
007A
0428
05D3
0572
0493
0483
0513
054A
04E3
0487
04A6
04D0
0481
040B
042D
04EC
0570
0532
04B7
04C3
0538
054F
04DC
04A6
0532
05E2
05CD
0528
050A
05B0
05B6
039A
FFB1
FC12
FA7C
FAB6
FB3F
FB23
FABE
FAC1
FB27
FB61
FB3A
FB1A
FB61
FBDD
FC0E
FBC9
FB56
FB06
FADA
FAB8
FAB2
FADE
FB07
FADF
FA7E
FA63
FAC4
FB1E
FAD4
FA33
FA7C
FCAA
0044
03A2
055A
055A
04A8
0444
0469
04B8
04D1
04AA
047A
0476
049F
04D6
04FF
0502
04C7
0464
043D
04A8
0567
05CD
0592
053B
0566
05CE
059C
04B5
0436
04E5
059E
043D
0059
FC35
FA5E
FAEF
FBE2
FBBF
FB09
FAF1
FB89
FBED
FBC0
FB82
FB86
FB61
FAC7
FA41
FA74
FB24
FB8E
FB70
FB31
FB17
FAF9
FABF
FAA9
FACA
FAC6
FA65
FA2C
FAAE
FB7B
FB8C
FAF6
FB5C
FE04
01F2
04C9
055A
049C
0422
045D
04B9
04D4
04EA
0527
0545
0519
04F2
051B
0557
054A
050B
04ED
04E1
04A0
044E
0475
0529
05BB
0590
04FC
04CB
0514
0521
04AC
0470
0505
058C
0454
00E9
FCE8
FA72
FA1F
FAD0
FB3C
FB20
FAE8
FAC9
FAA1
FA6F
FA74
FAC2
FB1B
FB49
FB63
FB88
FB93
FB4F
FADA
FA8F
FA90
FAB1
FAE2
FB38
FB8A
FB66
FACC
FA7E
FB16
FBED
FBBF
FA9C
FA88
FD50
0200
0589
0615
04E0
044C
04F2
0588
0529
048B
04AA
0541
0565
050A
0503
0582
05B1
050F
045C
047F
0529
055E
04EE
0496
04C4
0508
04EC
04B3
04C3
04E5
04B3
0481
04D9
0517
039C
FFFD
FC26
FA62
FACF
FB9B
FB83
FB0D
FB2E
FBAE
FBA8
FB03
FA93
FABF
FAF0
FA9F
FA32
FA49
FAC2
FB12
FB27
FB4B
FB71
FB4A
FB00
FB24
FBB7
FBEE
FB59
FAC4
FB22
FBF7
FBDD
FACF
FAD8
FDA1
01F9
04F6
0541
0451
0434
0514
059B
0526
048C
04AA
052B
053F
04E1
04C0
0518
0568
054A
04FD
04EE
0514
0523
050F
0500
04E6
0495
0437
043B
04A0
04D3
048E
046A
04F1
055B
03FE
0065
FC5E
FA47
FA8F
FB7A
FB6E
FAA6
FA56
FAD8
FB67
FB78
FB62
FB90
FBB3
FB48
FA92
FA56
FAC4
FB33
FB21
FAE6
FAFE
FB45
FB50
FB27
FB23
FB48
FB4C
FB3F
FB80
FBEA
FBC0
FAF7
FB0B
FD8E
01DC
054A
0608
0509
046B
04CA
0516
04A7
043A
049B
0550
055A
04BF
0478
04EB
0560
053C
04DF
04DC
04FE
04D2
048F
04BC
0528
0526
04AE
047A
04D0
04F4
0460
03DD
0468
0535
040F
0039
FBE4
F9DD
FA73
FB8E
FB8F
FAE1
FAB1
FB22
FB71
FB4F
FB2B
FB47
FB48
FAFA
FAC7
FB05
FB4E
FB24
FACA
FAE2
FB67
FBAC
FB69
FB1A
FB2C
FB61
FB55
FB44
FB9D
FC0B
FBBB
FAD8
FB0A
FDA9
01D9
0530
062F
058B
04E4
04DE
04FB
04D6
04BB
04F8
053A
050F
04A2
048A
04EC
0554
055E
052A
04FB
04CB
047F
0448
046C
04BE
04CA
0483
0461
049B
04C3
0486
0459
04CE
053F
0407
007D
FC3F
F9CB
F9E7
FB0D
FB7E
FB17
FAC9
FAF0
FB15
FAF6
FAF2
FB3F
FB6A
FAFF
FA5C
FA42
FAC6
FB43
FB5F
FB6E
FBAB
FBB7
FB4E
FAE3
FB09
FB82
FBA8
FB6F
FB67
FB99
FB5B
FA9D
FACF
FD6E
01CD
054E
062D
0549
04A9
04FE
056A
0540
04E3
04DE
0504
04EB
04B8
04D6
052B
0532
04E5
04D7
053B
0578
051B
049A
0498
04E5
04DB
0480
0475
04D3
04E6
0460
0417
04CF
0595
045F
00A1
FC60
FA21
FA47
FB2A
FB68
FB26
FB18
FB35
FAFB
FA80
FA6C
FAFE
FB93
FB80
FAEB
FA7B
FA74
FA98
FAAC
FABE
FADC
FAF2
FB00
FB2E
FB77
FB91
FB5B
FB31
FB72
FBCA
FB83
FAC5
FAF5
FD53
0153
04D0
0619
0574
0474
043A
04AC
052A
0566
0565
0529
04C3
0485
04BA
0531
0576
0560
0536
052D
051C
04DB
04AD
04DF
0536
0535
04E3
04D2
051F
0524
0486
0400
0469
050D
0408
009C
FC8B
FA5F
FA9D
FB81
FB7B
FAEE
FB02
FBAE
FBDB
FB2A
FA80
FAAA
FB37
FB37
FA9D
FA43
FAA4
FB42
FB70
FB2D
FAE5
FAC9
FAC7
FADD
FB0A
FB1E
FB08
FB1D
FB9B
FC0A
FBA6
FAB7
FAD5
FD4C
014E
047E
0562
04BD
043E
0484
04F3
04FB
04CF
04C5
04D2
04D1
04EA
053D
057A
053A
04AC
0472
04BD
0509
04FB
04E8
0536
0590
0562
04D0
0498
04EB
051D
04BD
046F
04E9
056D
0430
00A6
FC9C
FA70
FA87
FB4B
FB5C
FAFA
FB07
FB7F
FB98
FB17
FAB6
FAFD
FB77
FB60
FAC8
FA72
FAC3
FB58
FB9C
FB6C
FB08
FABD
FABE
FB15
FB78
FB6D
FAE1
FA7C
FAD9
FB8B
FB82
FABC
FADA
FD59
0187
04F1
05F4
0545
04AE
04E1
052A
04EE
0488
047E
04AA
04A7
04A4
050B
05A7
05C3
052F
0492
0484
04CC
04DB
04A8
04A0
04D6
04E6
04BD
04C5
0520
0544
04E7
04B0
0538
05A3
042C
0068
FC3F
FA12
FA30
FAEB
FAEE
FA9E
FAE3
FB8B
FBAB
FB22
FABF
FB04
FB76
FB71
FB0C
FACF
FADC
FAEA
FAEB
FB21
FB7A
FB7D
FB11
FAD2
FB28
FB99
FB85
FB2D
FB4D
FBC2
FB93
FA9A
FA7A
FCE9
0151
0507
0629
0574
04D9
050E
054D
050E
04D6
052C
059A
0567
04C2
0488
04EF
053E
04EB
046A
0465
04C4
04FC
04F3
04F6
0506
04D8
047D
0474
04CE
04E4
045A
03F9
049E
057D
047F
00E2
FC97
FA44
FA63
FB30
FB29
FA93
FA64
FAAA
FAB8
FA80
FAA5
FB47
FBA1
FB3A
FAAF
FACA
FB53
FB86
FB49
FB2E
FB62
FB6E
FB1E
FAFF
FB70
FBDD
FB87
FAD4
FADC
FB9F
FBD3
FB02
FAD6
FD36
0191
0526
061A
054B
04BC
0504
053B
04DC
049B
050E
059C
0566
04AB
0464
04D7
0551
0547
04FF
04E5
04DA
0498
0456
047F
04E5
04E8
047D
0456
04C7
052A
04E7
0483
04CC
0530
03FA
007D
FC6B
FA36
FA68
FB5B
FB6B
FABA
FA5D
FAAB
FB14
FB3B
FB5C
FB99
FB93
FB0F
FA85
FA8E
FB11
FB69
FB55
FB35
FB4A
FB59
FB41
FB54
FBB1
FBCD
FB38
FA89
FAB8
FB99
FBDB
FB06
FABD
FCFB
0150
04F7
05F0
0516
048D
04F9
054F
04E9
0480
04D1
055D
0536
0486
0459
0505
05A4
057A
04EF
04BC
04C5
0489
042F
0452
04E7
0539
04FC
04C0
04EE
0503
0472
03CD
0419
04EC
0453
013B
FD24
FA9C
FA78
FB59
FBBC
FB7F
FB49
FB44
FB1C
FAD1
FACC
FB18
FB35
FAED
FAB6
FAF6
FB53
FB45
FAF0
FAD8
FB0F
FB2B
FB14
FB23
FB71
FB89
FB2D
FAF9
FB92
FC72
FC5E
FB4D
FB0A
FD38
0125
0459
0541
04A0
042C
0485
04FA
04F7
04D1
0509
0567
0554
04C4
044B
0450
049F
04D2
04D7
04DA
04EB
04FB
0516
0550
0585
056C
04FF
048E
0452
042A
03FB
040C
0499
04FC
03EE
00EF
FD38
FAC2
FA54
FAF6
FB54
FB2A
FB08
FB27
FB2E
FAEF
FACD
FB1A
FB86
FB8A
FB34
FB11
FB54
FB8F
FB6C
FB27
FB17
FB1A
FAE3
FA92
FA87
FACE
FB17
FB40
FB72
FBA8
FB8A
FB2C
FB90
FDB8
0136
0440
0580
0556
04FC
04FE
050E
04FD
050D
0552
0565
04FA
046E
044F
0496
04CA
04C7
04E1
0534
0552
04F7
0491
04A1
04FC
0525
0510
0514
0524
04D2
042A
03FC
04B9
0560
043F
00F2
FD1F
FAD8
FA95
FB29
FB58
FAF9
FA98
FA94
FAD4
FB0D
FB19
FB0A
FB07
FB1E
FB3B
FB43
FB36
FB21
FB05
FAD8
FAA5
FAA3
FAF0
FB4D
FB56
FB0F
FAE7
FB1D
FB6F
FB8F
FB9D
FBDB
FC0E
FBBD
FB21
FB66
FD90
0127
0467
05D6
0592
04E3
04C3
0515
053C
0502
04C4
04DA
0525
053D
04FE
04B9
04C8
050F
0531
0516
0505
0523
0533
0500
04C0
04C7
04F9
04EA
048E
046D
04D4
0535
04DD
0423
0424
050C
0550
034B
FF54
FBA9
FA21
FA8C
FB5D
FB80
FB21
FADE
FAE1
FAF0
FAF4
FB0F
FB41
FB50
FB25
FAF1
FAF6
FB34
FB65
FB45
FAF1
FAD1
FB1B
FB6E
FB3F
FAA6
FA63
FAD9
FB74
FB63
FAD0
FAB6
FB6D
FBF8
FB6C
FAAD
FBCD
FF77
03BE
060C
05DD
04D5
0492
0515
0574
0544
04E3
04B3
04A0
0483
047E
04B8
0503
0512
04EA
04D1
04E7
0510
0526
0518
04E7
04B8
04B9
04E5
0502
04F7
04E8
04EB
04D1
048B
0481
051D
05C7
04EE
01B0
FD57
FA6D
FA1F
FB1E
FB77
FAD2
FA59
FAC2
FB6F
FB87
FB2E
FB22
FB84
FBAF
FB37
FA8C
FA5E
FAB7
FB16
FB38
FB4B
FB78
FB91
FB5D
FAF9
FAC7
FAF7
FB4B
FB58
FB15
FAF5
FB4A
FBA5
FB48
FA5B
FA50
FC88
0099
045C
05F7
05A0
0501
0518
0563
0521
0499
049C
0530
0581
0515
0470
0453
04BD
0512
0500
04D7
04F4
0530
0531
04FA
04DD
04EA
04D3
0467
03F9
040E
04AF
054B
055B
0513
0537
05EA
0606
0419
0037
FC54
FA6F
FA9E
FB46
FB27
FA8C
FA71
FAEE
FB37
FAE8
FA9C
FAEF
FB91
FBC6
FB75
FB29
FB2B
FB2D
FAEA
FAA2
FAB7
FB18
FB55
FB39
FB08
FB0A
FB24
FB0F
FAD3
FAC5
FB15
FB76
FB63
FABC
FA40
FB3B
FE49
0255
0542
05E0
050B
0482
04F4
0590
0573
04DD
04A8
04FE
0538
04F5
04A7
04C9
0517
050D
04C1
04B8
0507
0539
0506
04C6
04D9
0519
0517
04D5
04D0
0539
058A
052C
045E
040F
04B5
058B
0519
0290
FEBB
FB7E
FA3D
FAB0
FB67
FB66
FAF8
FAD8
FB12
FB17
FAC1
FA9D
FB0E
FB95
FB70
FABE
FA6B
FAE6
FB88
FB90
FB2D
FB18
FB6A
FB83
FB16
FAB3
FAF1
FB80
FB88
FAE8
FA7D
FAF4
FBC2
FBC2
FADD
FA87
FC4D
0010
03ED
05F1
05CF
04DA
047C
04EA
055D
0549
04F2
04D8
0503
0522
050F
04F2
04E9
04E5
04E3
050A
055D
0581
051F
0470
0417
044D
0498
0484
0454
0499
0543
0592
0515
0462
046F
054D
05C0
0457
00F4
FD19
FA9E
FA1E
FAB2
FB0D
FACB
FA83
FAC6
FB4F
FB6F
FB09
FAB4
FADA
FB2F
FB3D
FB17
FB1E
FB4E
FB40
FAE2
FABA
FB28
FBBB
FBB6
FB21
FACA
FB1E
FB8E
FB6B
FAF5
FAF8
FB86
FBC0
FB1B
FA6F
FB46
FE23
01CB
0468
053B
0509
0500
0583
0602
05E0
0532
0496
047A
04A8
04B5
04A0
04C0
0520
0552
050F
04AE
04B0
0502
0511
04AB
0454
048B
0508
0519
04A9
045F
049B
04E0
04AA
045C
04C2
0597
054F
02BC
FEA8
FB50
FA36
FADA
FB9D
FB93
FB10
FAC8
FAD6
FAE1
FAC8
FAC3
FAF2
FB1D
FB0B
FAE0
FAEB
FB33
FB5C
FB35
FB06
FB33
FBA3
FBD4
FB93
FB45
FB4C
FB75
FB46
FAD6
FAD4
FB84
FC17
FB8D
FA41
FA08
FC50
0069
0402
056D
050C
0480
04C2
0568
0593
0525
04C1
04DB
052F
0537
04E8
04B4
04E6
053C
0544
04F3
04AC
04B2
04CA
04A0
0448
042B
046B
04B0
04AA
0489
04A3
04DF
04CC
046F
046B
0520
05B2
04A0
016C
FD76
FAC3
FA25
FABA
FB2F
FB13
FAD6
FADE
FB0F
FB1C
FB05
FAFF
FB10
FB0E
FAEC
FAD8
FAF7
FB29
FB39
FB2D
FB3D
FB76
FB97
FB65
FB0E
FB03
FB5C
FBAE
FB90
FB3C
FB4E
FBD8
FC10
FB4A
FA2A
FA6C
FD21
014E
04AC
05CA
053E
04AC
04EE
057F
0590
051E
04C9
04E4
051A
0506
04C6
04BC
04F7
0525
0514
04FC
051B
054D
0537
04D5
0490
04AD
04E4
04C0
044E
041A
0469
04C7
04AA
0450
0480
054F
057D
03A3
FFE8
FC36
FA6A
FA95
FB3D
FB2E
FA97
FA54
FAA7
FB08
FB08
FAD9
FAD9
FAF9
FAED
FABE
FAC4
FB15
FB4C
FB14
FAB2
FAAE
FB12
FB5C
FB39
FAFD
FB24
FB97
FBC3
FB6F
FB22
FB69
FBF5
FBDB
FAEA
FA58
FBBC
FF46
0341
0594
05B3
04E2
04A4
0532
05A8
0563
04C9
049D
04FC
0560
0568
0545
0540
0541
0504
04AC
04AA
0512
056B
054D
04ED
04C3
04D3
04B9
0458
0425
0476
04E6
04C7
0423
03E4
049C
0577
04CF
01F3
FE05
FB01
F9FA
FA68
FB0C
FB31
FB02
FAE6
FAE9
FAD8
FAB1
FAAE
FAE9
FB28
FB28
FAF5
FAD1
FAD4
FAD3
FAB7
FAB5
FB06
FB7D
FBAF
FB81
FB58
FB82
FBC0
FB95
FB11
FAD6
FB44
FBD1
FBA8
FAEC
FAF8
FD16
00F1
0498
0638
05BD
04AA
046A
0502
0575
0527
0498
049A
0534
05AA
0585
0523
0513
0543
0532
04C6
047D
04AC
04FB
04E6
048D
047F
04D4
0503
04BF
0478
04A8
04FC
04C2
0421
0414
04F5
0580
03F6
0037
FC35
FA0D
FA0E
FADB
FB36
FB1A
FB1C
FB60
FB7C
FB30
FACA
FAB5
FAEB
FB0B
FAEB
FAD3
FB04
FB48
FB31
FAC0
FA7D
FACD
FB64
FB9F
FB5A
FB21
FB60
FBB7
FB82
FAE4
FAC1
FB73
FC1A
FBBC
FADB
FB4F
FE34
0267
0580
0634
055E
04AA
04BF
0506
04DF
0483
047F
04DE
0529
051B
04F2
0501
0531
052C
04ED
04D0
050A
054F
053C
04EF
04DB
050C
0505
0480
03F9
0422
04D4
051F
048B
03E6
0443
054E
0544
02D6
FECE
FB5D
FA02
FA69
FB36
FB7A
FB3D
FAF8
FAED
FB04
FB14
FB0E
FAFB
FAE9
FADD
FAD8
FADD
FAF4
FB18
FB2A
FB15
FB05
FB2A
FB5F
FB4E
FB00
FAEE
FB4D
FBA6
FB77
FB0E
FB2D
FBD1
FBFB
FB2C
FAA9
FC5C
005B
0450
05E8
0538
0437
043E
04E4
052E
0501
04F5
0537
055C
052B
0502
0530
0569
053C
04CD
049B
04C3
04E4
04C1
048F
049A
04D6
04F9
04EA
04E2
0511
054A
0524
047F
03D9
03E6
04B9
054D
0439
011A
FD43
FAB3
FA3D
FAEF
FB60
FB2D
FAF0
FB1C
FB65
FB5B
FB10
FAE9
FAFC
FB04
FADA
FAB8
FAD4
FB05
FB09
FAF1
FB0B
FB68
FBB6
FBAF
FB71
FB4F
FB61
FB6C
FB3B
FAF8
FB03
FB62
FB9E
FB5C
FB1B
FBF4
FE7B
01E3
0491
058A
0535
04A9
0484
049B
04AB
04C3
04FB
0516
04DA
047E
047B
04EA
0561
0570
051D
04C3
04A0
04AA
04BA
04C1
04BF
04AE
0490
047F
0498
04CF
04EE
04C6
0468
0436
048E
052A
04ED
02CE
FF2E
FBD8
FA64
FAB2
FB58
FB58
FAFD
FAFE
FB56
FB73
FB37
FB1E
FB57
FB6C
FB16
FACD
FB15
FB94
FB90
FB03
FAAE
FAF3
FB50
FB35
FAF2
FB3D
FC00
FC4E
FBA9
FAC5
FA8E
FAFA
FB4D
FB3E
FB37
FB73
FB8C
FB2E
FAE9
FBDB
FE78
01E3
0496
05A9
0561
04B8
0474
04AD
04F6
04F7
04C6
04BF
04F6
0521
0502
04C3
04B3
04DC
050D
051D
050C
04DC
0490
044F
0452
04A2
04F7
0506
04E0
04C6
04C3
04AC
0484
048E
04CE
04E2
049F
047D
04EE
055E
0463
0150
FD4D
FA79
F9EF
FAE8
FBC7
FBC7
FB55
FB1F
FB38
FB3F
FB00
FAAF
FA96
FABD
FAF7
FB27
FB56
FB92
FBBD
FBB3
FB79
FB3D
FB14
FAF5
FAE3
FAFC
FB3C
FB6F
FB67
FB3D
FB2E
FB41
FB48
FB3B
FB51
FB87
FB64
FABD
FA87
FC31
FFD8
03A5
058C
055F
04B9
04E4
0590
05B9
0536
04CB
04E4
0510
04E3
04A5
04C9
051E
0522
04E0
04D6
0523
054C
04F9
047F
0462
049C
04BD
04AF
04C9
0523
0545
04E0
046C
048E
0518
0533
049B
0429
04B5
05B0
055E
02A5
FE6E
FAFC
F9CE
FA69
FB38
FB46
FAE1
FABC
FAED
FB04
FAD7
FAC8
FB20
FB7D
FB4F
FAAC
FA4C
FA96
FB23
FB62
FB55
FB5A
FB7E
FB6F
FB1D
FAE7
FB08
FB2E
FAFD
FABB
FAF9
FBA4
FC03
FBBF
FB6F
FBA4
FBEA
FB76
FAB8
FB62
FE78
02BA
05A9
0619
0529
04A8
050D
0571
0532
04C7
04E7
0571
05A7
0544
04CA
04C2
050A
051E
04DB
0499
049F
04C9
04DD
04EC
0513
0521
04CF
044C
0423
0481
04E7
04DB
0492
0497
04DD
04BD
0412
03B8
0457
0500
03D2
004C
FC49
FA2E
FA69
FB5B
FB7E
FAED
FAA2
FAE4
FB1B
FAF2
FACF
FB0E
FB60
FB48
FAEE
FAE0
FB30
FB65
FB37
FAF6
FAFE
FB2B
FB24
FAF8
FB0B
FB69
FB9A
FB58
FB0D
FB46
FBD1
FBF7
FB81
FB1B
FB64
FBF1
FBD0
FAF9
FAD1
FCC9
0095
042F
05CF
058F
04F0
04F9
0554
0534
04A0
045C
04BF
053B
052F
04C7
04B2
0516
0566
053D
04F2
04FE
053A
051D
0497
043D
0473
04E2
04F8
04B5
0489
049A
049D
0473
0479
04DE
052C
04E1
045C
047D
052D
04EE
026C
FE56
FAFE
F9FD
FAAD
FB42
FAF8
FA91
FAE1
FB8F
FBAF
FB1E
FAA1
FAC7
FB36
FB4D
FB10
FB01
FB46
FB73
FB37
FADB
FAD7
FB22
FB4E
FB32
FB16
FB29
FB37
FB15
FB01
FB47
FBA6
FB93
FB10
FAD4
FB48
FBD4
FBA7
FB29
FBEB
FED6
02CF
05A7
064D
05A0
0518
0528
0540
04F7
04A2
04B1
0501
051D
04EE
04C5
04CE
04DE
04CE
04C9
04FF
054A
0557
0520
04F2
04F6
04FA
04CB
048B
0483
04A5
049E
0463
0456
04AB
04ED
048C
03CE
03B8
04AE
0578
043A
0088
FC35
F9A7
F99B
FABB
FB57
FB10
FAA8
FAB8
FB0E
FB38
FB31
FB35
FB41
FB1D
FAD3
FABC
FAFC
FB43
FB3C
FB08
FB08
FB4A
FB77
FB5F
FB3D
FB49
FB57
FB27
FAEF
FB20
FBAA
FBDF
FB68
FADF
FB0C
FBB4
FBCA
FB15
FAFC
FD17
0117
04BA
061F
059E
0502
054D
05E0
05C1
04FD
046B
047B
04D2
04FE
0509
051F
051A
04CA
046C
046E
04CA
0502
04D1
0498
04CD
0549
057B
0534
04DB
04C3
04B6
046B
0420
044A
04C6
04E1
0463
0416
04BF
05B6
0525
01FC
FD6D
F9F7
F911
F9FB
FAF4
FB17
FAD4
FAD9
FB1B
FB28
FAE9
FAC4
FAFB
FB52
FB6C
FB45
FB20
FB20
FB27
FB24
FB2C
FB44
FB3F
FAFD
FAB1
FAA9
FAE6
FB22
FB34
FB44
FB74
FB8E
FB5C
FB1A
FB42
FBCB
FC05
FB90
FB41
FC8C
FFD8
03B5
060A
0613
04F1
0449
04A9
055B
0589
052B
04CA
04B9
04D3
04D9
04C9
04C1
04BC
04A1
047C
047C
04B2
04F4
0512
0515
0520
0534
0536
0524
0514
04FB
04B6
0458
0436
0473
04A4
044E
03C1
03E7
04F5
0589
03D8
FFD2
FB9F
F995
F9F8
FB12
FB4F
FABC
FA5F
FAB6
FB4C
FB92
FB87
FB6F
FB5A
FB37
FB22
FB39
FB4F
FB21
FACC
FAC2
FB2A
FB98
FB95
FB3D
FB10
FB38
FB59
FB2C
FAF6
FB20
FB8B
FBB3
FB77
FB59
FBAD
FBFA
FB8E
FAC7
FB2D
FDDF
0206
0554
0632
0538
044B
0480
054D
059F
0541
04D0
04BE
04D8
04C9
04A9
04B9
04E7
04E7
04B8
04AA
04DB
04FF
04DC
04AA
04BE
04FA
04F0
048C
043B
044E
048C
049B
0497
04D4
052A
0500
0443
03D2
046B
0553
04B6
01A9
FD73
FA6E
F9C8
FA99
FB3A
FB05
FA8E
FA85
FADE
FB26
FB38
FB43
FB53
FB3F
FB06
FAF1
FB2C
FB74
FB6F
FB29
FB01
FB1E
FB3D
FB28
FB1B
FB61
FBBF
FBB4
FB44
FB0F
FB6E
FBE6
FBD5
FB6D
FB6A
FBD6
FBC8
FAD1
FA2E
FBBB
FFA5
03D2
05F6
05D3
0505
04E7
0561
05AB
0580
0534
04F4
049E
0442
043F
04B6
0538
0553
0524
050E
050C
04C8
0446
0411
0477
0505
050C
048E
042E
0445
046B
042F
03E4
0437
0514
057F
04E1
03FB
040F
051E
0579
0375
FF66
FB84
F9CB
FA3A
FB3F
FB8B
FB1D
FAB1
FAB2
FAED
FB17
FB26
FB2E
FB2B
FB18
FB0B
FB17
FB22
FB0D
FAF6
FB14
FB5F
FB84
FB59
FB1E
FB24
FB52
FB57
FB30
FB3B
FB9F
FBF4
FBCE
FB6E
FB80
FC0F
FC37
FB4C
FA1F
FA8F
FD8C
01D5
0501
05C3
04EC
0441
04A0
0579
05DE
0598
051F
04D4
04A8
0478
045B
047C
04C9
0501
0505
04ED
04D8
04C9
04BD
04C9
04F0
050C
04F2
04B9
04A0
04B2
04B2
0484
0465
0487
04AA
0467
03EC
03F8
04CE
056C
044D
011C
FD59
FAFC
FAA5
FB4A
FB94
FB2F
FAAC
FA8B
FAB9
FAE9
FB09
FB34
FB62
FB67
FB39
FB09
FAF7
FAEF
FACF
FAA5
FAA6
FAE1
FB2E
FB5B
FB5F
FB51
FB3C
FB23
FB1A
FB42
FB92
FBC7
FBBA
FB9A
FBA7
FBBC
FB6E
FAD4
FAF2
FCE3
0080
041B
05F1
05CF
0508
04DD
0546
0574
0510
0498
048E
04D4
04FE
04F2
04E9
04EF
04CF
0483
045C
0491
04E7
0504
04FB
051E
056B
0579
0517
04A8
0497
04B7
048B
0421
0417
04A4
0518
04C4
0412
0412
04D3
04D9
02BB
FEFD
FBB9
FA63
FA71
FA71
F9F3
F9BB
FA5A
FB40
FB8A
FB2F
FAE9
FB22
FB80
FB8B
FB5D
FB57
FB7C
FB79
FB36
FAFA
FAF5
FAFE
FAF5
FB0A
FB67
FBBA
FB91
FB0C
FADC
FB4D
FBC6
FBA3
FB31
FB52
FC11
FC5C
FB85
FA9B
FB85
FEB7
026F
0491
04DA
04B6
053F
0615
064A
05D5
056E
0568
054C
04BE
0427
0425
049D
04DF
04A4
0464
0498
050F
0539
04EB
0480
044D
044E
046D
04AF
04FE
050A
04B7
0470
04A5
0512
04F3
0421
0384
03F7
050B
0577
04CF
0422
0471
04FF
03F7
00BA
FCE3
FA9D
FA61
FADC
FAD3
FA6E
FA6E
FAE3
FB2C
FB0D
FAFC
FB58
FBC5
FBB9
FB51
FB26
FB6A
FBA8
FB7A
FB1D
FB02
FB29
FB35
FB0B
FAF1
FB0A
FB1F
FB08
FB03
FB48
FB8B
FB58
FAD2
FAA8
FB15
FB78
FB40
FADE
FB37
FC31
FC97
FBCC
FB10
FC54
FFD0
0382
054B
0517
047C
0497
050F
0521
04E1
04EF
055D
0585
0509
0462
0433
0475
04A8
049D
04A2
04DB
0501
04D3
048C
0490
04DB
0514
051B
0520
052E
0504
0497
0461
04C6
055E
055D
04AF
0429
0460
04CB
0494
03FE
042C
0547
05A3
037C
FF49
FB99
FA65
FB1C
FBBD
FB4A
FA8D
FA80
FAEF
FB04
FAA3
FA7D
FAED
FB6F
FB63
FAF0
FAB3
FAE8
FB37
FB52
FB4B
FB40
FB1A
FAD9
FACE
FB2C
FB94
FB79
FAEF
FAA7
FB02
FB80
FB7C
FB1B
FB09
FB5B
FB6A
FAEF
FAA4
FB3A
FC0D
FBCE
FA8F
FA54
FCEA
0180
0537
0629
0533
0480
04E8
057C
054A
04B3
04A6
053B
05AE
0586
051D
04F0
04F5
04E9
04DB
04FE
0526
04F0
0473
0448
04BC
054F
0553
04CF
0462
045A
046A
045A
0477
04FA
0569
051D
0450
03F9
0478
0502
04CA
044F
04AC
05AC
0567
0270
FDEB
FA9D
FA0A
FB0C
FB8C
FAE6
FA17
FA00
FA53
FA64
FA44
FA83
FB28
FB9E
FB8E
FB4D
FB3A
FB34
FAF4
FAAB
FAD0
FB53
FB94
FB42
FAD5
FAEA
FB63
FBA4
FB71
FB31
FB34
FB3D
FB0C
FAEB
FB45
FBD8
FBE4
FB48
FACD
FB09
FB71
FB2D
FAB1
FBA6
FEE4
0301
0599
05D0
04FC
04C6
054A
0588
051A
04B4
04F7
0584
0596
0522
04CA
04E5
0514
04EE
0497
046E
0475
046A
045A
0494
0514
0557
0507
0481
045D
04A7
04E2
04C7
049C
04A4
04A6
045A
0403
0420
0499
04CE
048A
0475
0502
054E
03CB
003C
FC71
FA82
FAA8
FB47
FB0B
FA47
FA0D
FA95
FB0E
FAE4
FA7F
FA88
FAF8
FB43
FB38
FB2C
FB60
FB9A
FB90
FB5E
FB4D
FB60
FB5D
FB3C
FB34
FB57
FB66
FB40
FB2E
FB74
FBD5
FBD2
FB6A
FB2D
FB6B
FBB7
FB90
FB30
FB43
FBC6
FBE7
FB51
FB1F
FCCC
004E
03C8
0574
056A
051D
0570
05DC
0593
04C6
0451
048E
04FB
050E
04E6
04EB
0522
0538
050E
04DC
04CB
04BB
049C
049E
04E5
052D
0515
04AA
0454
0442
043F
042B
0452
04E6
0576
054F
047C
03E1
0419
04A7
04B7
0462
0485
053A
0524
02DF
FEE8
FB71
FA25
FA9C
FB39
FB27
FADE
FAFD
FB51
FB47
FADC
FA93
FAB1
FAEF
FB0A
FB1F
FB53
FB6C
FB24
FAAD
FA8B
FAE0
FB3F
FB47
FB21
FB26
FB52
FB57
FB2F
FB2B
FB5B
FB58
FAEC
FA8B
FAC9
FB71
FBB0
FB44
FAE8
FB41
FBCA
FB86
FAB5
FB12
FDD9
0202
0510
05A9
04C4
0432
0495
052D
0544
050C
0500
0514
04F3
04B0
04B8
0512
0540
04F2
047E
0466
04A2
04BE
0492
0475
04A2
04DB
04D2
04AA
04B6
04E7
04E4
04A8
04A1
0504
0561
053E
04D7
04C8
0506
04D9
0407
0385
043C
0566
04F0
01DE
FDB3
FB00
FAAE
FB61
FB75
FAD9
FA98
FB16
FB89
FB35
FA74
FA25
FA8B
FB20
FB6D
FB84
FB94
FB7F
FB23
FABF
FAB4
FAF7
FB25
FB16
FB11
FB50
FBA0
FBB7
FBAA
FBBA
FBCC
FB7D
FADA
FA85
FAE1
FB70
FB78
FB11
FB04
FB83
FBB0
FAF1
FA53
FBBD
FF94
03CF
05F3
05A1
04A4
049C
054D
0582
04EA
046B
04BF
0578
05AC
052D
0498
046D
0493
04B7
04CA
04E3
04FA
04F8
04F2
0502
0505
04C2
0459
0441
04A0
0501
04EB
048D
047D
04D8
0516
04DE
0496
04BF
0515
04E0
042F
03FD
04C3
054F
03D0
0013
FC17
FA08
FA16
FAAF
FA9A
FA2B
FA50
FB0A
FB7C
FB31
FAAC
FAA1
FB0B
FB5D
FB4D
FB13
FAF6
FAF0
FAE5
FADD
FADE
FAC9
FA91
FA76
FAB7
FB23
FB42
FAF3
FAA9
FACA
FB26
FB47
FB2C
FB44
FBA8
FBD7
FB77
FAFC
FB15
FB95
FB98
FAED
FAD2
FCBA
0060
03C7
053E
050A
04B0
0511
05B0
05C8
056A
0531
0549
0548
04EF
0490
0490
04D3
04F8
04EF
0500
0549
058A
0585
055A
0547
054B
053D
051D
0516
0520
04FF
04AA
0477
04A3
04E8
04E1
04AA
04C4
053F
0575
04F5
0456
048F
0566
0535
02AF
FE9A
FB3E
FA1B
FAA0
FB40
FB4A
FB34
FB76
FBC0
FB94
FB17
FADC
FB0E
FB40
FB1A
FAD5
FAD2
FB08
FB21
FB01
FAE7
FB02
FB2D
FB36
FB27
FB28
FB31
FB26
FB15
FB22
FB35
FB0A
FAB3
FAA9
FB29
FBB5
FB9C
FAFF
FABC
FB36
FBA2
FB1F
FA48
FAF5
FE18
0252
0528
058D
04B0
0451
04D1
0547
050D
0488
046A
04B6
04EC
04CE
0495
047B
046C
0455
0460
04B3
0519
053B
0516
04F2
04EF
04E0
04A8
0478
0481
04A1
0498
047F
04B0
0525
055A
050D
04B6
04E8
055C
053B
0466
03E8
0495
0585
04B8
0163
FD2C
FA8B
FA4B
FB15
FB55
FAEC
FAC1
FB36
FBAB
FB7D
FAE1
FA7F
FA9A
FAEF
FB3B
FB7E
FBB2
FBB4
FB85
FB63
FB71
FB69
FAFA
FA5C
FA2B
FA9C
FB37
FB71
FB58
FB55
FB79
FB74
FB33
FB15
FB4E
FB7F
FB3B
FAD2
FAF7
FB98
FBB5
FAD6
FA33
FBB2
FF9C
03E9
0635
061A
0529
04D5
0508
04EE
0468
0423
047F
0502
0516
04D1
04B0
04D8
04FA
04E7
04CF
04DB
04DF
04B8
04A0
04E6
055C
057B
0520
04C1
04D0
051F
0534
0500
04E2
04FA
04F0
0491
043E
0460
04BD
04C7
049B
04F2
05D5
05E1
038F
FF42
FB5B
F9E9
FAA3
FB96
FB7F
FADC
FABD
FB33
FB7E
FB4C
FB21
FB67
FBC4
FBA9
FB36
FB08
FB4D
FB82
FB31
FA98
FA46
FA62
FA9F
FAC3
FAE9
FB1F
FB32
FB05
FAD6
FAEA
FB15
FAFA
FAA8
FA9A
FB00
FB6D
FB73
FB50
FB80
FBD2
FB8C
FABF
FAD5
FD29
0128
048A
05A2
0500
0473
04CC
0542
04F7
044D
0440
04EE
056F
0524
0482
0453
04A2
04CC
0486
0439
0450
0498
04A3
047A
048B
04FC
056D
0578
052A
04D6
04A7
0499
04B3
04F6
0524
04EF
047C
0456
04B7
051D
04FC
049D
04BF
053C
04AB
01EB
FDCF
FAA5
F9DB
FAA5
FB3C
FAFF
FAC7
FB4A
FBFF
FBED
FB1A
FA81
FAB8
FB40
FB5C
FB1B
FB19
FB80
FBC9
FB94
FB33
FB2D
FB7D
FBA9
FB7A
FB3F
FB4B
FB7C
FB87
FB66
FB51
FB5B
FB5C
FB40
FB24
FB18
FB0B
FB09
FB4A
FBC1
FBDC
FB36
FA95
FB95
FEE8
0322
05DE
061F
0522
04B5
0533
058E
0516
0466
0464
04F5
0536
04CD
0452
0460
04B7
04B7
0456
042A
0484
04FB
050F
04DF
04E0
051E
0529
04C1
0440
0423
046E
04C2
04E7
04FA
0517
051E
04EE
049B
044A
0404
03E0
0421
04DD
0592
0588
04C1
042C
0472
04C4
037A
000D
FC16
F9CE
F9D7
FADA
FB54
FB1D
FAFF
FB47
FB78
FB38
FAF9
FB41
FBD0
FBE8
FB57
FABC
FAA7
FAEC
FB02
FADD
FAE8
FB4D
FB9E
FB77
FB0A
FADC
FB11
FB50
FB4B
FB17
FAF0
FADD
FACB
FAC8
FAE6
FB04
FAF3
FAD3
FAFF
FB7C
FBCE
FBA2
FB5A
FB8B
FC0F
FC14
FB6E
FB50
FD27
00BF
041D
0579
04FC
043A
043C
04A3
04B0
0471
0483
04FF
0549
0501
0492
0498
0503
0543
051F
04F4
0512
053C
0511
04B1
049A
04F3
0554
0556
050F
04D8
04CB
04C4
04B9
04CA
04F0
04E7
0495
0446
0444
0468
0455
0415
041A
0484
04D2
04A4
0472
04F2
05C1
054B
027F
FE5B
FB31
FA57
FB04
FB8E
FB55
FAF8
FB04
FB2A
FAEC
FA78
FA68
FAD1
FB27
FB0A
FAC9
FAD2
FB02
FAE1
FA67
FA19
FA4D
FAB8
FAE1
FAC9
FACE
FB12
FB4F
FB4D
FB37
FB47
FB64
FB53
FB24
FB23
FB60
FB94
FB93
FB91
FBB7
FBC2
FB5E
FACF
FABE
FB38
FB63
FAAF
FA09
FB36
FEBE
02F8
0590
05D9
0524
04EF
0553
0582
052F
04E3
0507
0541
0517
04BD
04CA
0557
05D4
05D7
059E
0594
05A1
055D
04D0
047E
04BA
0532
0562
053A
050F
050A
04FE
04CD
04A1
04A3
04AE
0499
048A
04B9
04F8
04E1
0478
0450
04BC
0535
0504
0462
0450
0511
054E
0363
FF73
FBA2
F9F4
FA59
FB1D
FB05
FA61
FA1D
FA67
FAAE
FAA7
FAA6
FAEF
FB33
FB06
FA91
FA64
FAAC
FAFA
FAEC
FAB0
FAA4
FAC1
FAB1
FA64
FA3C
FA84
FB06
FB5B
FB6A
FB62
FB4D
FB0A
FAB4
FAA5
FAFA
FB4D
FB3B
FAF8
FB06
FB62
FB83
FB37
FB12
FB92
FC2B
FBD7
FAC3
FAAD
FD11
013B
04C5
0604
057E
04E2
0502
055B
0549
04FB
04F8
0542
0566
053C
0519
0539
055D
0535
04E5
04D5
051F
0571
0582
0567
0553
0542
050F
04CA
04B3
04D3
04EE
04D3
04A7
04A6
04C9
04D2
04B1
049D
04B3
04C4
04A1
047C
04A2
04F4
04F1
0481
0449
04D0
0564
0475
014B
FD2D
FA54
F9CD
FAA9
FB4C
FB27
FAD7
FAE6
FB18
FAF9
FAA4
FA8B
FAC2
FAEB
FACD
FAA5
FABC
FAFA
FB12
FAFF
FAF8
FB05
FAF1
FAB3
FA97
FAD1
FB22
FB34
FB16
FB25
FB71
FB9F
FB75
FB2E
FB25
FB48
FB49
FB2B
FB43
FB94
FBAC
FB5A
FB27
FB99
FC3C
FBFE
FAC2
FA13
FBAF
FF7D
036F
0581
0589
04E2
04AD
04E1
04F7
04D6
04D8
051F
0568
0573
0552
053D
0533
0511
04D6
04B3
04B8
04BF
04AC
04A6
04DF
0538
055B
052C
04F4
0500
0531
0529
04D1
047F
047D
04A2
049B
046E
0463
0489
04A0
0496
04B3
0512
0536
04B1
0402
0439
055E
05C9
03BB
FF92
FBBD
FA41
FAC1
FB65
FB2A
FAA6
FAB5
FB2F
FB56
FB06
FAD1
FB10
FB64
FB5C
FB1E
FB13
FB38
FB36
FAF7
FACC
FADE
FAEC
FABA
FA7B
FA90
FAFA
FB4D
FB43
FB0C
FAFE
FB24
FB4B
FB5C
FB6B
FB7A
FB65
FB30
FB11
FB29
FB43
FB20
FAE4
FAF6
FB62
FB8C
FAF3
FA27
FAA8
FD60
016B
04A9
05BA
052A
0495
04D5
0565
056A
04E9
049A
04D0
0514
04E6
0474
0448
0489
04E6
0516
0527
0535
052B
04F6
04C5
04DB
0526
0549
0518
04CB
04A7
04A8
04AD
04B9
04D6
04DE
04AF
0471
0475
04BD
04EB
04D0
04B4
04E4
051A
04D8
044E
0459
053F
05D4
047F
0115
FD48
FB02
FAA4
FB0A
FB11
FAAF
FA84
FADA
FB59
FB92
FB74
FB37
FB0F
FB0E
FB29
FB3D
FB26
FAE6
FAB5
FAC8
FB15
FB58
FB5B
FB24
FAE2
FAAF
FA93
FAA1
FAEF
FB66
FBB8
FBA8
FB5C
FB2E
FB3C
FB46
FB14
FAD2
FADB
FB2C
FB56
FB24
FB00
FB56
FBC2
FB6C
FA65
FA31
FC57
0071
0438
05BE
0546
049B
04D9
057C
0586
04EB
0468
0460
0486
048B
049A
04E8
053A
0534
04E6
04B6
04C1
04BC
047F
045C
049F
0508
051B
04CE
048B
048D
049E
0487
047C
04BD
0518
0512
04A7
045F
0492
04E9
04E3
04A1
04A9
04FC
04EE
042E
038A
0405
053F
0557
02DF
FEA4
FB1F
FA02
FAB2
FB5E
FB18
FA83
FA85
FB0F
FB61
FB2B
FAE1
FAF7
FB3C
FB3D
FAEF
FAB3
FAB8
FACB
FAC5
FACF
FB0D
FB49
FB39
FAFD
FAF7
FB3B
FB73
FB5F
FB30
FB35
FB5C
FB5A
FB30
FB29
FB4D
FB48
FAFD
FADE
FB4C
FBE4
FBED
FB6B
FB37
FBC2
FC48
FBD6
FAEE
FB6C
FE62
028E
0573
05E5
04F9
0471
04D2
054A
0525
04A8
0482
04D6
052D
0531
050C
0508
0528
053E
053B
0533
052A
050D
04E5
04DD
0505
0526
0506
04B9
0493
04B8
04F2
04FC
04DB
04BE
04AD
0492
047A
0492
04C9
04C4
045B
03FD
042B
04B4
04DE
0468
0407
0463
04CF
03AF
006C
FC7F
FA1E
FA01
FAE3
FB3B
FAD0
FA7D
FAC7
FB45
FB5E
FB1D
FAF8
FB1F
FB53
FB5C
FB44
FB24
FAF3
FAB3
FA91
FAB3
FAFA
FB25
FB24
FB23
FB3D
FB49
FB1C
FACF
FAAE
FADD
FB37
FB88
FBB8
FBBC
FB87
FB30
FB04
FB42
FBBE
FBFC
FBC7
FB81
FB99
FBDC
FBA9
FAFF
FB01
FCF1
00A5
0452
062F
060D
0539
04E2
050E
051B
04CE
048A
049C
04D1
04D8
04C2
04D4
050F
0532
0520
0501
04F3
04E2
04BC
04A7
04D2
0517
0520
04D8
048C
0487
04B4
04D0
04CA
04C0
04BD
04A8
048A
0491
04C3
04D9
04A3
045A
045D
0494
047B
03F2
03A8
0447
0546
050A
0285
FE8F
FB42
FA08
FA77
FB23
FB35
FAEC
FAD1
FAE0
FAC8
FA90
FAA4
FB29
FBB0
FBB7
FB42
FAD1
FABA
FADF
FB04
FB26
FB5B
FB87
FB76
FB36
FB1C
FB55
FBA6
FBB7
FB85
FB47
FB20
FB00
FAEB
FB01
FB4B
FB94
FBAB
FBA8
FBB4
FBBC
FB93
FB62
FB98
FC27
FC50
FB8F
FAB3
FB6C
FE7C
029C
058B
0630
0569
04C4
04D8
051A
04FF
04BC
04CB
0528
0559
0520
04CE
04D4
052D
0567
052F
04B3
045F
0461
0490
04B9
04D3
04ED
04FF
04F1
04C1
0492
0481
0487
0489
047E
0473
046F
046E
0476
048B
0498
0484
0461
045B
0473
047A
046B
0496
0518
0531
03A6
0023
FC1C
F9BC
F9D6
FB2C
FBED
FB8E
FAEF
FAE4
FB41
FB57
FAFD
FAAA
FABD
FB05
FB1A
FAF1
FAD0
FAE5
FB12
FB22
FB08
FAE3
FADD
FB05
FB3E
FB51
FB2E
FB01
FB06
FB43
FB87
FBA4
FB9D
FB8E
FB80
FB6A
FB53
FB59
FB85
FBB1
FBA7
FB63
FB1B
FB0B
FB44
FB93
FBAF
FB87
FB6A
FBA0
FBE4
FBA2
FAE1
FAC1
FC90
0040
040F
060F
05F0
0504
049E
04D7
0508
04F1
04E5
0521
0562
0555
050D
04DD
04E9
050A
050D
04F4
04DA
04CF
04D3
04E2
04E7
04D1
04AD
04A6
04C5
04D9
04C4
04A8
04B0
04C4
04B2
0480
046D
0495
04C7
04C7
049C
0484
049D
04C4
04D0
04BB
0491
0464
045C
0491
04D2
04CC
049E
04CD
0560
054A
034A
FF87
FBD4
FA0C
FA47
FB11
FB32
FACD
FAA3
FAE1
FB12
FAFE
FAEB
FB15
FB4E
FB4E
FB20
FB09
FB24
FB4A
FB4D
FB30
FB16
FB13
FB20
FB2F
FB34
FB34
FB4D
FB95
FBE4
FBF3
FBBE
FB92
FBA3
FBC0
FBAC
FB7B
FB6F
FB89
FB89
FB55
FB21
FB1B
FB24
FB10
FB00
FB29
FB60
FB52
FB22
FB49
FBB4
FB9F
FADE
FAB7
FCBE
00BD
0484
0613
058F
04B8
04BC
053A
0561
0531
052D
0561
055B
04FD
04AD
04B6
04DE
04CD
048C
046A
048B
04C1
04D6
04C9
04BB
04BC
04C9
04DE
04EE
04EC
04E6
04F2
0502
04E3
049D
0478
0498
04BE
04AD
0487
048F
04B6
04B4
047D
0463
048F
04B9
04A0
0482
04BB
0502
04C2
0430
0446
0526
054A
030B
FEDD
FB2B
F9D6
FA6F
FB31
FB2B
FADF
FAF4
FB37
FB27
FAE2
FADB
FB15
FB2C
FB09
FAF9
FB2B
FB67
FB75
FB60
FB4A
FB2C
FAF5
FAC0
FABF
FAF2
FB20
FB31
FB3D
FB4F
FB40
FB0F
FAF6
FB18
FB41
FB46
FB4D
FB80
FBB1
FB9A
FB58
FB42
FB67
FB72
FB3E
FB1B
FB49
FB7E
FB5B
FB26
FB70
FBFA
FBCE
FAE1
FAD3
FD38
016F
04FC
061B
0569
04B6
04DF
0550
0556
0517
050C
0530
0531
050C
0503
0522
0535
052E
0523
050F
04DF
04B1
04BE
04FD
0520
04FF
04D3
04DF
04FF
04E1
0492
0479
04B6
04EB
04D9
04C0
04DE
04FF
04D9
0494
048C
04B8
04BF
0496
0494
04D5
04F5
04AD
045D
0478
04B4
0471
03EB
0420
0511
0507
0267
FDFA
FA6C
F981
FA74
FB51
FB3F
FAE2
FAF2
FB38
FB2B
FADC
FABE
FAE9
FB13
FB13
FB05
FAFC
FAF6
FAFD
FB16
FB20
FB02
FAE0
FAF8
FB35
FB3E
FAF6
FABA
FAE8
FB4F
FB71
FB42
FB39
FB84
FBB9
FB81
FB2F
FB33
FB70
FB7E
FB5E
FB63
FB90
FB90
FB50
FB3A
FB8A
FBD3
FBAA
FB6E
FBC3
FC50
FC07
FAFD
FB12
FDD5
0248
05A6
0655
0555
049A
04D1
0534
051F
04E5
0504
0552
055F
0530
051D
0533
052F
0504
04DC
04CD
04C4
04C3
04DB
04F8
04EC
04C1
04BA
04E6
04FE
04C4
047A
048C
04E8
0508
04C4
0491
04BF
04F4
04C4
0461
0445
046F
047D
045B
045C
049A
04B9
0487
0466
04A9
04DC
046A
03C3
0400
04FF
04DA
0215
FDC5
FAA5
FA21
FB1A
FBAB
FB50
FAE0
FAF4
FB30
FB15
FAD1
FAC7
FAE7
FAE5
FAD0
FAEE
FB34
FB5B
FB5A
FB64
FB83
FB8C
FB6E
FB4E
FB3A
FB12
FACA
FAA2
FAD4
FB2F
FB55
FB46
FB5D
FBA2
FBAE
FB5B
FB1C
FB50
FBAB
FBB6
FB87
FB85
FBB0
FBA9
FB6C
FB65
FBB9
FBE0
FB7D
FB1C
FB72
FC08
FBBD
FAC6
FB1F
FE32
02A6
059B
05D2
04BB
0450
04DC
0550
051D
04CF
04F1
0536
0525
04E3
04DA
04F6
04DF
04A7
04A7
04E4
0505
04ED
04D9
04F0
0503
04E4
04BA
04C3
04E6
04D6
0493
046F
0485
048D
0469
0460
049E
04D5
04B5
0472
0465
047F
0478
045E
0478
04B7
04B4
0461
043F
0495
04D2
046A
03F0
046D
056C
04D6
017F
FD07
FA4D
FA46
FB56
FBA3
FB22
FAE3
FB3E
FB7D
FB32
FAD9
FAF6
FB44
FB44
FB17
FB22
FB52
FB47
FB08
FAF8
FB2B
FB4F
FB3A
FB2B
FB4F
FB71
FB4E
FB0B
FB00
FB22
FB17
FAD6
FAC8
FB13
FB52
FB3E
FB26
FB63
FBB6
FBB7
FB79
FB63
FB7A
FB6F
FB3F
FB53
FBC4
FC11
FBE1
FBA6
FBE8
FC28
FB81
FA7F
FB2B
FE91
02F6
058B
0584
048F
0465
04F0
0525
04D3
04BA
052C
0587
054A
04DC
04D1
04FC
04E2
049D
04A9
050A
0542
051B
04E5
04E8
0505
04FE
04D5
04B5
049C
0477
045F
0489
04D7
04ED
04C0
04AC
04CF
04D1
0481
043F
045A
0489
046D
043D
046A
04D4
04E5
0488
045F
04BC
0500
0496
0423
04A8
058B
04AA
0113
FCB3
FA51
FA7D
FB63
FB6D
FADF
FABC
FB11
FB24
FACD
FAAC
FB09
FB56
FB2A
FAFB
FB48
FBB2
FB8D
FAFC
FABD
FB09
FB5A
FB41
FAF6
FAE1
FB06
FB27
FB37
FB57
FB7B
FB69
FB2B
FB13
FB37
FB4D
FB32
FB30
FB6D
FB96
FB68
FB2C
FB39
FB5E
FB3C
FAFC
FB19
FB86
FBAA
FB56
FB32
FBAC
FC05
FB58
FA76
FB86
FF48
03AE
05FD
05C3
04CE
04A5
0511
0536
04FD
04ED
051A
0515
04C6
04A0
04CD
04DC
048A
0453
04AB
0535
0548
04F1
04C4
04F4
0524
0514
04F1
04E8
04D6
049A
046B
0491
04DC
04E4
04B4
04C1
0516
052B
04C3
0466
048E
04E2
04D7
048E
048A
04C3
04BD
046A
0453
04AC
04DD
047A
0435
04DE
05A1
046B
0096
FC38
F9FA
FA36
FB1B
FB39
FAD7
FAD1
FB2A
FB45
FAFC
FAC0
FACD
FADA
FAC7
FAE4
FB54
FB9F
FB62
FAF5
FAEA
FB35
FB5C
FB3E
FB2A
FB45
FB57
FB39
FB13
FB0A
FB01
FADB
FAC9
FB01
FB4A
FB3A
FAE7
FAE0
FB43
FB7E
FB37
FAE9
FB1A
FB84
FB8F
FB44
FB30
FB6E
FB84
FB44
FB33
FB99
FBC8
FB22
FA96
FC0C
FFE1
03F6
05E3
058C
04C3
04D4
0563
0595
055D
0538
0544
0535
0501
04F5
051A
0513
04C3
0497
04D6
051C
04F5
049B
048F
04CE
04E5
04B7
04A4
04E3
052B
0525
04EB
04D1
04E2
04E6
04DF
0505
0543
052F
04B9
046F
04AF
051C
052A
04F3
04E8
0510
050B
04C2
048E
048B
045E
03EA
03D1
0483
04FD
037C
FFB9
FBC1
F9E8
FA59
FB55
FB7F
FB14
FAEE
FB2C
FB47
FB0A
FAD4
FAE9
FB14
FB0E
FAEF
FAF4
FB11
FB1F
FB27
FB3C
FB3B
FAFE
FAB9
FABB
FB03
FB38
FB28
FAFC
FAEC
FAFB
FB09
FB16
FB33
FB4B
FB35
FB06
FB0B
FB4C
FB73
FB47
FB02
FAF7
FB29
FB6A
FBA7
FBD5
FBC6
FB73
FB48
FBAC
FC40
FC16
FB15
FAAD
FC88
0064
040B
05A2
0575
0517
0540
055F
04F4
047E
04AA
0546
058B
053B
04E8
0505
054E
054F
051A
050A
0521
0512
04D5
04BE
04EE
0515
04E8
0494
047C
04B1
04E6
04E9
04DC
04EA
04FB
04EB
04D7
04F2
051C
04FC
048F
0444
0472
04D7
04E4
048B
046B
04FB
059A
04DB
0202
FE0C
FAF7
F9F8
FA81
FB20
FB12
FABE
FACE
FB34
FB5C
FB15
FACA
FADB
FB16
FB19
FAEB
FAE2
FB10
FB2D
FB0D
FAED
FB0D
FB49
FB4E
FB1E
FB12
FB4B
FB7A
FB58
FB13
FB05
FB2A
FB39
FB25
FB2F
FB70
FBA3
FB89
FB50
FB46
FB56
FB2E
FAE8
FB0A
FBA6
FBEF
FB45
FA7A
FB57
FE92
02B1
0561
05C9
0519
04D7
0538
056C
0510
04B4
04E8
056C
0599
0550
0500
04F4
04F6
04C9
049D
04BE
050C
0516
04B7
0457
0460
04B6
04F3
04F1
04E3
04E7
04D5
0495
0466
0492
04FC
053D
0522
04E1
04B7
049B
047D
0486
04D9
0529
04FD
0478
0463
050B
0560
03D6
003E
FC5E
FA50
FA6F
FB49
FB77
FB00
FAC4
FB11
FB59
FB20
FAAC
FA8C
FACE
FB09
FB08
FB02
FB2F
FB63
FB5A
FB22
FB07
FB27
FB56
FB6E
FB79
FB8B
FB8E
FB6A
FB3D
FB3A
FB5F
FB71
FB55
FB30
FB2B
FB31
FB23
FB1A
FB45
FB89
FB8E
FB4B
FB2F
FB89
FBE4
FB8A
FAB4
FAD3
FD25
011B
049B
05FF
0590
04DA
04DB
0540
0552
0504
04D4
04EE
0500
04D0
04A1
04C2
0513
0533
0509
04DB
04D3
04CA
04A4
0493
04C3
04FE
04E7
048A
0455
047F
04B8
04A1
0462
046B
04C5
0500
04DC
04AA
04C0
04E9
04B7
0449
0436
04A4
04F9
04BE
0475
04E4
059B
04F0
01E5
FDB2
FABE
FA32
FB02
FB7F
FB30
FAD2
FAED
FB22
FAF6
FA9E
FAA0
FAF8
FB2E
FB15
FB08
FB48
FB8F
FB81
FB41
FB3D
FB81
FBA1
FB64
FB1D
FB2D
FB70
FB75
FB30
FB0B
FB47
FB99
FB9D
FB5F
FB3A
FB4A
FB4A
FB17
FAF5
FB21
FB69
FB70
FB4B
FB68
FBC9
FBCC
FB16
FA83
FB9B
FED5
02C3
0545
059B
04E7
04AC
0530
05A2
0574
0504
04E8
0516
0521
04F5
04EA
051C
0531
04E2
047C
0475
04BC
04D2
048D
045B
0496
04F7
0509
04D7
04CE
0503
050D
04AF
0443
043F
048D
04B9
04AB
04B4
04F1
0506
04C5
0497
04DC
0536
0505
047E
048B
055B
0592
0399
FFA9
FBE6
FA3D
FA94
FB5E
FB84
FB31
FAF9
FAF2
FADF
FAC6
FAE3
FB30
FB59
FB3E
FB29
FB59
FB98
FB8B
FB3A
FB08
FB22
FB4B
FB45
FB29
FB33
FB59
FB58
FB22
FAFB
FB1A
FB5D
FB7B
FB6F
FB70
FB87
FB7D
FB38
FB00
FB24
FB74
FB78
FB25
FB02
FB65
FBC3
FB57
FA6E
FA9F
FD29
0150
04D3
0617
0597
04ED
04F1
0533
0518
04C7
04C5
0509
0516
04CF
04A9
04E9
052E
0504
04A0
0492
04EA
0522
04E9
04A0
04BB
050D
050D
04B0
047E
04B9
04F8
04C9
046B
0470
04D7
0510
04D8
049A
04BC
04F8
04CC
045B
0443
049F
04CD
0470
0432
04CD
0594
04BF
017C
FD3B
FA6A
FA02
FAE0
FB63
FB29
FAE5
FB06
FB33
FB04
FAB3
FAB5
FB0A
FB45
FB34
FB15
FB26
FB43
FB2E
FAF9
FAEC
FB17
FB3B
FB2E
FB1A
FB33
FB5E
FB5A
FB27
FB0C
FB28
FB47
FB2E
FB00
FB0A
FB5A
FBA7
FBBB
FBAC
FB97
FB68
FB16
FAEB
FB39
FBBA
FBB5
FB03
FAC3
FC69
0008
03E0
05F0
05D9
04F3
04A0
04FE
054A
0520
04DA
04DC
0504
04FC
04C7
04B7
04E8
051A
051C
0506
04FE
04F4
04CA
049F
04AB
04E2
04FA
04DD
04CC
04FE
0539
051B
04AD
0462
047B
04B4
04B8
049A
04A4
04D1
04DC
04C3
04D8
0528
0531
049F
040B
0464
0569
0562
02E2
FE9E
FAF6
F99E
FA26
FAEB
FB03
FACA
FAD3
FB07
FB03
FACD
FAC4
FAFC
FB29
FB20
FB14
FB2D
FB42
FB20
FAE8
FAE6
FB15
FB23
FAF7
FAE4
FB2B
FB8B
FB91
FB3D
FB02
FB29
FB70
FB77
FB48
FB30
FB41
FB40
FB19
FB15
FB62
FBAA
FB7F
FB0F
FB04
FB8B
FBE6
FB62
FAA0
FB4D
FE4C
026E
056C
0618
0551
04B9
04EB
054E
0545
0502
0500
053B
054B
0513
04E9
0502
0522
0508
04DD
04F1
0532
0543
050C
04E2
04FE
051E
04F1
04A4
04A3
04ED
0510
04D1
048D
04A7
04F3
04FA
04BC
04AC
04ED
0507
04A6
0436
044F
04C2
04CF
045C
0448
051B
05C3
0472
00C9
FCA0
FA3F
FA23
FAEA
FB32
FAEB
FACA
FB0D
FB47
FB2D
FAFF
FB09
FB28
FB12
FAD5
FAC3
FAEC
FB01
FAD3
FA99
FA9D
FAD4
FAFB
FB06
FB24
FB5A
FB62
FB1A
FAD0
FAE6
FB40
FB5F
FB14
FACA
FAEA
FB4B
FB72
FB50
FB50
FB97
FBBA
FB6C
FB19
FB57
FBE4
FBC6
FAD2
FA75
FC66
007A
0478
0642
05D7
04E1
04A0
04E5
04F3
04B5
04AA
04F5
052C
0504
04C3
04CC
050C
0528
050B
04F0
04F4
04F3
04DF
04E5
0518
0537
0504
04B8
04C7
0535
057A
0535
04B8
0498
04E5
052A
051B
04F8
0504
0511
04CD
0467
0469
04E0
0525
04BB
0426
044C
050B
04E1
0285
FE8D
FB1D
F9D1
FA5B
FB2E
FB4E
FB01
FAF3
FB33
FB4C
FB0C
FAC6
FACD
FB05
FB1F
FB0A
FAF3
FAF9
FB11
FB30
FB51
FB5A
FB29
FAD5
FABE
FB17
FB91
FBA6
FB45
FAE4
FADF
FB07
FB08
FAEF
FB0B
FB53
FB60
FB13
FAE4
FB38
FBC1
FBD6
FB72
FB40
FB8D
FBB5
FB1B
FA73
FB5C
FE84
0295
0567
060F
056F
04E5
04E7
0516
0521
0521
0537
054B
0545
0543
0559
0563
0535
04EB
04CD
04E3
04E8
04B5
0480
048D
04C7
04E4
04D4
04CD
04ED
0502
04E0
04AF
04B0
04D5
04CC
0488
0460
0499
04EF
04F1
04A7
048A
04CD
04FE
04B4
044F
049C
0590
05D7
0419
0082
FCCD
FAA1
FA2B
FA72
FAA4
FAB5
FADE
FB00
FADC
FA93
FA87
FACE
FB0A
FAED
FAAB
FAAA
FAF0
FB20
FB00
FAC4
FAB8
FADD
FAFF
FB0C
FB20
FB42
FB5A
FB5E
FB69
FB82
FB88
FB6C
FB62
FB95
FBC9
FB90
FAF8
FA9D
FAE8
FB6F
FB86
FB2D
FB14
FB7C
FBB0
FB0B
FA3E
FAE5
FDAF
015B
03F8
04E1
04FA
0538
0584
054E
04AC
0462
04D5
057C
059D
0530
04C5
04C1
0505
054B
057A
058F
0572
0523
04D8
04CC
04F6
0512
04FD
04D1
04A9
047B
0459
0483
0511
0596
0582
04DC
044C
045D
04CF
0500
04C9
049F
04C6
04DD
047F
041A
048E
05CE
0665
04C9
0124
FD69
FB72
FB4A
FB7F
FAFC
FA22
F9FC
FABF
FB8F
FB97
FAFB
FA7E
FA85
FAD3
FB0D
FB32
FB5B
FB5F
FB06
FA8B
FA75
FAEF
FB7C
FB8E
FB2D
FAD8
FADC
FB17
FB4A
FB70
FB8F
FB86
FB40
FAF8
FAFE
FB48
FB79
FB6D
FB5E
FB64
FB3D
FAD5
FAAD
FB3C
FBF6
FBB8
FA70
F9D0
FBB0
FFC9
03B5
0566
0518
0487
04B7
053A
0557
0523
051C
054D
055A
0533
0530
0565
055D
04D2
043C
0449
04F4
058B
058E
052E
04DE
04BF
04AD
04A3
04C3
0504
0524
0502
04C6
04A1
0491
0491
04BC
0509
050E
0478
03B7
03C9
050A
065B
05FC
034E
FF8D
FCA3
FB6D
FB45
FB21
FAB4
FA6B
FA9B
FB0D
FB52
FB41
FB07
FAD6
FAC3
FADC
FB2C
FB8E
FBA5
FB44
FABB
FA9D
FB0E
FB97
FBAC
FB4D
FAF0
FADE
FAEC
FADD
FACA
FAFA
FB60
FB95
FB5A
FAE9
FAB1
FAE4
FB6D
FC08
FC4C
FBCD
FAA3
F9CF
FA9F
FD67
00F3
0396
04B9
050F
0566
05AF
057C
04EF
04A6
04E3
0543
055F
0555
0565
0562
04F3
0448
040C
0489
052C
0546
04E5
04A7
04C8
04EC
04C9
04A3
04D7
0539
0540
04D0
046D
0490
0506
0545
0517
04BF
0481
0466
0475
04D4
0566
0585
0467
01ED
FEE5
FC69
FB08
FA9A
FAB0
FAF9
FB41
FB55
FB20
FACD
FAA0
FAAF
FAD0
FAD9
FADB
FAFF
FB43
FB6C
FB54
FB28
FB26
FB4E
FB61
FB40
FB18
FB18
FB2E
FB29
FB0F
FB1B
FB5C
FB7F
FB3E
FAD3
FABA
FB10
FB66
FB61
FB30
FB2D
FB42
FB1E
FAFB
FBCD
FE38
0194
0458
058A
0586
053E
0527
0516
04F1
04F0
053A
058A
058A
054A
051D
051C
0511
04E4
04CF
04F7
0524
050A
04C4
04AC
04D3
04E8
04B7
0481
0498
04DE
04F3
04CC
04C2
04FE
052E
050D
04DD
04FB
052E
04DA
0409
03AF
0470
055E
049A
016D
FD56
FA9D
FA1A
FABE
FB22
FAF4
FABB
FAC2
FAC5
FA96
FA7C
FABA
FB13
FB1B
FADB
FAC7
FB15
FB6E
FB68
FB0A
FAB6
FAB1
FAE9
FB30
FB6F
FB90
FB7C
FB41
FB1E
FB39
FB6B
FB7A
FB6C
FB6D
FB6D
FB2F
FACB
FAD3
FB91
FC4D
FBED
FA86
F9DA
FBC0
FFF8
041E
05F7
0585
04A1
04B7
0578
05C2
0542
04BA
04D5
0555
058E
055A
051E
051D
0519
04D8
0494
04B7
0534
0587
0555
04DB
0499
04B7
04EB
04E9
04BA
049D
04AE
04C8
04BA
0480
045B
0493
0517
0559
04DA
03EE
03B8
04E5
0678
0647
0330
FE99
FB4A
FAAC
FB8B
FBCB
FADB
F9F5
FA3B
FB3F
FBB9
FB36
FA77
FA4B
FAA1
FAEA
FB02
FB35
FB90
FBAD
FB45
FAA9
FA72
FACF
FB5A
FB8B
FB4B
FAF4
FAE9
FB37
FB97
FBC1
FBB0
FB95
FB8C
FB67
FAFD
FA9B
FAD4
FBB5
FC5A
FBD1
FA68
F9C4
FB56
FEC0
0217
03CC
0412
0440
050C
05D7
05AC
049E
03C7
040E
0527
05F9
05D9
052D
04C1
04CC
04DD
04A1
046D
04BA
0562
05A9
052A
0467
0434
04AD
051D
04F4
0478
0449
0484
04BB
04B1
04B4
0508
0556
04FD
0406
0359
03D3
0536
063C
05B3
0380
009C
FE31
FCB9
FBD3
FAF3
FA28
FA0C
FAE9
FC14
FC72
FBA3
FA7E
FA1F
FAAD
FB4D
FB4E
FAF3
FAE1
FB29
FB47
FAFE
FAC4
FB16
FBB8
FBF5
FB85
FAE6
FAB5
FAF9
FB4F
FB80
FBA9
FBD1
FBBD
FB51
FAE6
FB03
FBB3
FC53
FC2A
FB2D
FA22
FA06
FB3F
FD5F
FF9A
0172
02FD
047B
05C6
064C
05BA
048E
03D3
041E
0504
059E
057F
0504
04BB
04BB
04C1
04B2
04BF
04FB
0523
04F3
049B
048A
04E2
0543
0548
04FD
04B5
0491
0471
0454
047D
0503
0573
0532
0454
03AF
0402
050D
05D6
05B1
04D3
03D2
02D0
0155
FEFF
FC33
F9FF
F94C
FA22
FB92
FC68
FC11
FB02
FA35
FA37
FAC1
FB37
FB54
FB43
FB2E
FB00
FABA
FAA9
FB0F
FBA0
FBBF
FB44
FAC0
FAC6
FB31
FB6A
FB46
FB31
FB72
FBA2
FB3B
FA7E
FA50
FB13
FC07
FC21
FB4D
FA84
FA96
FB49
FBCD
FBEE
FC85
FE95
0208
056D
0715
067E
04C6
03A6
03EB
04E8
0567
0506
0475
0474
04EC
053A
0524
050D
053E
0561
0504
0464
043D
04C9
055E
0543
04A7
045B
04B9
0539
0533
04BB
0470
049B
04DD
04C9
0483
0482
04E0
052F
0506
048B
0443
0464
0456
0316
0037
FC9B
FA02
F99C
FAE8
FC29
FC16
FB07
FA54
FAB1
FB73
FB9D
FB28
FAE2
FB3E
FBC1
FBBB
FB3E
FAF6
FB2D
FB74
FB50
FAE9
FAC7
FB0C
FB54
FB58
FB42
FB59
FB81
FB69
FB0F
FAD5
FAFD
FB45
FB47
FB09
FB03
FB77
FBFD
FBEB
FB25
FA81
FB35
FDC3
0163
0476
05C4
0569
0499
0478
0519
05AC
0585
04DF
047A
04B4
0528
053F
04E3
0481
0473
04AB
04E6
050B
052A
053E
0520
04D5
04A8
04D3
0528
053C
04EF
0492
047A
0490
048A
0474
04AA
0539
0582
04F1
03F3
03C6
04FF
0684
0663
03D0
000D
FD25
FBF8
FBBB
FB42
FA62
F9DB
FA3A
FB28
FBD8
FBD1
FB40
FAAA
FA7B
FAC6
FB46
FB8E
FB61
FAEF
FAA3
FABB
FB10
FB5C
FB7C
FB6C
FB22
FAB2
FA6E
FAB0
FB5B
FBD9
FBC0
FB52
FB1B
FB2B
FB18
FAD8
FB01
FBD8
FC7E
FBBF
F9DA
F8D1
FA60
FDF2
0130
02A1
0317
042F
05FC
06FC
062A
0468
037D
0411
053D
05DA
05B1
0544
04F2
04BC
04A0
04B3
04F0
0528
0544
0553
0551
051E
04CB
04B6
0511
0575
0547
0495
0420
0469
050E
055D
053C
0511
04EE
0476
03C7
03CA
0511
0695
066E
0406
00ED
FF0B
FE60
FD54
FB26
F925
F915
FADB
FC79
FC5C
FAF9
F9F5
FA26
FAFD
FB8D
FB93
FB62
FB35
FB0C
FAE7
FADF
FAF6
FB10
FB23
FB3B
FB3C
FAF2
FA6F
FA2E
FA8E
FB49
FBAD
FB72
FAFC
FACB
FAE6
FB10
FB49
FBB2
FC03
FB9F
FA83
F9C3
FA90
FCD7
FF46
00DD
0209
03CD
060F
0762
06AD
04AA
0344
0391
04DA
05AA
0574
04DA
04A1
04D0
04F7
04E8
04DF
0509
0538
052D
04F1
04C5
04C4
04DA
04F7
0520
0545
0529
04BE
045D
0482
052F
05C7
05AC
04E1
0402
03A8
03FA
04BF
058E
05DF
052C
035B
00F4
FEB7
FCE9
FB4E
F9E3
F944
F9FA
FB82
FC76
FBFC
FAAF
F9EC
FA51
FB41
FBD0
FBB9
FB4E
FAD6
FA6B
FA41
FA95
FB36
FB8A
FB45
FADF
FAEF
FB58
FB6F
FB04
FAB7
FB0B
FB91
FB73
FAB8
FA55
FAE4
FBC8
FC02
FB87
FB26
FB4A
FB71
FB28
FB0A
FC32
FED6
01EB
0448
059D
062C
060E
0547
0455
0404
0494
055E
05A1
0555
04F6
04BB
0482
045F
04B1
0564
05B2
0515
042A
040E
04E4
0595
0548
0484
0466
04FC
0541
04B0
041A
046F
0544
055F
0482
03DB
0459
0551
0564
0474
03D1
0457
050F
043C
0162
FDC3
FAFF
F9C2
F9C7
FA80
FB5A
FBBB
FB60
FABC
FA8F
FAFE
FB6C
FB59
FB13
FB20
FB61
FB44
FABE
FA88
FB12
FBC1
FBAD
FAF0
FA93
FB22
FBE9
FBEE
FB4E
FB03
FB72
FBE1
FB9A
FB08
FB22
FBEC
FC44
FB66
FA34
FA77
FCEB
0077
0360
04DF
0560
0589
0588
054A
04F3
04C9
04D9
04F3
04FD
0511
0537
0546
0523
04F9
04FC
050A
04D9
0478
0459
04B4
0527
0528
04BF
0471
047D
0488
0441
03FB
0441
04E6
050C
0453
038E
03D9
051C
05E7
04E7
0233
FEFE
FC59
FA9A
F9C4
F9E2
FAC0
FB9E
FBB1
FAF7
FA39
FA28
FAAB
FB1D
FB1B
FACE
FA93
FA98
FADA
FB42
FBA2
FBB3
FB61
FAFD
FAF9
FB5E
FBB4
FB9A
FB40
FB1D
FB45
FB57
FB23
FB0C
FB7D
FC1C
FC03
FAEF
F9DE
FA40
FC73
FF75
01FC
03A3
04CC
05B1
060A
05A1
04E5
0490
04E9
0586
05D7
05B3
0550
04F0
04B3
04A7
04C6
04E6
04DA
04A9
048A
04A1
04D0
04E8
04E0
04CD
04AD
0466
0413
0411
0499
0547
0560
04A8
03D4
03DE
04E6
05DA
0568
033A
0039
FD91
FBBE
FA91
F9E9
F9F3
FAAD
FB7C
FBA5
FB14
FA7C
FA86
FB0D
FB66
FB31
FAC1
FA97
FACE
FB16
FB2E
FB21
FB1E
FB37
FB52
FB4A
FB1E
FAFF
FB2E
FBA1
FBE7
FB93
FADB
FA93
FB3F
FC41
FC5D
FB2A
F9C9
F9CD
FB9D
FE37
007C
0248
040F
05BD
067F
05D0
045F
0392
0425
0578
0641
05D7
04C5
0427
0489
0565
05BF
053B
0472
043C
04B3
052F
0528
04DC
04DA
0524
0524
0497
0414
045A
053F
05C2
0538
042C
03BC
0456
0546
058E
04D7
036C
0195
FF54
FCC5
FA88
F977
F9E9
FB43
FC4D
FC23
FAF8
F9F6
FA26
FB5A
FC44
FBDA
FA91
F9E4
FA95
FBC2
FC00
FB1F
FA54
FA95
FB5F
FB8B
FAF3
FA9C
FB2F
FBF6
FBD7
FAE7
FA57
FAD9
FBBD
FBEC
FB55
FADA
FB02
FB67
FB94
FBFA
FD8C
0083
03E5
0646
06D9
05DE
0469
03B6
0453
059B
0640
059D
0483
0448
051F
05CD
0545
0413
03AE
048C
0596
059F
04DD
046C
04B8
050A
04C0
044A
047B
0539
058A
04EE
0419
0406
04B4
053A
0512
04B1
04B5
04D1
03EA
015B
FDCE
FAC8
F97D
F9FA
FB3E
FBF9
FB7A
FA42
F995
FA3C
FB9F
FC54
FBB2
FA95
FA59
FB2E
FBED
FB9E
FAB8
FA68
FAFA
FB85
FB47
FAB6
FABF
FB63
FBB6
FB3E
FAB5
FAF6
FBB0
FBC9
FAFA
FA4F
FAB5
FB9C
FBB6
FAE6
FABA
FCB0
0064
03E6
05A1
0597
04D2
043E
0430
04A0
0542
0593
0547
04BD
04B0
053F
05A7
0539
0459
0414
04B7
0562
053D
0496
0464
04DA
0529
04C0
042D
044C
04FE
054F
04E9
049E
052D
0602
05E2
04B1
03CF
0454
0570
0521
0272
FE8F
FB8C
FA6E
FAAA
FB27
FB49
FB10
FABB
FA8E
FAB6
FB18
FB53
FB23
FAC4
FAB3
FB08
FB53
FB34
FAE7
FAEF
FB56
FB9C
FB6A
FB09
FAF8
FB32
FB44
FAFF
FAC5
FAE9
FB24
FAEF
FA64
FA48
FB01
FBDD
FBC5
FABB
FA2C
FB93
FEE3
0284
04DB
0592
056A
0529
0503
04E8
04E8
0514
053E
0527
04DD
04B8
04E7
052B
052B
04E4
04A1
0490
049D
04B2
04DD
0520
0542
0517
04CE
04CA
0511
0534
04EC
0494
04B3
052A
0542
04B5
043C
04AF
05AA
059A
0367
FFC1
FC7F
FAD2
FA6D
FA6A
FA7A
FAD6
FB62
FB85
FAF6
FA48
FA53
FB22
FBE8
FBF4
FB6B
FAF4
FAE1
FAFA
FAF3
FAD4
FACC
FAE3
FAF8
FAF3
FAE1
FAD7
FAE0
FB02
FB35
FB59
FB48
FB16
FB10
FB61
FBB5
FB82
FAC0
FA39
FB03
FD7F
00ED
03EE
0592
05DD
0576
04FF
04BD
04B9
04F2
0548
0567
0506
0457
0402
0478
0554
05AF
052E
0475
0463
0500
057D
053F
0499
0452
04A7
0517
0524
04E3
04B3
04B4
04C1
04C4
04D0
04EA
0500
0518
053C
051F
0416
01B8
FE8F
FBCA
FA48
F9FF
FA67
FB12
FBB2
FBDF
FB5B
FA94
FA63
FB07
FBB0
FB6A
FA65
F9D9
FA88
FBC5
FC49
FBBD
FAFA
FAD1
FB1B
FB30
FAEF
FACD
FB0B
FB54
FB4A
FB19
FB21
FB54
FB50
FB0A
FAE9
FB15
FB22
FAC8
FAB8
FC24
FF42
02C2
0504
0596
0541
04D4
047D
043F
0469
051E
05C8
059F
04CD
045F
04ED
05B5
0592
0492
03E9
0461
0559
05B1
0537
04BE
04D4
051B
0501
04A4
048D
04D1
04F8
04CE
04B5
04F6
0531
04E0
0448
0443
04FC
0540
0398
0006
FC44
FA28
FA0F
FAE5
FB77
FB62
FAEB
FA72
FA44
FA9A
FB5C
FBEC
FBA8
FAB6
FA11
FA71
FB59
FBA9
FB11
FA6F
FAA1
FB5E
FBAB
FB30
FA97
FA89
FADD
FB0D
FB13
FB43
FB83
FB4D
FAAB
FA7A
FB36
FC0B
FBCE
FACE
FAEA
FD75
0181
04C0
05E6
05A0
053C
0520
04F4
04A6
0494
04D3
04FD
04E2
04EA
0567
05E7
05AE
04CD
0436
048F
0558
0595
0517
04A0
04C4
052C
0532
04D1
049F
04E7
0545
0542
04FE
04E4
04E9
049B
03FE
03DA
04AD
058D
04B5
0174
FD3B
FA64
F9FC
FB07
FBD6
FBB2
FB14
FAA0
FA7F
FA97
FADC
FB2A
FB28
FABD
FA60
FAA1
FB5C
FBC0
FB52
FA90
FA4E
FAB3
FB20
FB1C
FAEE
FB0F
FB69
FB7E
FB29
FAD7
FAE1
FB19
FB26
FB1C
FB56
FBCC
FBEF
FB7F
FB43
FC7E
FF7E
0300
0548
05BB
053E
0506
0557
0593
053E
049E
044D
0485
0502
056C
0599
0575
0509
04A9
04BF
0541
0599
0552
04B6
046B
0491
04A6
0463
043D
04BA
0581
05B5
052A
04A9
04BB
04D6
0449
0385
03B1
04DD
0556
035F
FF4E
FB6F
F9BC
FA24
FB1F
FB7A
FB2A
FABD
FA91
FAA5
FAC7
FAC4
FA8F
FA56
FA60
FAB6
FB0D
FB1F
FB09
FB28
FB94
FBF0
FBD5
FB60
FB0C
FB1F
FB5F
FB62
FB14
FACE
FAEC
FB57
FB9B
FB79
FB3E
FB5E
FBBF
FBD9
FB9F
FBFE
FE00
015D
0462
058F
0521
04A2
050F
05DE
0606
0571
04F2
0516
0585
05A4
0566
052B
051F
050D
04CE
0494
049B
04C9
04D8
04BA
04A0
04A3
04A2
0487
0471
048B
04CA
04F4
04ED
04C6
0498
045F
0423
041B
0468
048E
038F
00E7
FD69
FAC5
F9F9
FA71
FADB
FAA9
FA6C
FAB6
FB27
FB02
FA5D
FA1D
FAB7
FB82
FB9F
FB23
FADB
FB1F
FB73
FB5A
FB0D
FB10
FB5A
FB6F
FB27
FAEB
FB07
FB3D
FB38
FB1E
FB47
FB93
FB92
FB3A
FB0B
FB4A
FB9A
FB97
FBC2
FD31
0041
03C6
0600
0646
058A
0527
0583
05ED
05B4
0506
04A4
04DF
0533
0502
0479
044F
04BC
0523
04EE
0460
0431
0487
04CC
049E
0464
04AA
052B
0525
047B
03F7
0429
04A4
04C5
04B4
04F7
0534
0420
0118
FD3F
FA8C
F9D6
FA41
FA90
FA78
FA6E
FAA7
FAD9
FAD8
FADF
FB21
FB70
FB7D
FB47
FB16
FB23
FB59
FB82
FB93
FBAB
FBD2
FBDC
FBA1
FB3D
FB0A
FB3F
FBAB
FBDD
FBAD
FB6B
FB65
FB62
FAFC
FA90
FB57
FE16
01F3
04F5
05DE
053E
0497
04BF
054D
0584
0546
0502
04FB
0508
04F2
04C6
04AC
04AF
04B5
04A5
048C
048E
04B0
04C8
04B1
0485
0485
04BA
04DD
04BB
0483
0484
04AC
0498
0442
043F
04D6
0519
0382
FFD3
FBD3
F9B4
F9EA
FB02
FB74
FB19
FABF
FAD9
FB17
FB1B
FB02
FB0D
FB2C
FB26
FB0C
FB25
FB7C
FBC4
FBC7
FBA0
FB8C
FB92
FB7D
FB2D
FACF
FAB8
FB03
FB63
FB86
FB7B
FB92
FBC7
FB9B
FAD8
FA63
FBC5
FF79
03D5
065D
0635
04E5
046C
051D
05C3
0586
04E4
04C8
053F
0591
0550
04D1
0492
049B
04B4
04CD
04EF
04F1
04A1
0430
0416
047E
0505
052D
04EC
04AE
04CE
051D
051C
04A9
044C
0495
0529
04B2
022A
FE35
FAE6
F9D5
FA93
FB4F
FAFF
FA47
FA3F
FAE4
FB4C
FB08
FAA4
FAB7
FB0C
FB15
FAD3
FACF
FB42
FBB3
FBAA
FB50
FB21
FB34
FB3F
FB2D
FB3F
FB90
FBC2
FB75
FADD
FAA4
FB17
FBA8
FB85
FACB
FAD2
FCF1
00DE
0490
060B
054D
0424
042D
0531
05D4
057A
04EB
0502
0583
0599
051E
04B6
04CA
04FE
04DF
0498
049B
04D9
04D2
0474
0455
04CF
0551
0515
0441
03D4
0458
052D
0561
04F8
04D5
055C
058C
03E9
004C
FC73
FA6A
FA97
FB8D
FBC7
FB29
FAAA
FAE0
FB54
FB58
FAFF
FADF
FB1A
FB36
FAF4
FAB8
FAE1
FB25
FB0D
FABF
FAD1
FB54
FBA3
FB57
FAF8
FB47
FC0A
FC36
FB68
FA8D
FAB6
FB9A
FBE4
FAFE
FA0B
FAD4
FDE7
01EE
04D8
05A1
04FE
0468
04A0
0533
0547
04B6
0429
0437
04AD
04EA
04C3
04A3
04D4
0515
0517
04F8
0505
0531
0533
050B
04FD
050E
04EC
0478
0425
0461
04DA
04D4
0450
0437
0513
05F4
053B
0260
FE9F
FBCE
FAC7
FB09
FB81
FB89
FB2D
FAD9
FAD6
FB0D
FB2D
FB11
FAEF
FB19
FB88
FBDE
FBD9
FB95
FB47
FAF0
FA8C
FA4E
FA70
FAD3
FB1E
FB34
FB4C
FB86
FBA3
FB67
FB0D
FB00
FB2E
FB09
FA85
FAAF
FCBB
0083
0442
061B
05C4
0499
0423
04B0
0560
0565
04E9
04A4
04DD
051F
04F4
048D
0479
04DF
0543
0532
04D6
04AF
04D9
0500
04FA
0500
0530
053E
04ED
048C
048A
04CA
04D2
04A3
04D9
05A5
05F7
0454
00A1
FCA0
FA5A
FA3B
FB07
FB60
FAFE
FA83
FA86
FAF8
FB56
FB3C
FAD5
FA99
FABD
FAFB
FAF1
FAA9
FA8D
FADB
FB4C
FB76
FB52
FB2A
FB18
FAF4
FAC8
FADF
FB36
FB5C
FB1B
FAE7
FB32
FB89
FB26
FA5E
FADE
FDCE
0211
051B
0597
04AA
044B
04F3
0597
056E
04EE
04F0
0573
05BE
0567
04D5
04A6
04EE
0541
054D
052A
0520
0541
0564
0557
050D
04AF
0473
0472
04A0
04E0
050D
04FD
04B9
049E
0508
059C
0537
02EF
FF3E
FBE0
FA54
FA92
FB51
FB77
FB05
FA9D
FA94
FAB6
FAC2
FABE
FAD0
FAFA
FB1B
FB1A
FAFC
FADA
FAC4
FAB9
FABA
FAD1
FAF9
FB07
FADF
FAB6
FAE7
FB72
FBD1
FB8B
FAEB
FABF
FB39
FB82
FAED
FA60
FBB4
FF66
038E
05C0
0593
04B3
04A9
0547
0585
0520
04CD
04FA
053D
051D
04D4
04E1
053A
056A
0545
04FD
04C3
04A3
04B8
0514
0579
0573
04ED
046E
0483
0511
0571
053E
04B9
0469
0490
0507
053D
044C
019D
FDE8
FB0C
FA54
FB1C
FB99
FAF5
FA12
FA16
FAE6
FB7C
FB6B
FB3F
FB53
FB31
FA81
F9EC
FA54
FB78
FC29
FBCA
FB06
FABE
FAE6
FAD7
FA72
FA51
FAC6
FB46
FB2B
FAB1
FAA2
FB27
FB7C
FB0C
FA76
FB20
FDBE
0173
047C
05B4
0565
04B1
0468
0489
04B8
04D8
050B
054B
055B
0516
04B7
049A
04CA
04F6
04DF
04AB
04B2
0508
056B
058D
0565
051F
04ED
04E7
050E
054E
0579
0554
04D4
0464
049C
056A
059F
03D4
000E
FC27
FA34
FA83
FB81
FBA7
FB0B
FABE
FB1A
FB69
FB2D
FAE3
FB1A
FB73
FB3C
FA9F
FA7F
FB29
FBCF
FBA8
FB01
FABB
FB02
FB2B
FAD9
FA88
FAAB
FAEE
FAD0
FA91
FAD2
FB7A
FBA7
FAE4
F9F6
FA3A
FC52
FFA2
02DF
04EE
0570
04E2
0450
047E
0533
0590
053D
04D1
04E1
052A
051A
04C7
04C4
0521
053C
04BA
0428
043B
04C0
04EB
048F
045C
04BD
052A
0513
04D6
051F
05B0
0599
04BE
0441
0501
0609
0552
0218
FDE0
FAF7
FA3D
FAC3
FB32
FB16
FAC4
FAA1
FABB
FAE9
FB0F
FB2F
FB50
FB64
FB54
FB23
FAF9
FB05
FB4A
FB92
FBA6
FB84
FB5A
FB4E
FB58
FB58
FB3B
FB05
FAD0
FAD2
FB33
FBB5
FBC0
FB05
FA28
FA84
FCF3
00CD
043C
05C6
057E
04B5
0489
04EE
0523
04D4
046E
0475
04D1
050B
04FB
04EA
0506
0506
04A5
042F
0432
04B1
0514
04FE
04C5
04CF
04E5
049A
041E
042D
04EC
0586
0538
0480
048C
057B
05CB
03F9
004D
FCAC
FAB9
FA8D
FB1C
FB6B
FB3D
FAF0
FAEA
FB37
FB86
FB81
FB33
FAFE
FB27
FB73
FB71
FB1E
FAE7
FB0B
FB47
FB53
FB50
FB7C
FBB4
FBA8
FB5A
FB17
FAF8
FAD0
FAA8
FADF
FB7D
FBC4
FB0F
FA21
FAD3
FE05
024C
0536
05B1
04CD
0430
0471
0500
0534
0503
04BE
049D
049F
04B9
04DF
04F6
04F8
04FD
0513
051B
04F0
04A5
0474
047F
04BB
04FD
0516
04F3
04C2
04C4
04EB
04DA
0470
0437
04D0
05D6
05BB
0343
FF21
FB98
FA51
FADC
FB9B
FBA3
FB50
FB3B
FB57
FB3D
FADC
FA8D
FA8D
FABA
FAE1
FB05
FB3B
FB69
FB61
FB28
FAED
FAD5
FADD
FAF9
FB1C
FB3E
FB63
FB83
FB7F
FB40
FAF3
FAE8
FB18
FB14
FAB3
FABF
FC6E
FFE6
0398
058B
0556
0462
0432
04D6
055A
053E
04EA
04DF
0511
0533
0541
055D
0567
051D
04A5
0486
04F2
0568
0552
04CF
048B
04D6
053B
052D
04C4
0492
04DA
0531
0512
0495
045B
049E
04A8
0375
00D5
FDC3
FB80
FA85
FA66
FA8F
FAC9
FB1B
FB64
FB65
FB21
FAE6
FAEA
FB0C
FB1A
FB11
FB08
FAF7
FAD2
FAB5
FAD0
FB24
FB75
FB89
FB5F
FB24
FB04
FB06
FB0B
FAFC
FAE5
FAF4
FB38
FB6A
FB34
FAE2
FB97
FE35
020B
051F
0619
0586
04EA
04F0
051A
04F1
04BF
04E7
051A
04D3
045A
0482
055A
05EC
058F
04D6
04A7
04EE
04F2
0494
047A
04F4
056D
0542
04B2
0474
04AF
04EF
0504
0529
0514
03C2
00BD
FD26
FAB8
FA0A
FA4F
FAA8
FAEF
FB3C
FB4E
FAEB
FA77
FA8D
FB19
FB64
FB21
FAD8
FB03
FB4F
FB36
FAE1
FADA
FB22
FB3A
FB02
FAEF
FB46
FB96
FB6A
FB11
FB20
FB68
FB2F
FA9D
FB22
FDD1
01BA
04AE
058A
051D
04C8
04E8
04FC
04CE
04C7
0521
0571
0551
0505
0510
056A
0587
052E
04C9
04BF
04F3
0504
04E4
04CE
04D4
04CB
04B1
04C2
0503
0518
04D4
049F
04D9
04F0
03A7
009A
FD14
FAEC
FAA4
FB23
FB39
FAE0
FAB9
FAF0
FB21
FB1C
FB1B
FB32
FB0D
FA88
FA1C
FA50
FAF0
FB45
FB13
FAD6
FAEB
FB0A
FAED
FADC
FB29
FB84
FB73
FB2B
FB48
FBAF
FB80
FAA5
FAB0
FD39
018B
04F3
05B3
04CC
044E
04CB
0551
054A
0535
057C
0597
0502
0451
0483
0581
0623
05D3
0541
052B
054A
050B
04AD
04CD
0547
055A
04E9
04A9
04F0
051E
04AC
043C
04A2
052E
0401
008A
FCAC
FAB5
FAD4
FB63
FB3D
FACB
FAD2
FB2E
FB49
FB1D
FB17
FB41
FB28
FAB6
FA72
FA9F
FAD1
FAA6
FA76
FAB7
FB24
FB23
FACC
FAC5
FB23
FB2E
FA9D
FA49
FB06
FC1F
FC0C
FACD
FA88
FD11
017A
04EA
05C4
0506
0495
04FC
056E
0554
04FC
04D2
04B4
0479
0478
0507
05BF
05DC
054A
04BB
04BA
0510
0546
055B
058B
05B0
056D
04DF
0498
04C3
04D5
0480
045F
050A
05B6
04A5
013A
FD17
FA8C
FA37
FAC4
FADB
FA92
FAA4
FB1C
FB5F
FB35
FB05
FB16
FB2F
FB17
FB00
FB23
FB40
FB04
FAA5
FAA8
FAFD
FB11
FACA
FAC7
FB4C
FBA4
FB32
FA91
FACC
FBA4
FBB5
FAAA
FA5A
FCC4
013E
04D9
05B1
04DD
048D
0544
05D2
057B
04DD
04BC
04EB
04E3
04BE
04F1
0555
0549
04BD
046A
04B9
052C
0537
0512
052A
0548
04F8
0481
0495
0526
054D
04AD
0432
04B6
0557
0421
009A
FCAF
FA9D
FA9B
FB2B
FB37
FAF6
FAF2
FB20
FB35
FB42
FB76
FB94
FB44
FAB8
FA8E
FAE0
FB16
FAD9
FA9E
FAE0
FB42
FB1C
FA9A
FA8C
FB2B
FBB1
FB8C
FB3D
FB87
FC08
FBA0
FA5F
FA28
FCAD
0125
04E0
0613
0575
04E8
0534
0598
0548
048E
043A
0488
04FC
0520
04FE
04D4
04BF
04BE
04D4
04F6
0508
0503
0505
0518
050B
04BC
0471
0488
04D9
04D5
046C
0464
0536
05E9
04B9
0129
FCF0
FA5C
FA0C
FAB5
FAFC
FAD6
FADD
FB1E
FB2C
FAF9
FAF1
FB35
FB62
FB39
FB0D
FB35
FB66
FB27
FAAC
FAA3
FB21
FB67
FB0C
FAAA
FAEF
FB8F
FBC5
FB8E
FB94
FBE8
FBB6
FACF
FAAA
FCF6
0139
04D8
05DE
04FC
0448
04A2
0534
051F
04AB
0495
04F4
0545
053C
0509
04E1
04C0
04A9
04BD
04EF
04F5
04C9
04C7
0512
0541
0502
04B3
04D1
050E
04AA
03C1
037C
0471
0556
0425
0095
FCBC
FACF
FAE5
FB6E
FB5E
FB0B
FB19
FB69
FB72
FB25
FAEF
FB02
FB20
FB21
FB36
FB78
FB96
FB4A
FAD8
FAB4
FAD8
FAD7
FA97
FA85
FAED
FB7D
FBB5
FBA3
FBAE
FBD4
FB95
FAFB
FB31
FD68
013B
04AA
0602
0577
049E
048D
04F9
0517
04C7
0490
04B7
04EE
04DB
0495
0472
048D
04B7
04CA
04CB
04CD
04D3
04E5
0504
0516
0506
04F9
051F
0547
0502
0468
044C
0516
05B2
044D
0083
FC4D
FA25
FA6E
FB57
FB46
FA93
FA7B
FB30
FBBB
FB7C
FAEB
FABF
FAF1
FB0C
FB02
FB22
FB71
FB93
FB77
FB7C
FBBE
FBC5
FB4B
FACA
FAD8
FB3B
FB44
FAE6
FABC
FAFA
FB0B
FAAE
FAF2
FD34
0125
04A5
05F0
0567
04B4
04BD
0511
0515
04E3
04D6
04EB
04E4
04D1
04EF
0529
051F
04C2
0479
048A
04BC
04CD
04D6
04FB
04FF
04A8
0446
0460
04DB
050D
04C7
04CA
0598
062D
04B8
00DB
FC87
FA21
FA1A
FAE3
FB0C
FAB3
FABB
FB52
FBC5
FB91
FB09
FACC
FB00
FB54
FB84
FB86
FB57
FAFD
FAAE
FAAE
FAF8
FB37
FB3B
FB34
FB59
FB84
FB71
FB3E
FB46
FB6F
FB2F
FA8A
FAAA
FCD9
00CA
0479
060E
05A1
04C9
04B0
0518
0547
052A
052B
0554
0545
04E0
0487
0486
04A7
049A
0480
04A6
04FA
0516
04E9
04D0
04FC
0522
050C
04F2
04FF
04E2
0464
040D
048A
0547
0482
014E
FD25
FA9E
FAA3
FBA8
FBCC
FAFD
FA62
FA77
FAAB
FA96
FA9C
FB1A
FB9C
FB7B
FAE3
FA9C
FAEF
FB5A
FB69
FB4D
FB4E
FB40
FAF8
FACB
FB0B
FB63
FB4C
FAF5
FB0B
FB8D
FB9E
FAF6
FAE8
FD0D
0102
0461
0560
04B0
0446
04E0
0591
0579
04E8
04A9
04DF
051A
0525
0530
0544
051E
04C0
0497
04DD
0533
0533
050C
0523
0557
0536
04C7
0489
04A4
04A7
0462
047D
0574
0638
04D0
00C1
FC35
F9F3
FA7E
FBD9
FC0B
FB26
FA89
FAD3
FB58
FB5C
FB0E
FB02
FB44
FB63
FB2E
FAE5
FABC
FAA9
FAA4
FAC2
FAF4
FAF1
FAA6
FA78
FACA
FB61
FBAB
FB8D
FB74
FB78
FB1E
FA66
FA8F
FCF8
012A
04CA
05EF
0516
044B
04A2
054F
0538
0492
0458
04CB
053C
052D
04E2
04CE
04EC
04FB
04FB
0512
0526
0507
04E2
050C
0561
0562
050E
0505
056F
0582
04B2
03D7
042C
0532
04AC
014C
FCB5
F9F1
FA18
FB65
FBC3
FB30
FAF8
FB88
FC01
FBBD
FB24
FAD9
FADB
FADA
FAE5
FB36
FB8B
FB62
FAD1
FA85
FAC4
FAFF
FAC2
FA72
FA9F
FB15
FB38
FB17
FB42
FBB4
FBA5
FAF4
FAFA
FD37
012E
048D
059E
0501
0475
04AD
04F7
04C3
046F
0489
04EB
050B
04D4
04AB
04D0
0513
053B
054F
054D
050E
04A0
0472
04C0
0526
0520
04D4
04CD
050E
04FE
0471
0437
04FA
05D2
04D1
014B
FCFE
FA6F
FA5C
FB56
FBBB
FB58
FAF8
FB0A
FB34
FB21
FAFE
FB0D
FB2F
FB24
FAFE
FAFD
FB27
FB48
FB52
FB65
FB7C
FB61
FB0F
FADA
FAFE
FB3C
FB36
FB0F
FB2B
FB66
FB22
FA6F
FAA8
FD14
011F
0483
0592
04DE
0440
049F
0540
0533
04A7
046D
04C2
051D
051D
04F3
04EA
04F4
04E2
04C6
04CF
04E6
04C9
0478
0446
046B
04C0
0512
0555
056E
0522
048E
0454
04D3
0548
0446
0150
FDA5
FB26
FA8C
FB08
FB77
FB80
FB60
FB3B
FB09
FAE0
FAE3
FAF5
FAE4
FAC9
FAF8
FB6E
FBC0
FBAA
FB76
FB84
FBA7
FB6A
FAE2
FAB6
FB25
FB88
FB43
FAB3
FAAC
FB29
FB4C
FAD8
FAFF
FD1F
00E3
043B
057B
04F4
0443
0465
04FC
0544
051D
04EF
04F5
0505
04ED
04BA
0499
048C
047F
0479
049B
04E7
0529
0537
051A
04FD
04E9
04BD
046F
0444
049B
0546
0549
0390
0023
FC77
FA50
FA34
FB20
FBB8
FB88
FB17
FAEE
FB01
FB08
FAFF
FB19
FB4D
FB55
FB28
FB13
FB4F
FB9B
FB8E
FB2E
FAEC
FB09
FB39
FB1D
FADE
FAF5
FB58
FB66
FADF
FABB
FC60
FFF1
03BF
05CB
05B3
04D5
0493
04F2
051A
04BD
046D
04A6
0514
0525
04E2
04D3
051D
0549
0507
04AF
04C0
0518
0522
04BB
0473
04B7
051C
04F3
0463
0455
0518
057E
03EF
0053
FC89
FAA0
FAD9
FBA5
FB8E
FAB9
FA52
FAD9
FB8C
FB7E
FAC9
FA53
FA99
FB2F
FB7B
FB80
FB9B
FBC1
FB85
FADB
FA5F
FA94
FB29
FB73
FB5E
FB64
FBA6
FB93
FAE1
FA88
FC02
FF80
0348
054E
0538
046E
0452
04E5
054F
052E
04F8
0521
0573
0571
0519
04E2
04FD
0508
04A4
041B
0410
04A0
052B
0523
04C1
04A3
04E1
04F2
049A
046D
04EB
054F
0405
0096
FCAB
FA86
FAAB
FB8A
FB86
FAC2
FA83
FB36
FBE1
FB93
FAAA
FA3B
FA9A
FB14
FB19
FAF4
FB2E
FBA4
FBBC
FB52
FAF6
FB19
FB6E
FB70
FB36
FB46
FBA5
FBA3
FAF1
FA85
FBE1
FF4D
0330
0581
05B8
050E
04E5
0556
0583
0501
0461
0457
04D0
0531
0537
052E
0549
0540
04CC
0444
044C
04E8
055D
051B
047E
0446
048A
04AA
045B
0434
04C3
055D
046F
014E
FD49
FA8E
FA05
FAB1
FB16
FADB
FAB1
FB07
FB65
FB39
FAB8
FA96
FB00
FB61
FB3F
FAE5
FAE9
FB46
FB6D
FB29
FAF7
FB44
FBBC
FBBD
FB55
FB35
FB95
FBBB
FB12
FA6F
FB87
FEE3
02EC
055E
0591
04D2
04A4
052A
0589
054C
04E4
04D9
050D
051A
04F7
04F0
050E
0500
04AA
046F
04A9
0513
0516
0496
0429
044F
04BE
04CC
0473
0472
0530
05C5
04A3
0154
FD4B
FAAB
FA4B
FB1C
FB8E
FB2E
FAB5
FAC7
FB22
FB2C
FADB
FAB1
FAE7
FB23
FB0F
FAED
FB2E
FBB0
FBD2
FB58
FAD6
FAE8
FB61
FB97
FB5F
FB41
FB84
FB9C
FAFF
FA60
FB54
FE7F
027F
0526
059F
04F8
04A2
04E9
0524
04F5
04BB
04D9
051E
0527
0501
0505
0530
0517
049D
0444
047C
04F6
04FB
0476
0423
0488
0522
0509
0447
03FB
04DC
05EA
0536
01FC
FDB6
FAC5
FA37
FB15
FBB8
FB7C
FAF0
FAC4
FAF4
FB17
FB0E
FB16
FB4A
FB66
FB31
FAE5
FAE6
FB37
FB77
FB6F
FB5F
FB8D
FBC7
FBA6
FB3C
FB1C
FB7B
FBB3
FB1F
FA5B
FB0B
FE07
0218
04FB
059F
04FB
049A
04DF
0514
04C9
047B
04B7
052D
052B
04A5
044B
0483
04E4
04E1
0497
0491
04E3
04FE
0493
0420
0443
04D0
0503
04A1
0461
04DE
0578
04B4
01E6
FE24
FB5F
FA8E
FAFF
FB63
FB2E
FAD3
FAE1
FB44
FB82
FB66
FB2B
FB14
FB1F
FB2E
FB55
FBA8
FBE8
FBB6
FB23
FAC7
FB0B
FB8B
FB90
FB12
FAD5
FB52
FBDA
FB73
FA7A
FAB7
FD6F
01A2
04D0
0585
04A8
0423
04B2
0573
0574
04E9
04A7
04EC
0532
0514
04D8
04E1
0508
04E2
0473
043D
0487
04F3
0502
04C1
049F
04B9
04B5
0470
0467
050D
05CE
053E
028D
FEAB
FB9C
FA9F
FB29
FBBF
FB92
FB05
FAC4
FADD
FADF
FAA2
FA7B
FAAC
FAFC
FB0F
FAF4
FB00
FB37
FB38
FADE
FAA2
FB03
FBB7
FBE8
FB4E
FAA6
FABD
FB4E
FB5D
FAC6
FADD
FD03
00D4
043F
0591
0510
0454
046A
04FB
053E
0517
0504
053C
056A
0545
0501
04F5
0510
0501
04CA
04CA
0528
0578
0544
04BF
0496
0504
056F
0540
04C6
04D8
0574
054C
0314
FF36
FBBF
FA68
FAEE
FBA1
FB61
FA9A
FA52
FAC2
FB3A
FB32
FAED
FAE7
FB19
FB20
FAEA
FAD9
FB1D
FB5F
FB44
FAF5
FADF
FB04
FAF8
FA9E
FA6F
FAC9
FB3C
FB00
FA3E
FA56
FC83
0053
03D9
0583
056F
04E7
04D7
0518
0524
04F6
04F4
0538
055A
050B
0490
0470
04C1
0516
051E
0501
050D
052D
050A
04AB
048F
04F6
0569
0546
04C3
04C7
0591
05E3
041C
003B
FC45
FA5B
FAA8
FB85
FB87
FADA
FA85
FADC
FB40
FB2C
FAE4
FAE8
FB34
FB62
FB55
FB4C
FB56
FB26
FAA7
FA5D
FAC3
FB84
FBC4
FB4B
FADA
FB1D
FBA0
FB59
FA46
F9F1
FBDF
FFBF
037A
0544
052A
0499
049F
0507
051C
04C3
0488
04C8
0530
053C
04EA
04A8
04B9
04E7
04E6
04C9
04D5
0508
0516
04DF
04B1
04CD
04F1
04B3
044A
0471
054E
05B2
041D
008C
FCD4
FAE9
FAF6
FB86
FB68
FADA
FABC
FB28
FB62
FB04
FA8D
FA9E
FB18
FB60
FB51
FB57
FBA0
FBBE
FB52
FAC1
FAC3
FB51
FB9F
FB3E
FACB
FB13
FBCA
FBD3
FAE0
FA57
FBF0
FFA6
0371
0548
050B
043D
042B
04BC
0526
0525
0525
0563
0586
052A
0490
0454
0499
04E2
04C4
047B
0483
04D7
04FA
04B1
0465
0485
04D6
04CF
0481
04A2
0567
05B6
0412
006E
FC9E
FAA4
FAC6
FB93
FBB2
FB2A
FACE
FAF1
FB20
FB02
FAE3
FB27
FB96
FBA3
FB3D
FAF5
FB28
FB79
FB5C
FAEE
FAD3
FB41
FBA6
FB7D
FB1C
FB38
FBBA
FBB5
FACF
FA3E
FBBE
FF75
036C
0572
0549
0490
04A5
0543
0558
04AE
0430
0487
0532
053E
0492
03FC
0417
0493
04D0
04BB
04B7
04E4
04F6
04CF
04C9
0520
0569
0511
0459
0439
0507
059C
044C
00D7
FCF0
FAA4
FA6F
FB1C
FB5B
FB00
FAB8
FAE6
FB3F
FB60
FB5D
FB7B
FBB0
FBB4
FB7B
FB51
FB61
FB66
FB16
FAAA
FAAD
FB38
FBA7
FB6B
FAD8
FAC6
FB5A
FBB1
FB21
FA7F
FB87
FED5
02DB
054D
056E
048F
0451
04EC
0575
0555
04EE
04CC
04DC
04BB
0476
0473
04C3
04F3
04C6
049D
04E2
0551
0544
04B0
044B
0493
050B
04EB
0457
0453
0545
05F9
04AC
011C
FD18
FAD2
FACC
FBAA
FBE1
FB36
FA87
FA7A
FACB
FAE7
FAC9
FAE2
FB5C
FBC7
FBB1
FB3C
FAEE
FAFB
FB12
FAF3
FADC
FB25
FB9A
FBAE
FB4E
FB10
FB57
FBA4
FB4D
FAC1
FB78
FE44
0211
04C6
0569
04E7
04B0
0518
0573
0551
050A
0507
051F
04F9
04AB
049B
04D2
04EB
04BD
04A0
04DC
0521
04FA
048C
0471
04D3
0515
04AB
03F7
03EF
04D1
058E
04B1
01D7
FE1E
FB34
FA13
FA6E
FB32
FB7D
FB3C
FAF1
FAFC
FB3A
FB5C
FB55
FB51
FB57
FB3A
FAF7
FADD
FB22
FB76
FB66
FB08
FAEA
FB3A
FB7C
FB4F
FB13
FB4E
FBB5
FB7F
FAE1
FB6F
FE5C
029D
059A
05E5
049E
03DF
0452
04FC
04FA
04A1
04AB
0511
0533
04DC
0486
0490
04C8
04D9
04CD
04D3
04E4
04E9
04FE
0530
0532
04CB
0461
0494
050D
0457
0177
FD72
FA9F
FA38
FB33
FBBE
FB52
FACF
FAF1
FB6E
FBA4
FB79
FB4C
FB48
FB4C
FB43
FB41
FB40
FB24
FB0D
FB3E
FB98
FB98
FB24
FADA
FB26
FB7B
FB1B
FA94
FB98
FEE9
02FE
0566
056A
048E
0470
0500
053D
04E7
04A6
04CF
04ED
04AC
0472
04B5
0524
050F
047B
0416
0437
0477
0480
049D
0504
053E
04E4
0487
04F7
05A4
04B9
014D
FCF4
FA4F
FA36
FB1A
FB43
FAC2
FAA9
FB34
FB99
FB60
FB03
FB0A
FB49
FB59
FB4B
FB72
FBAE
FB9A
FB4C
FB4D
FBB2
FBDC
FB77
FB17
FB42
FB7C
FB0B
FA8D
FBB5
FF25
0332
0581
058D
04DC
04CF
052E
0526
04C4
04AF
04EE
04E5
0472
043B
04A2
051E
0508
049C
0491
04F1
050F
04AC
0465
04A1
04DE
0494
043B
0486
04DF
03A9
005A
FC95
FA89
FA97
FB45
FB50
FAF4
FAF4
FB44
FB5D
FB3C
FB4F
FB8C
FB6F
FAEA
FAA6
FB0C
FB92
FB7F
FB02
FAE5
FB4D
FB90
FB61
FB53
FBBC
FBE3
FB2B
FA98
FC11
FFE5
03F6
05DF
0581
04B3
04C5
0540
0531
04B4
0490
04E6
0524
050C
04FC
0529
0536
04E2
0487
0495
04D2
04B6
0457
0452
04B8
04D7
046E
0446
04F1
0565
03D7
001A
FC37
FA5C
FA9A
FB4B
FB44
FADE
FAD4
FB07
FAEE
FA94
FA7D
FAC6
FB07
FB0D
FB14
FB43
FB64
FB5C
FB76
FBDA
FC0E
FB8D
FABF
FA9E
FB3A
FB78
FAC8
FA7A
FC67
0074
0449
05CE
054A
049B
04D4
0565
0578
0530
0526
0562
0578
0554
0542
0546
050D
048A
042C
0440
0480
0496
04AA
0507
055C
0512
0465
045E
0539
0581
0382
FF86
FBCB
FA2E
FA69
FAF1
FAED
FABC
FAD4
FAF9
FAD7
FAA8
FAC5
FAFA
FAE3
FAA4
FAC3
FB4A
FBA8
FB87
FB45
FB51
FB78
FB45
FAE5
FAF2
FB5F
FB5C
FABC
FACC
FD00
00F8
048E
0604
05A2
04F2
04E5
0537
0557
053A
051C
0502
04D9
04C5
04E2
04FA
04DB
04B8
04DE
0520
0508
04A3
0492
050D
055D
04D5
0418
046A
05A9
05C6
0309
FE68
FABE
F9CB
FAA9
FB5C
FB20
FAB3
FAC1
FB08
FB0F
FAF7
FB1B
FB5A
FB4E
FAFE
FAD2
FAF4
FB2A
FB4B
FB6E
FB85
FB4A
FAC6
FA9F
FB3C
FBEC
FB9B
FA8E
FAA6
FD4E
018C
04DC
05CD
0534
04B8
04ED
053B
052A
04FC
0500
0507
04D1
0490
0499
04D9
0503
0511
0525
0522
04D5
047F
04AE
055B
05AC
050F
043E
0461
052D
04C6
01F5
FDE9
FB09
FA5D
FAD9
FB15
FAF6
FB21
FB9E
FBC0
FB4D
FAE6
FB0E
FB63
FB4C
FAE7
FAC5
FB01
FB2F
FB21
FB1C
FB3D
FB34
FADD
FAB4
FB24
FBA2
FB56
FAA2
FB3E
FE36
0254
0537
05CA
0514
0496
04AE
04CA
04A0
047D
0495
04AD
04A4
04BB
050F
053F
0500
04A9
04B3
04FA
04FC
04BD
04CB
0535
053E
047F
03DF
0474
0599
0516
01C5
FD4C
FA7D
FA4D
FB3F
FB95
FB32
FB06
FB5B
FB97
FB5F
FB1D
FB34
FB60
FB44
FB11
FB24
FB55
FB3D
FAF1
FAEC
FB39
FB51
FB08
FAF6
FB85
FC0B
FBA1
FAD1
FB7A
FE8C
0287
04FF
053C
04A4
04A9
0531
0550
04DA
0480
04AF
0502
0502
04D1
04C1
04C2
04AA
04A4
04E2
051E
04EB
0475
0452
0495
0499
0418
03DE
04AC
059C
04AE
013B
FD1E
FACD
FAB9
FB4F
FB3D
FAC9
FACC
FB3A
FB5E
FB13
FAF1
FB3E
FB79
FB3B
FAEB
FB10
FB71
FB73
FB18
FAF5
FB44
FB97
FBA8
FBC3
FC17
FC0B
FB24
FA58
FB7F
FF0F
031F
0551
0552
04B8
04C7
052E
051F
04BC
04BD
052F
0556
04E4
047B
04AF
051F
0518
04A0
045A
0482
04B6
04B5
04AE
04C2
04A5
043F
0423
04BE
0534
03E9
0083
FCC1
FABB
FAB6
FB44
FB3D
FADD
FAD7
FB23
FB35
FAF6
FAD7
FB09
FB2D
FB0C
FAFE
FB46
FB94
FB84
FB4E
FB64
FB9F
FB7B
FB09
FB00
FB97
FBEF
FB58
FACF
FC35
FFDB
03AF
0570
051C
047E
04BA
0542
0531
04BD
04B5
0528
055B
04FA
0493
04A4
04DE
04C3
047E
0483
04C0
04C3
048C
0491
04DC
04DF
046C
0444
04F7
0577
03E0
FFE6
FBBE
F9E4
FA7C
FB93
FBA3
FAFF
FABC
FB0E
FB51
FB30
FB08
FB28
FB54
FB49
FB30
FB46
FB64
FB55
FB44
FB6F
FB9B
FB69
FB11
FB2C
FBAD
FBB0
FADF
FA85
FC68
006F
044E
05EB
057C
04C9
04DC
0536
0525
04D2
04C5
04EB
04D0
0480
0479
04CC
04EF
04A6
0473
04BC
0516
04EC
047D
047C
04DC
04D8
044A
041E
04DE
0550
0392
FFA0
FBCF
FA45
FAB8
FB47
FB02
FAA1
FAE8
FB6F
FB6B
FAF1
FACC
FB3A
FBA2
FB92
FB52
FB45
FB49
FB1D
FAF7
FB26
FB76
FB7F
FB67
FBA2
FBFC
FBA6
FA9D
FA74
FCC4
00F6
0478
057D
04C8
044F
04C6
0551
0539
04E3
04E5
050B
04CE
045A
045B
04E3
053C
04F9
0495
049C
04DA
04D0
0492
048A
04A3
046E
0418
0464
0548
0541
02D8
FEBC
FB6A
FA89
FB4D
FBD7
FB7B
FAF4
FAE4
FB09
FB04
FB05
FB48
FB78
FB2A
FAAA
FAB0
FB42
FB9D
FB5F
FB18
FB4F
FB9E
FB6D
FB15
FB60
FC1A
FC16
FB15
FAC8
FD08
0148
04D8
05CD
04EE
043B
0473
04D1
04BC
049C
04E9
0550
0542
04E4
04C8
0502
050D
04B5
046F
0494
04D1
04CB
04B4
04D1
04D3
0458
03DD
0447
0552
0534
028C
FE52
FB17
FA4D
FB05
FB8B
FB5F
FB20
FB21
FB0C
FAC7
FAC5
FB36
FB94
FB5E
FAEB
FAEC
FB55
FB72
FB13
FAE1
FB49
FBBF
FB9F
FB3E
FB55
FBB1
FB72
FAB5
FB17
FDD7
01F5
04F7
059D
04F3
04A0
04F1
0527
04FE
04F3
053A
0553
04EA
047A
049E
0523
0551
04FF
04B1
04B5
04BA
0489
047F
04D7
0511
04AE
0430
0485
0555
04D9
01E3
FD9E
FA99
FA0D
FAE2
FB63
FB2E
FAF7
FB16
FB26
FAEF
FACD
FB0B
FB57
FB44
FAF2
FADA
FB0F
FB38
FB2F
FB34
FB58
FB4B
FB01
FAFC
FB7C
FBD0
FB3E
FA70
FB3D
FE83
02CB
0597
05ED
0505
048D
04DE
0543
054A
0524
0508
04DD
04A3
049F
04E7
0528
0513
04D6
04CD
04F2
04F5
04DA
04F6
053B
0513
045D
03F4
0496
056F
049A
014C
FD0D
FA4A
F9EA
FAC7
FB5B
FB4D
FB21
FB23
FB29
FB1E
FB27
FB41
FB2E
FAE9
FACC
FB04
FB47
FB3A
FB09
FB1A
FB58
FB45
FAD7
FAAE
FB1F
FB8A
FB40
FAE7
FC1C
FF76
0368
05B1
05A7
04A5
0441
04A8
050C
0500
04E5
050B
052E
04FA
04A4
04A8
0512
0565
053C
04D1
04A9
04E3
0516
04E9
0492
0497
050D
0526
03C2
00A0
FCF9
FA9C
FA4F
FB29
FBAD
FB56
FAD4
FAD5
FB22
FB19
FABA
FAA8
FB22
FB93
FB69
FAEC
FAD5
FB35
FB5E
FAFB
FAA4
FB03
FBB3
FBA7
FABD
FA5F
FC1C
FFC8
0377
055E
0562
04C8
04A9
0501
052E
04ED
049D
04AC
050D
0555
0544
0500
04D4
04D5
04DB
04D2
04D3
04EC
04E9
049F
0463
04CC
05BD
05FA
0429
0062
FC79
FA61
FA69
FB35
FB73
FB19
FAED
FB38
FB76
FB38
FAD0
FAD9
FB5C
FBBC
FB87
FB04
FAC9
FAFB
FB35
FB24
FAF4
FB03
FB43
FB40
FAD0
FAA8
FBEB
FEF9
02BA
055E
05F8
053B
0496
04B5
051D
051E
04CB
04B8
0505
052A
04D2
0464
0472
04DD
0500
04A7
0466
04BB
053E
052E
04A1
0490
055F
05DD
0452
008E
FC7D
FA52
FA6F
FB55
FB7D
FAE1
FA8A
FB01
FBB4
FBCD
FB46
FAD2
FAE8
FB43
FB5F
FB32
FB24
FB5A
FB7D
FB40
FAF4
FB1C
FB8E
FB74
FA89
FA04
FBA1
FF9A
03E7
060E
0599
0456
042C
051F
05C6
0556
0489
046C
04F3
0533
04C8
0453
047C
04FF
051E
04BC
047C
04B8
04F5
04AA
043A
0486
0584
05BD
03C2
FFE9
FC40
FA95
FAD5
FB85
FB87
FB0B
FAD4
FB0C
FB2C
FAE3
FA98
FAD1
FB6F
FBC7
FB84
FB0F
FAFC
FB43
FB61
FB1F
FAEB
FB2D
FB8E
FB55
FA93
FA8B
FC8D
005B
040B
05BB
0549
0434
03EE
048A
0524
052E
04FA
0509
054B
054A
04F2
04B2
04D4
050C
04ED
0499
049A
050C
0554
04F4
045C
047B
0554
0584
0395
FFC1
FC01
FA3C
FA90
FB88
FBCB
FB4A
FACF
FAD3
FB13
FB20
FAF8
FADF
FAF0
FAFF
FAF0
FAE9
FB0E
FB39
FB28
FAE9
FAE1
FB46
FBAE
FB7C
FACD
FAC0
FC83
FFFB
038E
0581
0587
04D1
049C
04FE
053A
04F3
04A3
04D0
0540
054D
04D5
046F
0499
0512
0547
0524
0512
0537
0527
0497
040D
0450
052F
0543
034E
FFB9
FC57
FAB5
FAC6
FB4F
FB5C
FAFC
FAC3
FAE3
FB0B
FAF9
FAD7
FAF5
FB4D
FB85
FB62
FB0D
FAD5
FACC
FACD
FAD0
FB0D
FB93
FBEA
FB80
FA9D
FA92
FC98
005A
03F1
0595
053F
046F
046F
0518
0579
0532
04D5
04EC
053F
053B
04DB
04AD
04F5
0547
0524
04BA
04A2
04F8
0524
04BC
0440
0481
0559
0564
035F
FFA9
FC24
FA7B
FAAE
FB67
FB8B
FB23
FADE
FB00
FB24
FAF3
FAAD
FAC7
FB35
FB6B
FB1F
FAB9
FAC9
FB3F
FB78
FB29
FAC9
FAE8
FB4A
FB33
FAA3
FAD5
FD01
00C1
0428
0597
053B
048A
0482
04E3
0506
04E8
04FF
0559
0571
0508
049B
04BF
053F
0553
04BA
042B
0465
052A
0584
051A
04B5
0526
05EF
057B
02CF
FED0
FB8F
FA5C
FAC4
FB60
FB60
FB0E
FB03
FB45
FB5A
FB0E
FABB
FACB
FB19
FB29
FAE1
FAB3
FB05
FB8B
FBA1
FB22
FAA6
FABA
FB16
FB07
FA94
FAE0
FCFE
0092
03E9
058B
0584
0504
04F6
053B
053C
04D6
0478
047D
04C1
04F0
04F3
04F7
050B
050C
04E9
04D6
0501
0538
0516
049F
0470
0507
05DA
0579
02E7
FEE4
FB81
FA42
FAC4
FB62
FB1B
FA73
FA75
FB3A
FBD9
FBAC
FB1B
FAEB
FB2D
FB4C
FB0C
FAEC
FB49
FBAB
FB64
FAA7
FA63
FAEF
FB61
FAC9
F9CD
FA5B
FD7C
01DF
0509
05C6
0511
049A
04F0
0557
0521
048F
044F
048B
04D8
04E1
04D2
04F1
052B
052A
04DD
049E
04B6
04F6
04F2
04B2
04D0
05AB
0684
05C9
02A4
FE2D
FAB9
F9CA
FAB9
FBA1
FB70
FAC0
FAAE
FB4F
FBC0
FB75
FAEF
FAEA
FB4D
FB60
FAE9
FA8A
FAD2
FB66
FB7E
FB0C
FACF
FB33
FB94
FB23
FA46
FA97
FD30
0139
048F
05C4
054E
04A4
04A0
04F5
0506
04C9
04AB
04D5
04FA
04D8
04A8
04CA
052E
055C
051B
04C8
04D4
051B
0511
049D
0465
04F3
05A5
0500
023E
FE63
FB6E
FA7D
FAF4
FB72
FB54
FB04
FB0A
FB48
FB4B
FB07
FAE7
FB20
FB5E
FB3A
FAD3
FAAE
FAFE
FB60
FB63
FB22
FB15
FB52
FB57
FACA
FA4B
FB21
FDEB
01BC
04B9
05BA
052F
0477
0471
04DD
050D
04D6
04A5
04CF
0526
0542
0516
04E9
04E3
04D9
04A7
0481
04A9
04FC
050C
04C4
04AB
0530
05BF
04FD
022B
FE3C
FB2C
FA36
FACF
FB78
FB61
FAF5
FAEC
FB45
FB68
FB14
FAB3
FABE
FB12
FB35
FB11
FB06
FB4B
FB85
FB50
FAE6
FAE2
FB4B
FB63
FAAD
F9F9
FADE
FDFB
0206
04E5
05A3
0514
04A5
04D8
052B
051C
04D5
04C4
04EC
04F1
04B7
0492
04C7
051C
0523
04D4
049A
04BB
04F1
04D2
0484
04B2
0591
062F
0516
01D1
FDAE
FAC4
FA1E
FAF2
FBA7
FB74
FAD6
FAA5
FB06
FB6F
FB78
FB4B
FB3F
FB4C
FB32
FAF6
FAEF
FB40
FB8E
FB78
FB28
FB1F
FB63
FB53
FA93
F9FC
FB1A
FE75
02A7
0576
05ED
0511
0482
04BD
0505
04BA
0443
0461
050B
0575
0528
049D
0485
04CF
04D5
0465
041C
047E
051D
0529
04A5
0489
0558
0607
04D6
0151
FD16
FA5D
F9E9
FAB0
FB4A
FB5B
FB5D
FB96
FBAF
FB55
FACF
FAAF
FB08
FB5E
FB57
FB35
FB6F
FBEC
FC0D
FB7E
FACA
FABE
FB51
FB93
FAE9
FA34
FB33
FE9D
0304
05FA
065C
0530
044F
0476
04F5
04FF
04B6
04B9
051B
0549
04F5
048F
0499
04DC
04BC
0431
03F3
0474
051C
0507
0459
0433
051F
05E8
04A8
0100
FCCF
FA6B
FA5E
FB34
FB62
FAD5
FA82
FADF
FB53
FB2F
FAAB
FA8D
FB13
FBA4
FBA6
FB43
FB16
FB49
FB67
FB29
FAF9
FB5E
FC0B
FC09
FB0C
FA4A
FB7D
FEEF
02EA
054D
0591
04F8
04E3
055E
0591
0523
04B1
04D3
053A
0530
04AF
046F
04DF
0574
055E
04B0
044F
04B7
0542
0507
0432
03E4
04AE
0581
0497
0169
FD6A
FAAC
F9FF
FA83
FAF1
FAE4
FAD0
FB09
FB4A
FB2F
FAD9
FABF
FB05
FB45
FB25
FADE
FAED
FB53
FB88
FB39
FAD6
FAFF
FB8F
FBA8
FAF1
FA6C
FBAA
FF02
02EB
0564
05D0
0537
04E1
0509
0519
04CF
049B
04EA
0572
058C
0516
04A2
04AE
0502
0515
04D5
04BD
0508
053E
04D5
0422
0420
0511
05B5
0451
00AE
FC9E
FA56
FA55
FB3A
FB84
FB15
FAD5
FB33
FB9C
FB62
FAB7
FA68
FAC6
FB53
FB80
FB64
FB6B
FB90
FB5E
FABE
FA55
FAB7
FB6D
FB63
FA77
FA28
FC2B
004E
0449
05F0
054A
0437
042C
04D6
0517
04B6
0481
04F0
056E
0546
04AD
0463
0493
04AC
0469
044C
04CD
0579
0583
0504
04DA
051E
0485
01E5
FE0A
FB32
FA9D
FB55
FB97
FAFA
FA80
FADF
FB84
FB8E
FB13
FAD7
FB20
FB73
FB70
FB57
FB77
FB98
FB64
FB09
FB00
FB34
FB18
FAB5
FB2A
FD77
0108
0408
053D
0522
04F1
0516
0515
04AD
0469
04C0
0542
052F
048E
0437
049A
0521
0510
0494
046E
04C5
04F7
04B5
049E
0533
058A
03F0
001D
FC09
FA11
FA7A
FB72
FB68
FAAF
FA88
FB32
FBC0
FB8A
FB10
FB13
FB78
FB99
FB57
FB32
FB5B
FB5E
FB00
FAD3
FB4F
FBCA
FB3F
FA23
FA8C
FDDF
02BA
0616
0672
0530
0490
0510
0576
04FB
045D
048F
0541
0560
04B2
041E
044C
04CF
04EA
04AE
04AD
04EB
04E7
049F
04CA
0593
05A1
0361
FF24
FB47
F9D3
FA6E
FB2E
FAFE
FA84
FAB5
FB5E
FB98
FB2E
FAD3
FB01
FB60
FB72
FB57
FB6B
FB87
FB43
FACE
FAD8
FB70
FBA9
FAEB
FA44
FB92
FF41
036C
05C4
05DA
051F
04E6
0528
0535
04F4
04D5
04F5
04F8
04BC
049D
04CC
04E4
0491
0443
049B
0555
0571
04AD
0422
04CF
05D1
0501
0188
FD33
FAAB
FAA2
FB72
FB69
FAAA
FA6C
FB07
FB92
FB5A
FAD9
FAE5
FB69
FB9D
FB40
FAF0
FB2D
FB8F
FB7D
FB27
FB34
FB8F
FB63
FA97
FA9D
FD01
0145
04F1
0613
0530
044C
047E
0518
0524
04CC
04D0
0536
054D
04CF
045E
048E
050F
0530
04E4
04B2
04BF
049D
0436
043B
050A
058E
040D
0051
FC4B
FA3F
FA79
FB5D
FB76
FAE8
FAA4
FAF5
FB4E
FB42
FB0B
FAFF
FB06
FAF0
FAE5
FB22
FB6C
FB4B
FAD9
FACE
FB75
FBFF
FB85
FA9E
FB33
FE54
02A6
0590
05E5
04E4
0477
0504
0581
0535
04AA
04A9
050B
0513
04AB
0484
04FA
0575
054D
04C6
04A0
04F0
0512
04CD
04C4
0542
052C
02FF
FEF2
FB3A
F9D2
FA6D
FB32
FB11
FAA1
FABF
FB37
FB4A
FAF9
FAF1
FB5F
FB95
FB26
FAA3
FAC4
FB45
FB57
FAE8
FAC5
FB3C
FB79
FAD9
FA5C
FBDE
FFAF
03CA
05E1
05BC
04FC
04E3
052E
0527
04E9
0506
0568
055A
04B4
043C
0496
0549
056F
04FE
04BD
04FF
0527
04C6
047D
0519
05F3
0524
01C7
FD6D
FAAF
FA7A
FB5D
FB8E
FAE8
FA80
FADA
FB48
FB22
FAC1
FADF
FB6A
FBA1
FB36
FABE
FACC
FB24
FB34
FB00
FB05
FB39
FB01
FA58
FA84
FCD9
00E6
047D
05D2
0538
0469
047C
050F
054F
0523
04FA
04F2
04CA
047C
0464
04A8
04ED
04E3
04C7
04F4
052F
04F4
0474
0496
059C
062C
0479
0076
FC49
FA35
FA6F
FB53
FB7D
FB0E
FADC
FB15
FB3B
FB13
FAF7
FB2A
FB69
FB6B
FB63
FB9F
FBDC
FB8F
FAD8
FA93
FB22
FBA6
FB21
FA2A
FABE
FDEE
024E
053B
05A1
04CE
0487
04FF
0532
04B1
0448
04AD
0567
0582
04EB
0474
0487
04A3
0449
03E3
041F
04CD
0510
04B7
049A
0530
0559
0370
FF84
FBC2
FA3B
FACB
FBA8
FBA6
FB34
FB28
FB68
FB4E
FAD0
FA94
FADC
FB23
FAFF
FAD1
FB23
FBB4
FBD2
FB74
FB53
FBAF
FBB8
FADB
FA22
FB77
FF3D
036C
0591
054E
0452
0420
0497
04D9
04B9
04BD
0509
0520
04D2
04A9
0518
05A9
059F
050B
04AE
04C6
04B2
041F
03E0
04D1
0618
0580
0201
FD5A
FA70
FA51
FB6D
FBCF
FB49
FAFD
FB66
FBC2
FB67
FAD3
FAE2
FB76
FB9F
FB01
FA59
FA66
FAEA
FB32
FB32
FB67
FBBE
FB73
FA7B
FA54
FCA4
00FB
04CD
0604
0519
042B
0467
0509
04F1
044B
0414
0491
0502
04DA
0489
04B6
053A
0568
0516
04C4
04BD
04AF
0470
0481
0532
058E
0403
0059
FC6E
FA75
FAB4
FB8E
FBA2
FB2A
FB1A
FB8D
FBC6
FB6E
FB14
FB3A
FB8A
FB68
FAEE
FAC0
FB0B
FB47
FB26
FB1F
FB97
FBFA
FB73
FA85
FB0F
FE28
0271
0543
057E
047F
042F
04CD
0531
04B9
0422
043E
04C5
04E7
0495
0483
04F1
053F
04F2
0486
049E
04F0
04B9
041A
0426
0523
0578
0350
FF0F
FB51
FA24
FAEA
FB8C
FB20
FA98
FAF9
FBD5
FC15
FB91
FB21
FB47
FB8E
FB6C
FB19
FB13
FB41
FB35
FB10
FB5E
FC03
FC05
FAFE
FA40
FBBD
FF9E
03B5
05B2
0579
04C1
04C9
0528
0501
0473
044D
04B3
04F2
04A9
0463
04B6
053C
0525
047C
0424
0481
04D7
047E
040D
048C
0587
0507
01DE
FD79
FA90
FA42
FB34
FB92
FB23
FAE9
FB4E
FBA2
FB5A
FAEA
FAF3
FB41
FB37
FAE4
FAF0
FB77
FBC4
FB6B
FB11
FB76
FC1E
FBD6
FAA8
FA6C
FCC8
00FD
0482
05A9
051A
048A
04AF
04F9
04D6
048B
0497
04EC
0525
0528
0529
0525
04E0
046C
0441
0496
04EA
04AF
0429
043C
0512
0570
03DA
0058
FCBB
FAD3
FAC6
FB46
FB4A
FAF8
FAF7
FB4F
FB6E
FB1A
FAC6
FADC
FB1F
FB1A
FAEE
FB1F
FBA6
FBD5
FB5F
FAEB
FB28
FBA7
FB65
FA95
FAFD
FDF4
0259
0572
05D6
04C1
0444
04D1
0550
050F
04A4
04C6
0529
0511
0491
0469
04C4
04F1
0489
042A
047A
050E
0500
0471
047B
055D
0582
0330
FEE1
FB25
F9FC
FAD7
FBB0
FB78
FADE
FACF
FB2A
FB3F
FAFE
FAF6
FB5A
FBA7
FB72
FB12
FB18
FB70
FB8B
FB4C
FB38
FB84
FB8C
FAD8
FA5D
FBD4
FF9D
03CD
05F8
05AD
049F
046D
04FC
0539
04DE
049C
04D0
04EE
048B
042F
0484
0530
0544
04A4
043F
04A6
052A
04F9
0485
04DC
05AC
050A
01D2
FD70
FA8B
FA1C
FAC6
FAEA
FA89
FA92
FB2D
FB90
FB53
FB0E
FB4B
FBA5
FB78
FAFE
FAF7
FB6F
FBA2
FB2F
FABE
FAFB
FB70
FB21
FA3A
FA66
FCFE
013E
04D3
0627
05B7
050F
0504
0540
052B
04CB
048E
049E
04C2
04C9
04CD
04E9
04F6
04D2
04AC
04CA
050C
0508
04C0
04C7
0561
059E
03FC
003B
FC22
F9FD
FA4B
FB72
FBBB
FB15
FA9C
FAE4
FB64
FB74
FB2C
FB0A
FB20
FB21
FB01
FB0E
FB4D
FB5D
FB1C
FAF8
FB3C
FB69
FAEC
FA57
FB38
FE4C
0250
0514
05A6
0500
0497
04C5
04F3
04CE
04B2
04E6
0519
04E5
0486
0482
04DF
0513
04D2
048E
04C8
053E
053F
04C1
0497
051C
0538
035F
FF94
FBD2
FA15
FA68
FB40
FB77
FB44
FB4D
FB78
FB43
FAD2
FACC
FB44
FB86
FB37
FAF1
FB47
FBBD
FB7F
FAC7
FAA3
FB46
FB87
FAAF
FA1F
FBF9
0038
0439
059D
04CE
03F9
0440
04F2
0521
04EC
04DF
04EB
04B6
046A
0487
04FA
051F
04CC
0497
04D0
04F3
04AD
0496
052A
0568
03A8
FFD7
FC08
FA58
FAC2
FB8F
FB97
FB31
FB14
FB32
FB2D
FB25
FB5E
FB9D
FB80
FB29
FB02
FB0B
FAFC
FAF5
FB5D
FBF7
FBD6
FAD4
FA7F
FC9D
00C5
0463
058D
04EF
0470
04C1
0527
050F
04CE
04CB
04D2
04A2
0478
04A5
04E6
04CD
0491
04B8
0517
04F4
0469
0485
0573
0578
02DF
FE7C
FB17
FA5C
FB3A
FBAA
FB22
FAA6
FADC
FB42
FB46
FB2A
FB52
FB7B
FB4B
FB08
FB17
FB3D
FB19
FAF5
FB4E
FBBA
FB4C
FA4C
FAA0
FDB0
0243
0575
05E0
04E0
046F
04D9
0527
04F6
04BE
04C5
04C1
049B
04A1
04E4
04F7
04AC
0488
04EE
054C
04EC
044D
049E
0592
050A
01BB
FD3F
FA78
FA53
FB35
FB6B
FAFD
FADA
FB28
FB45
FB07
FAF3
FB2E
FB3C
FAF4
FAED
FB6A
FBBE
FB62
FAF1
FB2A
FB8E
FB23
FA6E
FB64
FEEE
0342
05AB
0585
049E
0493
051A
052A
04C8
04B0
04FC
0523
0507
0508
0530
0515
04A9
0477
04BA
04E3
0487
044E
04F8
05A3
0448
006B
FC41
FA53
FAB2
FB70
FB4F
FAD6
FADF
FB3E
FB4F
FB12
FAFD
FB1B
FB07
FAD3
FAFC
FB73
FB83
FB0D
FAEB
FB7F
FBCF
FB0E
FA6E
FC11
002B
0443
05E0
0534
0463
04A6
053F
0533
04C7
04B7
04EB
04DF
04AE
04CB
0513
0502
04AF
04B6
0519
051D
0488
0445
04F3
0552
035D
FF1A
FB2C
F9EA
FAD3
FBAD
FB70
FAE9
FAF2
FB3D
FB32
FAF5
FB09
FB5B
FB69
FB2C
FB17
FB3B
FB27
FAD6
FAE3
FB61
FB74
FACD
FAD5
FD2F
0162
04EB
05F4
0525
0468
0485
04CB
04A9
0486
04CD
0517
04ED
049D
04AC
04EE
04ED
04C7
04EB
0534
0519
04BA
04E1
0582
0510
0230
FDDD
FAC2
FA46
FB28
FB81
FB20
FB0F
FB98
FBE9
FB8D
FB19
FB29
FB7A
FB74
FB23
FB00
FB1A
FB15
FAFB
FB29
FB65
FAFC
FA44
FB01
FE46
029F
055B
0585
04A7
0489
0522
0552
04CE
046C
04A3
04E7
04B8
0479
04A7
04F7
04ED
04BD
04D6
0501
04C9
0480
04D9
056A
0484
0140
FD1A
FAA2
FAA3
FB80
FB90
FAFD
FAD1
FB25
FB49
FB13
FB0A
FB57
FB7F
FB40
FB00
FB1A
FB45
FB25
FB05
FB4C
FB8E
FB22
FAB7
FC13
FFB1
038F
054E
04EC
0451
04A7
053F
0523
04A1
049F
0512
0529
04B3
046C
04AF
04E8
04A9
0477
04C4
050F
04CB
0481
04E6
052E
0392
FFBF
FBDE
FA4D
FAFF
FBDE
FB9A
FAE9
FAD8
FB30
FB31
FAF6
FB12
FB66
FB58
FAF9
FAF4
FB69
FBAD
FB6A
FB32
FB71
FB8F
FAF7
FAB0
FC97
00B5
0489
05D3
050D
0454
0497
0507
04EA
04AF
04E6
053A
050F
0495
047E
04D5
04FB
04CE
04D2
0511
04D8
041D
03FC
04EB
054D
0323
FEDE
FB3E
FA39
FAFA
FB7D
FB2B
FAF9
FB5C
FB91
FB19
FAAE
FAF7
FB69
FB3B
FACA
FAE4
FB56
FB45
FAC1
FAC5
FB8F
FC00
FB78
FB5C
FD95
01B1
04F2
0590
04B4
0473
050B
0542
04B6
0459
04BE
053F
0523
04B8
04B3
0509
0523
04F8
04FB
051A
04C6
0430
0454
051C
04A9
0197
FD3E
FA83
FA7F
FB8A
FBAF
FAF5
FAA8
FB2C
FB99
FB5C
FB03
FB19
FB49
FB24
FAF5
FB18
FB2D
FAD7
FAA1
FB2C
FBE5
FBAA
FAD4
FB72
FEC3
032A
05BA
058B
0476
0461
0513
0551
04F5
04C4
04EC
04E3
0490
0482
04E7
0524
04D5
0480
04B7
0510
04D2
0457
0498
0533
0433
00A4
FC5C
FA25
FA89
FBA0
FBB9
FB12
FABF
FAF4
FB11
FAE5
FAEB
FB4B
FB83
FB45
FB00
FB18
FB49
FB4A
FB60
FBB1
FBA9
FAF0
FA97
FC4C
0027
040F
05D7
056F
048A
0464
04B7
04D7
04CF
04EF
050A
04DE
04B3
04DF
051B
04F6
04A9
04BD
050C
04E4
0448
0437
0518
0579
0370
FF3B
FB68
FA04
FA8C
FB32
FB3B
FB2C
FB50
FB4B
FB05
FAFE
FB6C
FBB7
FB5D
FAD7
FAE8
FB60
FB66
FAF5
FAF1
FB86
FBA1
FAD1
FAA5
FCFA
0147
04E3
05FE
0560
04DD
0505
051A
04C1
048F
04D6
0502
04AD
0460
04A7
050F
04F1
0494
04AF
051F
051A
049E
049B
053B
04FB
0254
FE11
FAD1
FA15
FACB
FB2D
FAF0
FAE9
FB47
FB6F
FB34
FB1D
FB63
FB81
FB21
FABD
FAE2
FB48
FB49
FB09
FB31
FB9B
FB59
FA94
FB22
FE4F
02C2
05B1
05FE
0519
04CB
052E
054B
04DE
048E
04AF
04C0
047A
0459
04B9
0527
0521
04F6
0518
0536
04D0
0454
049D
0542
0475
012B
FCDA
FA29
FA05
FAED
FB2E
FACD
FABA
FB1A
FB4E
FB28
FB1D
FB5A
FB7F
FB52
FB18
FB08
FAF0
FAB9
FAC7
FB50
FBAB
FB26
FA8F
FBD2
FF87
03B7
05DB
059C
04B9
04A2
051E
054C
0509
04D0
04D0
04CA
04B3
04C8
04F7
04DB
048A
049A
051A
0546
04C2
0469
04F6
056C
03E7
0020
FC29
FA44
FA82
FB34
FB33
FAE3
FAE6
FB09
FAE7
FAC7
FB12
FB72
FB56
FAED
FAE2
FB48
FB88
FB67
FB59
FB8A
FB60
FA96
FA6B
FC85
009A
0433
0564
04CE
0460
04CB
0542
052E
0502
0537
057B
0550
04F3
04F5
053F
0538
04D0
0496
04AC
0488
041E
044B
0548
0585
033D
FEFA
FB63
FA61
FB2F
FBC6
FB65
FAEC
FB0B
FB45
FB01
FA95
FA98
FADA
FAD4
FA9A
FAAC
FB08
FB40
FB48
FB77
FBB5
FB67
FAAA
FAEF
FD83
0199
04BD
057C
04CE
0478
04E2
0537
050B
04D1
04E3
0504
04F6
04F7
0542
0587
055A
04EA
04B6
04BE
049F
047F
04EF
0594
04D7
01C6
FDB0
FAFB
FA92
FB37
FB61
FAF4
FABC
FAF9
FB27
FB07
FAFD
FB3F
FB61
FB1B
FAD2
FAE6
FB13
FAFD
FAEA
FB2B
FB4E
FABA
FA24
FB52
FEF1
0335
0586
0555
0473
0494
0564
05A1
0515
049C
04AD
04DF
04D2
04BE
04DF
04F8
04BE
046B
0465
04A7
04E9
0543
05E3
060E
0460
0093
FC76
FA4E
FA7E
FB70
FB9B
FAFB
FA79
FA8D
FAF8
FB5C
FB9D
FBA2
FB4F
FADC
FAC6
FB22
FB80
FB9C
FBB3
FBCF
FB69
FA61
F9F6
FBC8
FFCF
03E0
05C6
056B
0486
0472
04F8
0547
052F
0500
04CF
0480
0447
0474
04E4
0523
0510
04ED
04D4
049A
0456
0486
052B
051E
0312
FF60
FC0E
FAB8
FAFC
FB60
FB33
FAE7
FAE2
FAED
FAD3
FAE2
FB59
FBCD
FBAE
FB27
FAF1
FB45
FB93
FB75
FB37
FB24
FAF7
FAA1
FB14
FD69
012E
046B
0597
0521
049C
04D1
053E
0548
051C
0515
0507
04AA
0446
0451
04B3
04E5
04C4
04A7
04B2
04A5
0484
04CC
0581
0568
0317
FEF7
FB5A
FA19
FAAD
FB38
FAE4
FA72
FAAA
FB2C
FB36
FADE
FAD4
FB41
FB8C
FB61
FB33
FB73
FBC7
FB9D
FB1D
FAE6
FAFC
FAC1
FA2E
FA71
FCB9
0092
0400
056D
0523
049E
04D0
0563
0592
052F
04AF
0484
04B7
0507
052C
0505
04A8
045F
0479
04F7
056D
0569
0504
04D4
051F
0535
03F1
00F9
FD6B
FAFE
FA76
FB0D
FB7B
FB4F
FB0D
FB2F
FB7D
FB81
FB35
FAF0
FAE4
FAF6
FB13
FB43
FB61
FB24
FAAB
FA98
FB41
FBE8
FB88
FA7D
FAA9
FD66
01A9
04E7
05C1
0526
04C1
04EE
04E1
0452
0407
048C
0547
0552
04D0
04A4
050C
0556
0507
049B
04B0
04F9
04C0
0434
045E
0571
05DE
03E1
FFC3
FBD6
FA19
FA65
FB25
FB50
FB26
FB37
FB72
FB6E
FB2E
FB0F
FB29
FB2F
FB02
FAF4
FB3B
FB80
FB59
FAFA
FB03
FB84
FBB8
FB12
FA6A
FB6E
FEBE
02DF
0586
05CC
04D1
043E
0497
052A
0546
0502
04CF
04D3
04E9
04FE
0510
04F4
0490
043E
0488
0548
0590
04DA
03F6
042B
0546
054F
02B1
FE62
FB1A
FA6D
FB4E
FBB7
FB1B
FA84
FAB6
FB2D
FB23
FAC7
FAD1
FB4A
FB86
FB4E
FB37
FB94
FBC5
FB33
FA79
FABA
FBD3
FC41
FB49
FA78
FC0C
000B
03EC
0568
04E1
045F
04DA
0573
053B
04A5
04A7
0532
055B
04D7
0463
0488
04C3
047B
0419
046E
053F
0564
048A
03F0
04AD
05BE
04DA
0147
FD05
FAAE
FAB2
FB6A
FB6F
FAFF
FAFA
FB61
FB84
FB30
FAEF
FB17
FB51
FB51
FB5F
FBC6
FC17
FBB7
FAF7
FAE1
FBA8
FC19
FB28
F9C7
FA44
FD9C
0217
04FE
0562
04A1
0464
04D6
0517
04C5
0468
0484
04E0
04F5
04B8
047E
046D
045C
0448
046D
04C5
04D5
0462
0409
049E
05C8
05DB
037B
FF5E
FBDB
FA9B
FB1D
FBAA
FB65
FAEE
FB0F
FB95
FBC1
FB6F
FB38
FB73
FBB1
FB78
FB0B
FB03
FB5C
FB82
FB45
FB35
FBA4
FBF4
FB74
FACB
FBA9
FEC7
02B1
0521
0558
049C
0464
04C6
04F1
049A
0441
043E
044F
0438
0444
04C3
0559
0565
04F5
04C0
0505
0511
0459
038E
03D6
04F7
050E
029F
FE85
FB40
FA5F
FB1F
FBB4
FB67
FAF2
FB14
FB98
FBD5
FBAD
FB82
FB86
FB7A
FB31
FADC
FAB4
FAA6
FAA1
FAEB
FBBB
FC7F
FC3A
FAF5
FA5E
FC46
0070
046C
05F8
053E
043D
045A
050D
0525
0486
0420
046E
04D6
04B6
0457
046D
04FF
056F
056E
054B
0537
04E3
043A
03F6
04B3
0586
047B
00E6
FCA0
FA44
FA6A
FB60
FB7A
FAE1
FAB5
FB31
FB89
FB55
FB2E
FB88
FBDD
FB7F
FACC
FAB5
FB3E
FB66
FAB9
FA25
FAAF
FBC5
FBEE
FB12
FB13
FD93
01B2
04E6
05C3
0538
04E6
052E
054F
04EA
0482
0487
04AC
0485
044D
047D
04EF
0508
04BD
04BB
0559
05E7
0586
047D
0400
0480
04C1
0326
FFB1
FC33
FA6E
FA6C
FAEB
FAFA
FAC5
FAE0
FB53
FBA6
FB93
FB56
FB3F
FB4D
FB52
FB44
FB29
FAE8
FA83
FA52
FAC3
FB99
FBF4
FB61
FAD4
FBF9
FF49
0330
0582
05A7
04EF
04C1
051B
0526
04AF
0469
04BB
0517
04D8
044A
043A
04C3
052C
0511
04EB
0529
0556
04D4
0418
043E
052E
0510
0259
FE00
FAC5
FA32
FB21
FB8E
FB0D
FABF
FB3B
FBB1
FB51
FA9B
FA9E
FB5C
FBC7
FB57
FAC3
FAD4
FB3E
FB3B
FADE
FAEC
FB81
FBB1
FB10
FAD2
FCA0
0069
0418
05BF
057C
04D9
04C7
04F1
04D4
04A8
04DB
053C
0537
04CB
048F
04CE
0513
04EF
04AD
04DE
0554
054C
04AB
045D
0504
05AB
0482
010C
FCFC
FA8F
FA51
FAFE
FB47
FB19
FB0F
FB3E
FB38
FAE6
FAC1
FB02
FB36
FAF3
FA93
FAB1
FB2C
FB46
FACC
FA87
FB09
FB99
FB24
FA1F
FA95
FDC1
0235
0523
0562
0466
042D
04EB
0564
04F8
0467
0488
0515
0548
0512
0505
054D
0574
0541
0521
055E
057D
04FE
046E
04D4
05F1
05E2
0335
FEE8
FB9B
FAC4
FB6B
FBC2
FB52
FB02
FB60
FBD0
FB91
FAE4
FA9E
FAED
FB32
FAFB
FA99
FA83
FAA4
FAA8
FA9F
FAE4
FB55
FB42
FA7E
FA25
FBB5
FF44
030E
0518
0513
0458
042B
0487
04A8
045C
043B
04AE
054B
0568
050E
04DC
051C
056B
0561
0527
0519
0523
04F8
04CB
052B
05DC
056F
02AE
FE6A
FB15
FA50
FB54
FC21
FBD5
FB36
FB2A
FB75
FB67
FB05
FAEA
FB2E
FB37
FACA
FA82
FAE0
FB65
FB4B
FAC4
FAB3
FB30
FB3F
FA6E
FA21
FC2F
0062
0438
058E
04D7
041D
0464
04EC
04E5
04B8
051D
05B8
0589
048C
03EF
0469
052E
0517
0456
042A
04F2
05A4
055E
04C5
04F0
0569
0459
00EE
FCD8
FA98
FAC4
FBB1
FBC5
FB2D
FAF9
FB45
FB2B
FA53
F9A5
FA0F
FB3A
FC04
FC00
FBBE
FBBA
FBAD
FB44
FAE8
FB25
FB97
FB55
FA87
FAD4
FD8E
01CA
0504
05BB
04D7
043D
049A
0524
0528
04FA
0532
059D
0592
0501
048F
04A4
04E9
04E9
04BA
04A9
0494
042F
03CE
0434
0543
0574
034F
FF54
FBD0
FA8C
FB12
FB9A
FB3A
FA9F
FAA9
FB2A
FB4E
FAF0
FABC
FB1A
FB87
FB56
FAA4
FA2B
FA4F
FACE
FB57
FBE9
FC5F
FC31
FB34
FA7B
FBB5
FF43
0361
05B5
05A4
04B1
0487
053E
05BE
0569
04BD
0468
0466
045D
0452
0498
0523
0574
0557
0526
052F
0528
04BE
0459
04A9
055F
04EC
0225
FDEA
FA8E
F98C
FA37
FAE7
FADF
FAAD
FAE3
FB48
FB61
FB44
FB5A
FB9B
FB8E
FB18
FAC5
FAF8
FB50
FB3B
FAE3
FAF2
FB69
FB6B
FAA2
FA57
FC49
0070
0484
0646
05C7
04F8
0528
05C9
05AD
04D9
0451
0487
04D8
04AE
0464
049E
052E
055C
0509
04D2
0504
0513
049E
0450
04EC
05A8
0485
00C6
FC56
F9EF
FA34
FB54
FB7A
FAC5
FA6B
FACE
FB30
FB19
FAFE
FB51
FBA1
FB5C
FAD5
FACF
FB3E
FB4E
FABB
FA63
FAFC
FBCD
FB94
FA92
FAC3
FD98
01FC
0553
0634
0583
04E4
04E9
0509
04E1
04C1
04FA
0554
056E
0552
0549
054D
0514
04A9
0482
04D2
051E
04E0
045E
0466
050C
051C
0338
FF8F
FBFF
FA54
FA95
FB49
FB4A
FACE
FAB1
FB24
FB7D
FB2F
FA7C
FA08
FA0C
FA49
FA87
FAC7
FAF9
FB00
FB00
FB51
FBDD
FBF4
FB45
FACD
FC25
FF95
0357
053F
0500
0431
043E
04EA
053B
050B
050D
0582
05CF
0581
0519
054D
05E4
0600
056C
04EF
051C
0569
050C
044D
0436
04D9
04B8
0264
FE68
FAFF
F9E2
FAA9
FB95
FB8A
FAE2
FA83
FAB3
FAFA
FAEF
FAA9
FA87
FAA8
FAD6
FADD
FAC5
FAB4
FAAD
FAA1
FAA9
FAF2
FB53
FB47
FAA0
FA2B
FB4C
FE86
0293
0557
05D7
050B
049A
0514
05B5
05AB
0525
04DD
0511
054A
0527
04EB
050D
057E
05B3
0562
04E1
04B2
04DB
04FB
04E4
04EA
0558
05AB
04B3
01C7
FDC7
FAA3
F9AD
FA66
FB2B
FAF9
FA44
FA1C
FABC
FB63
FB69
FB09
FADD
FAF5
FAEC
FAA6
FA96
FB08
FB90
FB8B
FB0A
FAC9
FB24
FB86
FB3C
FAB5
FB66
FE33
0236
055E
065B
05B6
0500
0522
05A9
05AA
0500
0462
0464
04CD
04FF
04D3
04B7
04F6
0542
052F
04DD
04CA
04FE
04ED
045F
03FD
047D
0545
0496
017F
FD46
FA60
F9F4
FADE
FB48
FACC
FA74
FAFB
FBC9
FBE4
FB54
FB03
FB5D
FBB7
FB56
FA8D
FA58
FAFD
FB9F
FB70
FACC
FABE
FB84
FC28
FBCC
FB0D
FBA3
FE7B
0280
0588
0654
057F
0492
0471
04D1
04FF
04C7
0482
0481
04B0
04D7
04EC
0504
0512
04EB
049D
0485
04D9
053A
050F
045C
03F5
0479
0532
0474
0165
FD47
FA7A
FA2A
FB41
FBD6
FB4D
FAA8
FAEB
FBBF
FC07
FB67
FAAE
FAA5
FB1F
FB64
FB41
FB26
FB50
FB63
FB18
FADF
FB50
FC20
FC3C
FB3B
FA59
FB6C
FED6
02D9
053B
0562
048E
043D
04A5
04FB
04C4
0468
0482
04FC
0537
04EE
0487
047F
04C5
04EC
04D1
04C2
04E7
04EC
0477
03E4
0406
0507
05BF
049E
0154
FD61
FAD4
FA7A
FB63
FC16
FBF2
FB64
FB09
FAF8
FAF0
FAE0
FAFB
FB53
FB9E
FB8E
FB40
FB1C
FB44
FB67
FB39
FAF5
FB14
FB88
FBA4
FB03
FA72
FB71
FE96
0299
0551
05B6
04AF
03F1
043E
0500
0564
054C
052A
0530
0522
04DA
0495
0492
04A2
0471
0421
043E
04F0
058F
055E
0495
0447
04F9
05A4
048C
0134
FD2A
FAA5
FA72
FB68
FBE5
FB70
FAC6
FAA0
FAE2
FB03
FADF
FACD
FAFC
FB31
FB37
FB41
FB95
FBF7
FBD2
FB0A
FA5D
FA91
FB61
FBB1
FAFB
FA51
FB78
FEEB
0312
05AD
05EB
04E4
0430
045A
04D1
0505
0509
0524
053B
0506
04A5
048F
04E2
0520
04D9
045C
0463
050B
058E
0541
0493
049B
058D
0613
0480
00B8
FC8D
FA20
FA07
FB10
FBBB
FB9C
FB47
FB43
FB66
FB4A
FAF8
FADD
FB25
FB77
FB71
FB2F
FB10
FB1E
FAFE
FA94
FA5B
FAC6
FB61
FB34
FA26
F9AA
FB73
FF7D
03BD
0602
05F0
04F3
0474
0492
049F
045A
0430
0479
04EA
050C
04DA
04B4
04C7
04D6
04B6
04AC
0515
05BE
05F9
0573
04C9
04E5
05C0
0604
043B
0070
FC6D
FA2C
FA1E
FB0D
FB98
FB7F
FB62
FB97
FBBF
FB76
FAFF
FAEC
FB42
FB71
FB2D
FADF
FB09
FB6C
FB4B
FA86
F9F0
FA49
FB26
FB60
FAAA
FA4E
FBEA
FF8E
036C
058B
058C
04A9
0430
0461
04AD
04B6
04AE
04D1
04FC
04E7
04AB
04A3
04E8
0523
050C
04DE
0508
0578
0591
0501
0460
0493
057F
05B9
03D9
001B
FC63
FA8A
FAC1
FBAF
FBFE
FB87
FB09
FB08
FB4D
FB63
FB3A
FB1E
FB31
FB3F
FB18
FAE0
FAD5
FAEB
FADA
FA9D
FA9A
FB16
FB9C
FB66
FA84
FA4E
FC31
0009
03E1
05B6
0552
0444
040E
04B7
053F
050C
0490
0473
04B9
04EC
04DE
04DB
0511
0530
04EF
0497
04B9
054F
059A
0521
0477
049A
0581
05B3
03B8
FFD6
FC0D
FA3D
FA7E
FB66
FBAC
FB45
FAED
FB0B
FB54
FB59
FB1C
FAEC
FAEF
FB06
FB17
FB31
FB60
FB75
FB42
FAEE
FAE3
FB3E
FB84
FB20
FA53
FA5E
FC6F
0043
040B
05E7
0596
047D
041E
04A6
052A
0501
048E
048E
0511
056F
0537
04B7
047E
049F
04C0
04B9
04BD
04DF
04D2
046D
0431
04C6
05D7
05E1
039A
FF80
FBB1
FA09
FA82
FB8D
FBCE
FB44
FACE
FAEB
FB4A
FB65
FB34
FB14
FB2E
FB4D
FB3F
FB25
FB3C
FB6F
FB6C
FB2C
FB16
FB69
FBB6
FB4E
FA64
FA55
FC6F
005B
041F
05DC
0582
0496
0471
0507
0571
0535
04B7
047E
0489
048A
047B
049F
0500
053D
050E
04B5
04AB
04F1
0506
04AC
045F
04C3
058D
0564
0330
FF67
FBE8
FA4E
FA8E
FB49
FB55
FAC3
FA6E
FAC9
FB6A
FBB1
FB8A
FB5B
FB65
FB74
FB49
FAFC
FAD6
FAE3
FAEE
FAED
FB1F
FB8F
FBBB
FB21
FA39
FA73
FCE1
00DD
045C
05CA
0565
04AA
04A1
0509
0525
04D1
048F
04AE
04E3
04CC
0486
047B
04C3
050E
0525
0535
056A
057A
0500
0435
03F5
04BF
05D3
059A
0327
FF44
FBDD
FA58
FA89
FB33
FB6A
FB3E
FB39
FB7B
FB9A
FB4C
FAE3
FAEA
FB63
FBB9
FB7E
FAF4
FAA7
FAB5
FAC4
FAAE
FAC2
FB34
FB86
FB18
FA46
FA86
FCF6
00EA
0454
05AF
0545
048C
047E
04DE
04FD
04B5
046C
0469
0487
0492
04A3
04E5
052F
0526
04C6
048A
04E0
0585
05C6
055E
04EB
0529
05CD
0572
0305
FF1C
FBAA
FA3B
FA9A
FB53
FB59
FAE2
FAB9
FB26
FBB9
FBFE
FBEE
FBB6
FB5A
FAE2
FA9D
FAE2
FB86
FBD3
FB58
FA82
FA2F
FA9A
FB04
FAAE
FA05
FA82
FD2A
0144
04C5
0619
057C
0478
0445
04C5
0515
04C4
043C
0410
0448
0483
049E
04CC
051A
0536
04EC
0497
04B9
053B
0572
0513
04BE
0530
05FD
0593
02D8
FE98
FB02
F9AC
FA4B
FB62
FBDA
FBC2
FBA8
FBBA
FBB3
FB73
FB3B
FB4A
FB79
FB71
FB2B
FAFA
FB10
FB2E
FAF9
FA94
FA89
FB0A
FB7F
FB38
FA8C
FAEC
FD71
0174
04E2
0623
0587
049E
0472
04AF
0492
041F
040D
04A4
0545
0536
049B
043B
0474
04D7
04E7
04D0
0508
0572
0569
04C6
0455
04D5
05A6
050E
021E
FE02
FB06
FA5D
FB27
FBB3
FB5E
FADE
FAFB
FB85
FBBD
FB60
FAEF
FAEA
FB38
FB6D
FB6C
FB73
FB96
FB84
FB07
FA82
FA8F
FB28
FB80
FB09
FA76
FB4C
FE3C
021C
04D9
0576
04DA
0494
0519
0590
0535
0463
040D
0477
04FA
04FB
04AE
04A1
04E1
04EF
0496
0454
04A7
054E
0592
0544
04FB
0531
055B
0446
0178
FDEF
FB4F
FA6A
FAB1
FB0C
FB05
FAF1
FB2E
FB8F
FB9A
FB3C
FAE2
FAED
FB3A
FB60
FB49
FB35
FB44
FB3A
FAEC
FAA6
FACB
FB2A
FB19
FA6F
FA26
FB8E
FED3
028C
04FE
05A8
0560
0527
052B
0506
0498
0448
0479
0500
0551
052C
04DF
04CC
04EA
04E8
04BB
04BE
0525
0585
0541
047C
0434
0500
05EA
051F
01F8
FDEB
FB25
FA65
FAAD
FACB
FAB0
FAE8
FB73
FBAC
FB53
FAF2
FB06
FB4F
FB4D
FB0B
FAF5
FB1E
FB2F
FB0E
FB0E
FB4F
FB6A
FB07
FA8E
FA9F
FB13
FB2F
FB06
FBD6
FE80
0213
0493
0522
04B8
04A8
051A
0553
0507
04B1
04B2
04CF
04C4
04BB
04E8
050D
04E9
04BF
04F1
054A
0540
04D7
04AA
04F7
0520
04AF
044A
04D2
05AF
04F1
01B5
FD98
FB17
FADB
FB72
FB6F
FAEC
FABF
FB04
FB28
FB01
FB05
FB63
FBA4
FB78
FB41
FB5E
FB7A
FB22
FAA4
FAAF
FB32
FB60
FAF3
FAA5
FB05
FB66
FAE9
FA46
FB73
FF15
0334
053B
04D2
03E3
040A
0500
0596
0573
0525
0504
04D3
047E
0466
04B2
04E5
049A
0435
044C
04C0
0505
0512
0559
05D2
05C4
04F1
044F
04C9
0585
0471
00D8
FCAD
FA82
FABA
FB8B
FB71
FAC7
FAB1
FB52
FBC3
FB76
FADE
FAAA
FAEB
FB4F
FBAE
FBF1
FBDD
FB63
FAEF
FAEF
FB26
FB05
FA9A
FA97
FB27
FB64
FAA9
FA12
FBAB
FFD7
044A
0656
05B4
046B
0430
04C5
0503
04A5
0460
049F
04FE
050C
04EA
04DE
04CE
0498
047D
04BD
050C
04F3
049C
04A4
0515
053E
04CE
048A
0520
05A1
0426
0048
FC21
FA20
FA76
FB4C
FB45
FAC8
FAD3
FB60
FBA7
FB6A
FB38
FB63
FB84
FB46
FAFC
FB07
FB2A
FAFD
FAB4
FAD0
FB3D
FB64
FB2B
FB2B
FB9E
FBC2
FB07
FA7E
FC0B
FFE7
03DD
059F
053F
049D
04DC
055D
0531
0495
0465
04BE
04F9
04CA
04A9
04EB
0532
051C
04EA
04FE
0519
04D3
046D
0489
050F
052E
04A7
045E
04F7
0560
03B6
FFD0
FBE6
FA35
FAA2
FB56
FB37
FACC
FAE5
FB4E
FB60
FB1D
FB15
FB69
FB98
FB58
FB08
FB01
FB08
FAD2
FA9B
FAC1
FB10
FB15
FAF4
FB38
FBC9
FBC9
FAFA
FABA
FCB9
00BB
046E
05DC
0560
04C5
04F3
0555
052C
04B3
048D
04CB
04F5
04D4
04A5
0498
0498
04A4
04F0
0562
057C
0514
04B3
04D2
050A
04B0
0415
044E
056D
05AE
0341
FEC3
FAF6
F9E0
FAC7
FB87
FB2E
FA91
FAA1
FB29
FB6B
FB42
FB1A
FB23
FB2B
FB24
FB4A
FB96
FB9A
FB2F
FAD3
FAF0
FB37
FB26
FAED
FB1F
FB96
FB79
FAB1
FABD
FD2B
0169
04F4
0604
054B
04B2
04FA
055D
052B
04CE
04E8
053E
0522
0486
0419
0441
04A5
04D8
04EB
0510
0519
04D9
04A3
04D2
051D
04EF
0478
0495
0552
0529
0297
FE49
FADC
FA10
FB02
FB92
FAFF
FA54
FA8E
FB51
FBAC
FB72
FB3A
FB56
FB76
FB4F
FB09
FAE1
FACC
FABE
FAEB
FB59
FB9F
FB7D
FB57
FB9D
FBDF
FB45
FA2A
FA73
FD88
023F
05AB
062C
04F9
044D
04D0
056F
054F
04CF
04A7
04CE
04CC
0497
0491
04D0
04FD
04F7
0502
0526
0502
047F
0434
048C
04FE
04CF
045A
04A6
058D
052F
0216
FD70
FA32
F9E4
FB1B
FB97
FAF6
FA8C
FB18
FBC4
FB91
FACA
FA7F
FB01
FB9D
FBAD
FB59
FB1C
FB14
FB23
FB45
FB6F
FB6A
FB2C
FB1B
FB71
FBAA
FB28
FA80
FB59
FE8F
02C4
058A
05EA
0524
04DA
0532
054A
04D2
0466
0482
04DB
04FB
04EB
04EE
04F3
04BF
047E
0491
04E8
04FC
04A7
0469
0489
0493
0433
0406
04BF
059B
04AD
012A
FCD6
FA57
FA60
FB3B
FB39
FA92
FA76
FB14
FB82
FB40
FAE3
FB10
FB86
FB9D
FB4B
FB16
FB37
FB60
FB5D
FB68
FB97
FB99
FB58
FB51
FBC9
FC1A
FB8A
FAC8
FBA1
FEE4
0305
0591
05BB
04E5
04A1
0505
053D
0504
04DA
04FF
051B
04E3
048C
0463
045B
044D
0453
0493
04D0
04B7
0482
04B4
0521
04FA
0417
0399
045E
0555
044A
009D
FC69
FA50
FAA8
FB85
FB58
FA95
FA73
FB08
FB62
FB17
FAC5
FB01
FB8E
FBD7
FBC4
FBA6
FBA1
FB92
FB71
FB64
FB5B
FB22
FAEC
FB3A
FBF0
FC20
FB50
FAA8
FBFA
FF8B
0369
0568
0556
04C4
04E7
056E
057F
0510
04B8
04B3
04BA
04A3
0495
049D
0488
0458
0465
04CD
0515
04CE
0455
0460
04DC
04E7
0441
03E6
0498
054C
0406
005C
FC59
FA57
FA86
FB32
FB18
FAAA
FAD3
FB71
FBA9
FB44
FAE8
FB04
FB45
FB38
FAFF
FB05
FB50
FB87
FB80
FB65
FB4D
FB2C
FB2B
FB9D
FC4A
FC51
FB61
FAB2
FC13
FFC9
03DD
05FD
05BF
04B3
0460
04D1
0525
04F6
04A8
04A9
04F1
0537
054A
0523
04D7
049F
04A8
04CE
04BE
0473
0464
04D2
0533
04CC
03E4
03B0
0495
051E
0362
FF6F
FB98
FA0D
FAB1
FBA6
FBA5
FB16
FAE8
FB2B
FB43
FB02
FAD3
FAFE
FB3B
FB37
FB08
FAF5
FB0D
FB34
FB66
FBA4
FBBB
FB7B
FB29
FB41
FBA8
FBA7
FB16
FB23
FD33
0102
047D
05CE
052F
045B
0478
0515
053F
04DB
0491
04BA
0507
0519
04FB
04EA
04F3
04FA
04EF
04D3
04A6
047F
0492
04DD
04FB
0498
041B
044A
050F
0507
02DD
FF07
FB96
FA32
FA9B
FB51
FB5D
FB02
FAE1
FB11
FB43
FB4E
FB3B
FB06
FAB7
FA94
FADB
FB58
FB92
FB64
FB2B
FB2C
FB2E
FAF8
FADD
FB4B
FBE0
FBBA
FAE5
FAEB
FD33
0124
047F
05B2
053B
04AC
04BF
0503
04FB
04DC
04F9
0522
0500
04B9
04AF
04E9
0511
050B
050B
051A
04F8
04A0
0485
04E7
0541
04F6
045E
0479
053F
0512
0289
FE6B
FB21
FA2D
FACE
FB52
FB1B
FAD1
FAFE
FB4B
FB3D
FAFF
FB00
FB41
FB69
FB60
FB46
FB15
FABA
FA76
FAB0
FB43
FB7F
FB19
FABA
FB13
FBAC
FB72
FA95
FAEA
FDCA
0217
0538
05E3
0531
04DB
0533
0557
04D8
0451
045C
04BA
04E9
04E8
04FC
0514
04F2
04BE
04D3
051E
0529
04E8
04E2
0553
059B
051D
0468
0495
0565
04F9
0203
FDB0
FA9C
FA08
FADA
FB57
FB1A
FAE3
FB22
FB73
FB79
FB68
FB77
FB6E
FB20
FAE2
FB0A
FB4B
FB25
FABD
FAB2
FB15
FB37
FABA
FA48
FA9D
FB4B
FB46
FABD
FB6C
FE73
0290
0546
0599
04D7
04A6
0528
0569
04FF
047D
0469
0490
0496
0491
04B6
04CC
0497
0463
04B2
055A
05A9
055E
050B
0532
0578
053F
04C2
04C9
052E
047C
01A9
FDB2
FAD5
FA35
FAE7
FB57
FB09
FAA7
FAC0
FB1E
FB52
FB5C
FB72
FB8F
FB84
FB57
FB3D
FB43
FB46
FB36
FB1E
FAFA
FACC
FAC2
FB10
FB74
FB47
FA6A
F9F7
FB73
FF0F
0312
0569
0592
04C6
0469
04C6
0545
055F
0514
04A8
045B
0459
04A2
04EA
04D9
0484
0467
04BC
051F
0519
04D1
04C8
0504
04FF
0490
0468
0517
05C9
04C2
0160
FD33
FA93
FA48
FB14
FB71
FB27
FAFD
FB50
FB9F
FB6B
FAF9
FAE0
FB31
FB6B
FB41
FAF6
FAED
FB1A
FB34
FB2F
FB3F
FB6E
FB6C
FB11
FABC
FAF0
FB89
FBC1
FB33
FAB7
FBC4
FED5
02A0
052C
05A3
04E8
045E
0482
04D4
04E1
04D5
0501
0539
0513
04A4
0477
04CD
0532
051C
04B6
04A6
0519
0578
053C
04AD
0479
04B6
04D0
0486
046D
0505
0598
0490
014B
FD2D
FA7E
FA3A
FB50
FC05
FBB8
FB10
FAD1
FAFC
FB27
FB32
FB52
FB89
FB84
FB1E
FAB3
FAB3
FB06
FB2D
FAFB
FAD0
FB02
FB4F
FB41
FAF3
FB04
FB99
FBEB
FB51
FA8C
FB65
FEA7
02DE
0595
05D1
04D5
0465
04D9
0531
04CC
0440
045E
0504
055C
0513
04B4
04C8
051B
052A
04F5
04E6
0516
051C
04C2
047D
04C5
0540
0524
0464
03FA
0495
055F
0490
0177
FD7B
FAD1
FA57
FB0A
FB77
FB3A
FAF3
FB10
FB43
FB22
FAD9
FAE4
FB4A
FB7E
FB2C
FAB6
FAB9
FB33
FB8B
FB66
FB18
FB0F
FB2D
FB06
FAB2
FAD4
FB97
FC22
FB99
FA9B
FB05
FDEF
0223
052A
05C5
04FA
0491
050B
0586
0545
04AC
0489
04E4
0516
04CB
046D
0476
04C5
04E9
04D0
04C2
04D3
04BD
0468
0441
04A1
0528
051B
0478
042C
04E0
05C7
0526
0236
FE33
FB47
FA7B
FAF7
FB49
FAF9
FAA7
FAE0
FB5A
FB74
FB21
FAED
FB2F
FB8A
FB77
FB08
FAD0
FB19
FB87
FBA3
FB7C
FB73
FB91
FB77
FB08
FABD
FB00
FB6D
FB44
FAAC
FB02
FD72
015E
04B7
05F0
056B
04AE
04A6
0504
0530
0535
056D
05B5
0586
04CE
0434
0448
04CA
0503
04B8
0461
0466
0497
049A
048C
04D1
054F
056A
04EB
0484
04F6
05BF
053F
0276
FE61
FB40
FA69
FB25
FBBD
FB58
FA8B
FA41
FA98
FAF5
FAF7
FADB
FAF9
FB40
FB5F
FB4A
FB4B
FB81
FBAB
FB82
FB24
FAEE
FAF9
FB05
FAEE
FAE8
FB1D
FB38
FACD
FA46
FAE8
FD93
0178
0496
0596
050B
0490
04EE
0581
056D
04DC
04AA
051F
058F
054F
049F
0441
046A
049B
047C
0463
04B6
052E
052F
04BB
048C
0506
058F
055C
04AD
048A
052A
0528
02F7
FEE9
FB3C
F9DB
FA82
FB5D
FB3B
FA92
FA6C
FAE7
FB43
FB10
FAC0
FAE1
FB4D
FB73
FB2F
FAF7
FB25
FB78
FB7F
FB40
FB23
FB49
FB62
FB32
FB02
FB27
FB66
FB2F
FAA6
FAF5
FD31
00F1
045E
05E5
05A6
0507
050D
0578
0584
0510
04AC
04B4
04E2
04D1
049F
04B2
0504
051C
04C6
046D
0487
04E6
04F9
04A9
047D
04C9
051E
04EB
047D
04AB
0575
0574
0342
FF58
FBE4
FAA3
FB29
FBAE
FB32
FA5C
FA42
FAEA
FB6E
FB4B
FAF2
FB01
FB62
FB8A
FB57
FB32
FB5E
FB8D
FB5F
FB09
FB0D
FB72
FBA3
FB4A
FADD
FB04
FB97
FBB4
FB19
FAE5
FC91
001F
03C2
0591
0560
049E
0491
051F
0569
051B
04B9
04BE
04F9
04F3
04A6
0471
047B
048E
048C
04A6
04F5
051E
04C9
0446
044E
04FD
0584
052D
0470
0467
0524
052A
0305
FF2F
FBD8
FAA8
FB32
FBC3
FB6D
FABE
FA9B
FB00
FB37
FAF7
FAB6
FAE9
FB5C
FB92
FB78
FB67
FB84
FB82
FB28
FAC9
FAE4
FB69
FBAB
FB47
FAB4
FAB1
FB38
FB83
FB37
FB35
FCD5
0038
03C8
05AB
058F
04C0
0491
050C
055B
0511
049F
0490
04C9
04CD
0480
043C
0441
046C
0491
04CA
0528
0559
0502
0462
0430
04AF
0536
0509
0468
044D
04EF
050F
0342
FFB9
FC4F
FAAB
FAB6
FB18
FAEF
FA8E
FAA3
FB28
FB82
FB68
FB36
FB4F
FB8C
FB8A
FB46
FB1E
FB40
FB67
FB4A
FB0E
FB16
FB69
FB9A
FB70
FB41
FB74
FBC6
FB7F
FA9B
FA57
FC24
FFED
03CF
05C5
0593
04B2
048E
0520
057A
0531
04C8
04CD
0511
0505
0499
0443
0449
046A
0461
0456
048B
04D3
04C1
0466
045E
04F3
0589
055D
04A6
0473
052C
05A2
042B
00A4
FCDF
FADA
FAD9
FB74
FB63
FAB7
FA56
FAA8
FB2F
FB53
FB1D
FAFB
FB17
FB37
FB35
FB40
FB83
FBCD
FBC1
FB60
FB17
FB29
FB4B
FB15
FAAA
FA94
FAF8
FB3A
FAE0
FA90
FBB8
FEE9
02D9
0573
05D1
04EE
0452
047A
04D6
04ED
04EF
0527
0557
051F
04AD
0496
04F7
0538
04E4
0457
043E
0495
04B0
0450
0419
04A2
0570
0579
04A3
0419
04BF
05AE
04E8
01A3
FD69
FAA2
FA41
FB2A
FBC6
FB99
FB3C
FB2A
FB32
FAF9
FAA1
FA8D
FAC9
FAF9
FAE4
FAC4
FAEB
FB4A
FB8E
FBA0
FBBB
FBF5
FBFA
FB7B
FACD
FAA2
FB23
FB95
FB4A
FAC7
FB83
FE41
01F6
04A5
055C
04E9
04A5
04EB
051A
04CC
046D
0486
04EF
0514
04DC
04C8
051A
0560
051E
0494
046D
04BE
04DF
0468
03E1
040E
04C7
051C
04AF
0451
04D7
0598
04D6
01CE
FDE0
FB47
FAD4
FB66
FB83
FAFA
FAA7
FB00
FB82
FB83
FB1D
FAE5
FB09
FB28
FB00
FAD9
FB07
FB55
FB46
FAE2
FACE
FB69
FC2A
FC3A
FB94
FB11
FB37
FB7D
FB1E
FA82
FB2F
FE0C
0201
04DD
0582
04D8
0479
04DF
0545
0506
0482
0474
04E5
0535
0507
04AE
0494
04A9
04A9
04A3
04DA
0528
0509
0464
03E0
041F
04C8
04E7
044F
0400
04CF
05E6
054E
0225
FDDE
FAF2
FA73
FB47
FBB5
FB41
FAB5
FAC3
FB29
FB4B
FB1A
FB0B
FB50
FB8E
FB6F
FB2D
FB3B
FB97
FBC8
FB92
FB53
FB76
FBC8
FBBA
FB41
FB08
FB7C
FC05
FBB6
FACC
FAEB
FD67
017F
04D6
05CE
0509
0457
049A
0524
0516
049E
0484
04EE
0534
04E9
0477
046E
04B1
04BA
0475
0455
048B
04A6
0451
03FA
044B
0515
0564
04D1
042F
0474
0527
04A1
01F7
FE40
FB86
FABA
FB07
FB28
FAD0
FAA0
FB04
FB9F
FBDB
FB97
FB2C
FAE8
FAD6
FAE4
FB10
FB51
FB76
FB5D
FB2E
FB40
FBAB
FC0D
FBF9
FB80
FB34
FB75
FBDA
FBAC
FB00
FB20
FD53
0136
04B5
05FB
053F
0457
0489
0550
0567
049B
03EF
0425
04D0
051D
04FF
0506
054C
0545
04B0
042A
0455
04E2
04F5
0466
03FE
0438
0483
0434
03B9
041B
0538
055E
0316
FF0D
FB8C
FA28
FA6F
FAF6
FB0A
FAF9
FB19
FB3F
FB2D
FB04
FAFF
FB11
FB0A
FAFF
FB2A
FB79
FB86
FB28
FACB
FAEC
FB75
FBE0
FBE3
FBC2
FBDE
FC27
FC27
FB94
FADF
FB19
FD1F
00B0
0444
0618
05B1
045B
03D7
049A
0590
05A2
04FD
0493
04C1
0501
04DA
048E
048F
04BF
04B0
046E
0474
04D0
04F0
048D
0432
046B
04D2
049A
03E8
03D0
04A6
04FB
0319
FF44
FBC4
FA77
FAFB
FBA0
FB89
FB2B
FB1A
FB2A
FB06
FAE0
FB14
FB71
FB6E
FB0A
FAE1
FB45
FBB9
FBAB
FB4D
FB3C
FB95
FBDB
FBB9
FB64
FB3B
FB4E
FB7F
FBC6
FC03
FBD8
FB2B
FACC
FBFC
FEF6
0261
0495
052D
04FF
04DD
04DA
04C9
04C6
04F6
0517
04DE
0489
04A2
0521
0557
04E9
045A
0442
047C
0487
0478
04C5
054C
0543
046B
03B7
041B
0513
053F
046F
03FE
04AD
0514
0333
FF34
FB97
FA68
FB20
FBC8
FB7E
FB07
FB29
FB8D
FB92
FB61
FB7B
FBBA
FB8F
FB08
FAD6
FB43
FBB2
FB8C
FB1F
FB1B
FB8A
FBCC
FB99
FB5C
FB6D
FB89
FB75
FB84
FBF0
FC1F
FB67
FA79
FB23
FE3B
0246
04DC
052A
0477
043F
0498
04C3
0491
0479
04A8
04D1
04D3
04F7
054D
0562
04EC
0462
046B
04DE
04FA
0494
045E
04C9
0537
04EE
043D
0406
0468
04A5
0481
04B9
05A1
05EA
03D8
FFAD
FBE6
FA95
FB3D
FBDA
FB79
FADF
FAE1
FB30
FB1F
FACB
FADB
FB58
FB97
FB4B
FAF8
FB1B
FB6B
FB69
FB38
FB4F
FBA1
FBB1
FB65
FB35
FB5D
FB7D
FB41
FB0A
FB49
FB83
FAEA
F9FB
FA9E
FDEE
0273
056E
05C0
04CE
0476
04FC
055C
0516
04B8
04C2
04E8
04C0
048E
04CD
0551
057B
0522
04B8
0493
0489
046C
0469
04AD
04F2
04E3
04BA
04EB
0542
0514
0478
0476
056C
05D8
03C3
FF5C
FB44
F9D6
FABA
FBBE
FB9C
FB06
FB05
FB63
FB4D
FAB9
FA5C
FA81
FAB5
FAA4
FA9D
FAF8
FB71
FB93
FB69
FB4D
FB39
FAE7
FA96
FAE6
FBBC
FC08
FB38
FA42
FA6E
FB6C
FBAE
FAE2
FAF3
FDC7
0273
05DC
0637
04D5
0423
04BB
0564
0543
04E2
04FD
0558
054E
04F0
04E5
054E
0598
0565
050A
04E6
04D9
04BA
04C8
052A
055E
04DC
040C
03E3
0481
04FA
04BF
0496
0548
05D1
041B
FFCE
FB57
F968
FA0C
FB20
FB2B
FAB7
FAC9
FB35
FB22
FA8D
FA4A
FAA6
FAFA
FAD7
FAB8
FB15
FB75
FB2F
FAA0
FAB6
FB85
FC1B
FBEE
FB9F
FBD7
FC1D
FB92
FA83
FA2F
FAE0
FB6A
FB29
FB75
FDFD
0222
053F
05BC
04C8
0487
0554
05CA
0529
0461
047B
050C
0509
0473
0442
04E2
05A3
05C5
0558
04DB
047A
0431
042B
048B
04EC
04C1
0443
0434
04A5
04B4
040C
03C0
04C3
05E4
04A7
0061
FB92
F959
FA18
FB7A
FB91
FAD5
FABB
FB76
FBFA
FBB2
FB16
FAB9
FA95
FA84
FAB4
FB3E
FBB0
FB91
FB26
FB1C
FB74
FB85
FB1F
FAF4
FB7B
FC0F
FBDF
FB30
FAED
FB26
FB06
FA86
FB2B
FE3E
02AF
05C6
0623
0512
048E
04E5
050A
0499
045C
04D8
0573
0564
04E6
04C5
0518
052C
04B4
0447
0473
04E8
0504
04BD
0472
0445
0422
0438
04BF
054F
0532
0489
0478
0578
0605
03F9
FF69
FB1F
F9AF
FAC2
FBEA
FBAF
FAC0
FA5E
FAA5
FAE1
FADE
FAFC
FB4C
FB5D
FB14
FAF6
FB4C
FB98
FB60
FB00
FB1B
FB8E
FBAB
FB5C
FB3F
FB90
FBA9
FB13
FA86
FAED
FBCD
FBB8
FAB0
FAD6
FDE4
0296
05C6
05FB
04CB
0482
055B
05D8
053A
0474
048D
052C
0555
04F0
04B8
04FE
053F
0509
049D
0478
04AF
04FF
0533
0532
04DB
044D
0419
04A3
0552
0519
040F
03B1
04DF
061B
04DA
00A4
FBFE
F9C6
FA3D
FB4B
FB50
FAB0
FA85
FADC
FAF4
FAA4
FA81
FACE
FB0A
FAD2
FA8F
FAD7
FB87
FBF3
FBD6
FB99
FB95
FB9D
FB78
FB52
FB5C
FB62
FB31
FB10
FB56
FBA6
FB4A
FA83
FAE2
FD9F
01DB
052D
061C
0573
04F3
0545
05BD
05B9
0568
0539
0525
04EB
04A2
04A1
04E9
0517
04E8
0486
0431
03F8
03E9
042B
04A5
04D8
0484
0421
0455
04F2
051D
0490
042F
04BB
0551
040A
005A
FC1E
F9CA
F9E5
FAE2
FB31
FAC8
FA88
FAD6
FB47
FB68
FB3F
FB06
FACE
FAA8
FABF
FB17
FB68
FB7E
FB85
FBB2
FBD7
FBAA
FB58
FB57
FBAF
FBCB
FB58
FAD8
FAEB
FB44
FB12
FA86
FB1F
FDE5
01DA
04DC
05E5
05C0
0590
056C
04E3
0434
042D
04DF
0563
0521
04A7
04BA
0519
04EC
0424
03AF
0424
04F4
053C
04F4
04C1
04E3
04F9
04D6
04D3
050C
0508
0495
0460
04F0
0555
03D2
001C
FC29
FA34
FA5F
FAF9
FADB
FA8E
FAED
FBA0
FBB2
FB16
FAB4
FB12
FBB8
FC07
FC04
FBF2
FBB7
FB24
FAA1
FAD4
FB98
FC01
FB98
FAFD
FAD2
FACA
FA5E
F9FF
FA91
FBD1
FC4A
FB76
FB10
FD48
01D3
05CE
06EC
05CD
04B9
04C0
0513
04C8
041D
03CD
03EF
0428
0465
04CD
0526
04F7
0469
0442
04C6
0533
04E0
0451
047C
0554
05D5
0575
04CC
0491
0492
0455
0424
0497
0516
03E7
005D
FC29
F9C3
F9D1
FAE4
FB80
FB8C
FB9B
FBB1
FB6B
FAEC
FAD2
FB30
FB5F
FB0E
FACE
FB24
FBA1
FB89
FB05
FAF1
FB8E
FC1D
FBF1
FB49
FAD4
FAC0
FACC
FB01
FB8B
FBEB
FB4F
FA1F
FA4D
FD4C
0203
05AD
06B6
0602
0550
052C
0504
0496
0458
047B
0482
0435
042C
04DE
05AB
059D
04CE
0446
0487
04FF
050F
04EB
0508
052A
04CE
0442
045F
0517
054A
0490
041D
04F6
05E0
0469
0015
FB70
F956
F9E5
FAF8
FB1D
FAE2
FB27
FB8A
FB45
FAA3
FA94
FB23
FB6E
FB1F
FAF2
FB78
FC18
FBE6
FB0B
FA88
FAC3
FB25
FB49
FB89
FC03
FBFE
FB0B
FA22
FA77
FB9B
FBE9
FB17
FB2A
FDF8
026B
057A
05BC
04D0
04CA
0591
05B0
04E2
045D
04CE
0558
0513
047A
0494
0545
0571
04B6
0402
0425
04B3
04EA
04DC
0503
0530
04E4
0465
0483
052D
053E
0445
039D
049B
0614
0525
00D0
FBAF
F923
F9A8
FAFA
FB53
FB15
FB3C
FB84
FB0F
FA20
F9F4
FAEC
FBF2
FC06
FB8B
FB68
FB96
FB6D
FAE1
FA99
FACD
FAFA
FACC
FAAD
FAF3
FB2C
FADD
FA8D
FB25
FC4F
FC9B
FBC0
FB9A
FDF9
01FD
04DA
0526
0449
0452
0556
05CE
0513
0435
0450
0505
054E
0506
04D5
0502
052A
050C
04E1
04E3
04F9
0518
056F
05E3
05D9
0507
0435
045F
052A
0539
0448
03DC
0500
062C
04B3
003F
FB9A
F99B
FA23
FAF1
FAC1
FA53
FA8D
FB02
FB05
FB03
FBBF
FCBD
FCBB
FB9C
FABC
FB10
FBC8
FB86
FA5B
F9A9
FA27
FB0D
FB5E
FB27
FAEC
FAB1
FA50
FA3A
FAE5
FBC2
FBBF
FB0C
FB5E
FDED
01AC
0465
0549
0573
05DE
0614
056D
0482
0466
04F7
0518
0473
03ED
042C
0490
0446
03B1
03D1
0499
050C
04FA
055D
067E
06FB
05CB
042E
042C
0592
060F
04B0
0390
04AF
0618
0358
FB25
F1BE
EC90
EC97
EE68
EED9
EDEF
ED45
ED56
ED6F
ED48
ED56
EDA7
ED99
ECF6
EC85
ECE8
EDA9
EE04
EDFB
EDF7
EDDB
ED4C
ECB1
ECE1
EDD1
EE64
EDF3
ED5A
EDB7
EEA5
EEB6
EDA2
ECCD
ED3A
EE2A
EE6D
EE36
EE70
EEEC
EEA5
EDBF
EDC3
EF3A
F05F
EFA4
EEEC
F239
FA84
039B
0850
07E7
0606
05D2
06F0
0769
06D9
067E
06F4
0768
0726
06B6
06CA
070A
06C2
062E
062A
06D2
074E
070F
0679
0638
0656
066B
064D
062F
0635
0656
0689
06A3
0608
0444
020A
00D8
0128
01CB
0194
00F7
0112
019F
013E
FFEF
FFB9
019D
02DF
FF64
F712
EEF1
EBF0
EDA3
EFA0
EF2D
EDB6
EDC0
EF42
F037
EFB0
EEC1
EE80
EEA1
EE84
EE7B
EF03
EF98
EF64
EEA5
EE74
EF33
F01E
F084
F09C
F0EB
F15F
F197
F19C
F1B1
F196
F0E6
F02B
F089
F1F7
F2D9
F218
F0B2
F04E
F0F8
F174
F165
F1B1
F271
F221
F03E
EFA5
F429
FD7E
0664
0A10
090A
0779
07B7
0886
083C
076F
0783
080A
0747
04F8
02EF
028E
030D
0300
0282
02A8
037D
03E9
0379
02FD
0324
0366
02E4
01D7
0152
01CE
02AD
033A
0365
0355
02F3
026E
026E
032B
03CD
0380
02B7
0291
0318
0336
0296
026E
0362
0374
FFBC
F87E
F1EA
EFD2
F179
F2FC
F230
F0A7
F0B2
F217
F2B9
F1C0
F088
F07B
F145
F1C8
F1DB
F220
F2AC
F2DD
F26E
F1E1
F1AB
F1A0
F17C
F170
F1C7
F23F
F255
F217
F20F
F261
F28E
F263
F262
F2D7
F325
F2A4
F1B3
F13A
F161
F17E
F14B
F147
F191
F15B
F079
F0F6
F565
FD49
047C
0733
05DC
03FB
03E3
04CC
0500
045A
03FB
045B
04D8
04F8
04FF
051E
04F1
0459
03FC
044B
04B7
049A
0450
0495
0521
04FB
042A
041F
05DE
0876
0A01
09E3
092D
08E2
08E8
08EC
092E
09BA
09DD
0930
088B
08CF
0951
08C8
07AC
0801
09F5
0A12
04A8
FADE
F275
EFC4
F16F
F30A
F299
F1BA
F21C
F303
F2F5
F233
F23A
F351
F414
F383
F259
F1D6
F207
F21B
F1C2
F161
F136
F120
F125
F175
F1DC
F1DA
F174
F168
F228
F30F
F321
F26F
F1F2
F223
F275
F276
F28F
F314
F362
F2DD
F241
F2CA
F40B
F41A
F288
F228
F64A
FE48
055B
0793
05F6
04C0
0651
0933
0ADE
0AE1
0AA0
0AF5
0B5A
0B34
0ADA
0ADC
0B02
0ABB
0A14
09A8
09BD
0A09
0A3F
0A61
0A76
0A5B
09FF
0998
095D
0947
0936
0941
0985
09D8
09FE
0A1B
0A6D
0A99
0A03
0902
08C9
09A6
0A1D
08BD
0671
0580
0605
04D5
FF35
F6FE
F148
F0C0
F2EB
F3C1
F283
F17E
F213
F2FF
F2BC
F1D3
F1C2
F29A
F310
F2A8
F260
F2DD
F352
F2EB
F246
F275
F33D
F378
F2EA
F28B
F2F2
F37C
F368
F306
F323
F3B8
F408
F3EF
F412
F49A
F4CD
F457
F3F2
F434
F48F
F472
F485
F57D
F64D
F53B
F32E
F438
FB25
053C
0C42
0D12
0A96
0985
0AE6
0C3D
0BF1
0B30
0B72
0C14
0B9F
0A4B
09BB
0A84
0B54
0B00
0A38
0A55
0B3F
0B89
0A62
0865
06A0
0590
0534
0575
0608
065A
060B
056C
0531
059E
064B
06BA
06C2
0666
05C0
0546
0585
0641
0677
05CD
0566
065B
076E
0588
FF39
F722
F1D2
F13F
F340
F491
F44D
F3BC
F3C1
F3CA
F344
F2C2
F322
F433
F4F3
F4F5
F4C3
F4E7
F532
F53F
F524
F521
F514
F4C0
F45E
F459
F495
F48B
F42A
F41F
F4F0
F622
F6B1
F633
F52D
F453
F3F9
F431
F4DB
F56C
F54D
F4D2
F50B
F61B
F67A
F502
F387
F5D9
FD4D
0627
0ADA
09CF
06A9
059A
06F6
082B
07CE
06FD
0709
0790
077E
06E2
06B8
0741
07A8
075C
06DD
06D1
071C
0753
076D
0771
070F
0646
05FD
0705
08AB
0937
0807
0670
060D
06BA
0709
067E
0633
0735
092A
0B0E
0C59
0CCE
0C17
0AA2
0A0F
0B5E
0C93
09D3
01D9
F86C
F30C
F342
F58C
F60C
F4BD
F426
F53E
F664
F61E
F51C
F4DF
F584
F5DE
F563
F4E1
F530
F5FE
F662
F619
F595
F531
F4E9
F4B4
F4AC
F4CF
F4FD
F52D
F55C
F55B
F509
F4B5
F4E7
F598
F5F7
F568
F477
F442
F4F8
F5AE
F5CD
F5CD
F606
F5A9
F421
F320
F5DA
FD43
05EF
0AD3
0A42
074A
05F3
0716
0886
087F
079A
0765
082A
08CA
0863
0769
0713
0810
0A07
0C05
0D44
0D8E
0D38
0CB9
0C45
0BD5
0B8C
0BAA
0C1F
0C80
0C94
0C97
0CBC
0CC1
0C65
0C05
0C33
0CC2
0CDB
0C4D
0C1B
0CF3
0DAE
0CAD
0AAB
0A7B
0D05
0EC0
0AFA
0198
F7F8
F387
F470
F690
F6B6
F562
F47B
F44B
F3EA
F355
F37C
F47A
F529
F4BE
F3DB
F38D
F3E8
F43B
F440
F45D
F4BC
F4ED
F4A3
F43D
F42A
F44F
F47A
F4D8
F573
F5BA
F534
F46F
F46A
F528
F595
F512
F464
F482
F517
F52E
F508
F5D9
F772
F7D3
F644
F5B2
FA0D
032B
0BF8
0F97
0E5A
0C8B
0D01
0E89
0EBD
0D95
0CE4
0D56
0DBC
0D2C
0C63
0C73
0D13
0D28
0C86
0C27
0CA0
0D3C
0D22
0CA0
0CAD
0D72
0E18
0DEA
0D2C
0C99
0C88
0CAB
0C76
0B8E
0A0A
086F
0758
06FD
070B
072D
0775
07E3
07D3
06C3
05A4
0635
085D
0918
054C
FDAE
F69D
F3BE
F47D
F59F
F56F
F4F1
F53D
F58F
F4DA
F3E5
F44F
F602
F713
F659
F4E6
F470
F51A
F5A5
F568
F50C
F53F
F5B7
F5F8
F639
F6D1
F75C
F737
F686
F60A
F626
F69A
F71C
F799
F7EA
F7D7
F790
F794
F7D7
F785
F64F
F571
F636
F7B4
F789
F59E
F588
FAA9
03A1
0B3C
0DF0
0D11
0C2C
0CAA
0D57
0D55
0D7D
0E6F
0EEC
0D7A
0ABB
08C7
0889
08F3
08D7
085C
0848
08A1
08C0
0867
0810
0822
086B
08A1
08D0
0906
0902
08A3
0850
087B
08F0
092E
0924
091A
090B
08A7
0819
080C
08A4
08F4
0848
078B
084A
09F5
095B
040B
FBC3
F55A
F3E0
F5D3
F784
F75B
F6B8
F70C
F7B0
F742
F604
F592
F68B
F7A2
F774
F65E
F5C6
F61E
F682
F649
F5F9
F648
F6F0
F722
F6C6
F67D
F69E
F6CB
F6AB
F67B
F6A6
F717
F76A
F783
F794
F7A2
F780
F749
F74A
F753
F6D8
F5F3
F57F
F5C1
F5DF
F58B
F686
FB1A
02B4
095F
0B8C
09E9
0850
0919
0AE5
0B4F
0A40
0974
09B2
0A10
09BC
0920
08F1
0911
08FA
08BD
08E2
0967
099D
0926
0881
085C
08CC
098F
0A82
0B6F
0C05
0C62
0D29
0E7F
0F7C
0F38
0E1C
0D67
0D88
0DC0
0D7D
0D37
0D68
0D63
0C6F
0B8B
0C72
0E50
0D45
06AC
FD05
F5FF
F4A4
F6C0
F835
F78C
F670
F683
F756
F7A1
F741
F71F
F7A6
F844
F84A
F7AE
F6DE
F656
F654
F69E
F69F
F611
F579
F59E
F687
F753
F73E
F683
F5FA
F601
F628
F609
F5F3
F65C
F70B
F746
F6D0
F63F
F63F
F6CC
F752
F76F
F758
F769
F789
F73D
F66B
F5BD
F5D7
F666
F677
F5C6
F530
F590
F69C
F76A
F7CB
F84D
F8D3
F82B
F614
F517
F8C1
0163
0ABE
0FE6
100A
0E7A
0E5B
0F90
101A
0F3D
0E42
0E6B
0F49
0F99
0F04
0E63
0E7B
0F19
0F85
0F56
0EC8
0E67
0E7D
0EC2
0EAA
0E1C
0DA6
0DDF
0EB8
0F8F
0FD1
0F62
0E88
0D92
0CA1
0BA9
0AA8
09D4
0984
09D1
0A3B
09F8
08E9
0805
0844
0944
09A5
08D5
07C4
0775
07C2
07FF
0832
08C3
0964
0944
0863
07D2
0821
0887
0853
0872
09D9
0AB3
0756
FF1A
F687
F2EF
F4A9
F74D
F75D
F5CF
F57B
F6DF
F7F5
F78A
F6C4
F6FF
F7C8
F7F4
F796
F794
F7F6
F7F4
F779
F755
F7E0
F85F
F82C
F7C2
F801
F8D3
F935
F896
F791
F70A
F71F
F75B
F78C
F7C6
F7F3
F7E2
F7B9
F7C8
F808
F823
F803
F7F5
F831
F887
F88F
F82F
F7C8
F7D3
F847
F88C
F828
F75D
F6F3
F747
F7C2
F78A
F6B7
F657
F6D7
F71D
F647
F5FF
F969
010A
08F0
0C5D
0ADD
0875
08C0
0B20
0C80
0B97
0A0D
09A7
0A0B
09FD
0984
099C
0A62
0AE2
0A99
0A1B
09FC
09EC
0966
08BD
08CF
09CA
0ACB
0AF6
0A8F
0A9A
0B9A
0D0D
0E1D
0E7B
0E69
0E4B
0E4A
0E54
0E5B
0E76
0EB2
0ECD
0E71
0DBD
0D43
0D6D
0E0F
0EB7
0F22
0F4B
0F40
0F13
0ECF
0E54
0D7F
0C9A
0C6A
0D63
0ED0
0F69
0EFD
0ECB
0F36
0DDB
07CA
FE05
F5EC
F3EA
F6A4
F8F2
F7FA
F5B0
F51C
F625
F671
F54C
F499
F5BA
F77E
F816
F79E
F766
F7A2
F76D
F6AE
F662
F6F0
F760
F6D1
F5DF
F5C3
F68C
F719
F6C8
F634
F609
F60B
F5DD
F5EA
F6AF
F7B1
F80E
F7CD
F7BC
F823
F868
F811
F777
F727
F711
F6E6
F6E6
F7A2
F8D1
F93C
F84B
F70B
F6EB
F7CF
F83C
F774
F695
F728
F8FF
FA2D
F966
F829
F9DE
004E
0933
0FEF
11CA
101C
0E35
0DE2
0E73
0EB7
0EBC
0F22
0FA4
0F69
0E93
0E5F
0F4D
1033
0FD8
0EB1
0E35
0ECB
0F5D
0EDC
0D77
0C19
0B53
0B19
0B3F
0B95
0BB5
0B3C
0A5A
09B0
0976
094E
0919
0948
09F8
0A70
0A10
0951
0907
0919
08BD
07E7
07A1
0897
09FD
0A87
0A23
09E9
0A54
0A8C
09DB
08F3
08E5
0979
0982
08C8
0889
09C0
0B6B
0B0C
0700
004A
F9F9
F6B5
F6AD
F7DB
F829
F748
F67A
F6B0
F754
F73A
F669
F620
F712
F862
F8E5
F892
F82D
F805
F7D0
F79B
F7F7
F90C
FA18
FA37
F96F
F882
F7E4
F76D
F709
F705
F776
F7DA
F7CB
F790
F78B
F795
F765
F74A
F7C9
F8A9
F90C
F884
F7A8
F73C
F745
F748
F73C
F77F
F7EC
F7C5
F6E5
F654
F6FD
F838
F887
F79B
F6D1
F75A
F87C
F867
F6C9
F607
F933
0092
08A2
0D17
0CD7
0A9C
09B6
0AAE
0B88
0ADE
09B5
09DC
0B40
0C13
0B59
0A19
09AA
09FA
0A53
0ADE
0C4D
0E47
0F6A
0F0C
0E20
0DE5
0E49
0E64
0E17
0E35
0EFB
0F7F
0F19
0E69
0E51
0EA3
0EB5
0E98
0ECE
0F24
0ED9
0DE6
0D46
0D96
0E2A
0E22
0DD8
0E40
0F23
0F3A
0E3F
0D97
0E27
0EC9
0E18
0CE2
0D38
0F26
1022
0E55
0B58
0A46
0B64
0B39
0689
FE54
F6F2
F3AD
F416
F578
F5DC
F562
F53B
F5FF
F705
F750
F6C5
F63A
F657
F6D2
F6FF
F6C1
F688
F68A
F669
F5E9
F588
F5EC
F6C8
F70E
F658
F589
F5A2
F679
F70F
F6D8
F62B
F5A4
F596
F606
F6BF
F762
F7A4
F7A4
F7BF
F801
F801
F78F
F739
F7A3
F87A
F8D0
F881
F87B
F935
F9C5
F933
F811
F7C8
F88D
F91F
F8C4
F874
F947
FA64
F9F5
F850
F8C7
FE40
0761
0F56
1273
1156
0F61
0EEB
0F92
0FD4
0F54
0EFB
0F4A
0F62
0E3E
0C48
0B06
0B34
0BE1
0BC2
0ADA
0A46
0A88
0ACC
0A2D
0916
08BA
095A
0A09
0A25
0A27
0A95
0B05
0AD9
0A58
0A3F
0A8A
0A88
0A0F
09DB
0A65
0B07
0ADA
0A0C
0996
09C2
09E5
09A8
0993
09E4
09F3
095E
08F2
0982
0A8B
0B12
0B65
0CAD
0EB6
0F92
0E4A
0CBC
0D47
0ED9
0D57
06A6
FDCD
F7D7
F68E
F7A8
F852
F7EB
F743
F6D8
F69D
F6A8
F722
F7B3
F7C4
F768
F749
F78F
F791
F716
F710
F84C
F9FE
FA84
F95B
F7AD
F6DB
F731
F803
F899
F8B3
F87E
F83B
F7F9
F799
F6FC
F644
F5D9
F604
F691
F6FC
F720
F74C
F7B4
F818
F834
F812
F7BE
F73C
F6E1
F727
F7D4
F7FA
F73E
F682
F6AD
F73C
F6FE
F61A
F627
F7B8
F8E2
F7D0
F637
F846
FF63
07A8
0BEE
0B47
0921
08BD
0A3E
0C0D
0D63
0E77
0F3B
0F3F
0EB7
0E8D
0F12
0F7F
0F43
0EF2
0F4B
0FE5
0FCC
0EF4
0E3B
0E26
0E67
0EA0
0EE8
0F61
0FBF
0F91
0ECD
0DF3
0D8D
0DB7
0E21
0E6D
0E7D
0E94
0F1A
100A
1095
0FE8
0E67
0D86
0E16
0F3F
0F8B
0E74
0C8E
0AB7
0993
095B
09A0
0985
08BD
0820
089C
09A2
0981
07D0
0686
075C
0896
0648
FF6F
F7FB
F49E
F5A8
F77F
F767
F603
F545
F58E
F5DD
F5B9
F5B6
F62C
F69E
F6A7
F6A0
F6DA
F6FE
F6D1
F6D6
F769
F7D2
F730
F5FB
F598
F692
F7F1
F889
F848
F7F7
F81A
F873
F88D
F852
F7FD
F7BA
F7A1
F7CD
F837
F8A4
F8E3
F8F8
F8E1
F88B
F821
F7FB
F810
F801
F7CD
F7E5
F845
F84E
F7D8
F7B8
F883
F96D
F949
F873
F885
F9C4
FA46
F8F7
F880
FCE0
05C9
0DAB
0FA8
0CD3
0A05
09CE
0AAC
0AA9
0A34
0AA1
0B96
0BA8
0AD2
0A8A
0B49
0B9C
0A6F
08E3
08AF
09B4
0A75
0A61
0A36
0A71
0A96
0A44
09ED
0A14
0A6B
0A4D
09C3
097E
09C2
0A01
09C2
096B
09A1
0A2B
0A32
0968
0883
0884
09C9
0BC5
0D65
0DF9
0DCC
0DB6
0E01
0E35
0E02
0DC5
0DE8
0E44
0E83
0EAF
0EE8
0ED5
0E28
0D8B
0E1E
0F4D
0E25
0849
FF7C
F8A6
F6AF
F7BA
F831
F72C
F66D
F704
F7E9
F7F0
F782
F79F
F823
F82E
F7BF
F7C7
F889
F907
F88F
F7D0
F7B3
F7E4
F78D
F6C9
F669
F699
F6B8
F67A
F646
F678
F6D8
F70D
F725
F75F
F79E
F788
F710
F69D
F674
F67E
F6AD
F720
F7A5
F7AF
F72F
F6DB
F723
F780
F74C
F6BA
F67F
F6DD
F79D
F87F
F92C
F918
F812
F6EC
F6C5
F77E
F7C7
F77E
F91E
FF32
0844
0F49
10E3
0EE5
0D8E
0E80
1007
1074
1030
1049
10A7
1094
102C
1016
1020
0F4E
0D9D
0C8E
0D48
0EF3
0FCF
0F52
0E5E
0DDC
0DF4
0E68
0EDF
0EEE
0E6E
0DCC
0D96
0DD5
0E21
0E40
0E5D
0E94
0EB7
0EB0
0EC7
0EFC
0E6D
0C3C
0926
0730
0756
086E
08EC
08D0
0905
09A3
09E8
0994
0945
0960
0988
095E
093C
099B
0A2E
0A46
09F0
09D2
09E9
096D
0855
07E6
08E7
0A3D
0A4A
0923
084E
0894
092A
0912
0872
0825
0878
08DD
08D4
088A
0867
0871
0868
082C
07E7
0810
094C
0BA6
0DDD
0E66
0D73
0CE7
0D7C
0CF9
0892
00AD
F91F
F554
F527
F601
F62F
F61D
F697
F74C
F792
F77C
F765
F718
F65C
F5C2
F603
F6D1
F72A
F6B5
F616
F5F8
F650
F6B4
F6FE
F733
F739
F70A
F708
F78F
F835
F827
F766
F6F0
F746
F796
F6FA
F5EA
F58E
F60A
F667
F60C
F58B
F5AE
F64B
F686
F60A
F571
F565
F5D2
F633
F660
F698
F702
F76F
F791
F73F
F6B0
F66E
F6DD
F790
F7A3
F6E8
F63B
F668
F715
F74D
F6D8
F66F
F6A7
F725
F739
F6D7
F68C
F697
F6B4
F6C4
F6F6
F739
F73E
F736
F7D0
F906
F9C3
F969
F8E4
F956
FA44
FA33
F919
F8BD
F9F9
FAEC
F98B
F785
F96D
0129
0ADE
10DB
1198
1056
105B
117D
11CB
10D3
0FEA
0FDF
1003
0FA8
0F4C
0F99
1018
0FE5
0F25
0ECB
0F17
0F42
0ECE
0E4C
0E6B
0EDF
0EDF
0E56
0DF5
0DF7
0D9B
0C47
0A9C
09D0
0A15
0A67
09FB
0944
0931
09D3
0A66
0A6E
0A46
0A5F
0A7B
0A1A
0962
0913
0978
09F5
09DC
095B
092C
0978
099F
0920
0845
07A3
0757
0725
0721
07A9
089A
091D
08A6
07C8
078E
0820
089E
0863
07D7
07A5
07BA
07A8
07C6
090C
0BA2
0E27
0F09
0E43
0D32
0CDF
0D15
0D3B
0D3E
0D40
0D15
0CB7
0CBD
0D97
0E82
0E3E
0D0C
0CC6
0E05
0E03
0913
FF7F
F669
F2CA
F46D
F6FE
F758
F63B
F5DA
F679
F6AA
F5E6
F54A
F5A8
F651
F65F
F631
F696
F748
F751
F6AD
F666
F6FF
F7AF
F788
F6C6
F653
F66C
F66E
F608
F5C5
F622
F6AE
F6A1
F5F1
F535
F4D2
F4C5
F524
F61B
F76D
F856
F83E
F754
F653
F5D6
F5F0
F655
F6B1
F6CC
F69B
F64A
F619
F617
F619
F610
F620
F650
F65E
F623
F5DA
F5D1
F5FF
F63A
F67A
F6CB
F712
F737
F75A
F7AA
F814
F84E
F841
F826
F82E
F837
F81E
F826
F88F
F8F4
F8AD
F7E2
F789
F813
F8CE
F8FE
F8CA
F89B
F847
F799
F725
F787
F80C
F76F
F672
F86A
FFA2
0991
1089
11A6
0F92
0E91
0F7C
101A
0F43
0E6F
0F1A
107A
10C9
0FD6
0F09
0F30
0F75
0EC3
0D40
0BC4
0AAC
09EB
09A1
09D7
0A08
09BA
0940
093F
09A2
09BE
0954
08DC
08C1
08D8
08CD
08BF
08F9
0953
0953
08FA
08D4
0918
0944
08F9
088C
0872
0898
08CF
0940
09E8
0A2E
09A4
08E1
08D1
0953
094E
0859
078D
080F
0947
098A
088B
080C
098B
0C2C
0DD1
0DB6
0D0C
0D31
0E2E
0F07
0EF2
0E12
0D33
0CFE
0D60
0DC1
0DC8
0DA9
0DA7
0D92
0D09
0C45
0C15
0CCA
0D8F
0D86
0D2C
0D91
0E5A
0E0F
0CB5
0C5A
0DD6
0E56
0A10
014E
F8F3
F569
F632
F783
F72E
F64F
F662
F6DE
F697
F5D9
F5A2
F5BE
F535
F423
F3B8
F467
F53D
F55B
F51E
F545
F5A4
F57A
F4CA
F470
F4C4
F51B
F4F9
F4DB
F53F
F5AC
F58B
F549
F5AA
F662
F661
F56B
F47B
F470
F4FB
F55C
F591
F62A
F713
F763
F6A9
F5B2
F580
F603
F674
F67E
F67F
F6BD
F712
F750
F784
F7B9
F7E0
F7F3
F810
F84A
F88C
F8A5
F87F
F830
F7DF
F7A3
F78C
F796
F7A1
F78F
F77D
F7A7
F7F3
F807
F7CA
F786
F76F
F784
F7E3
F8A6
F94D
F8FF
F7D0
F713
F7B3
F8BE
F894
F770
F763
F928
FA4F
F874
F5B1
F76F
FFCC
0A40
105C
10B3
0F17
0EC7
0EDB
0D19
0A1A
0894
0965
0A78
0A03
08FD
0941
0A9D
0B52
0AC6
0A11
0A0F
0A3C
09D5
091D
08CA
08EF
0913
0921
097B
0A15
0A51
09F7
09A8
09DB
09FF
0961
086B
0832
08E8
098E
095A
08A7
084C
0866
086B
0828
081F
08A2
0917
08BE
07F6
0826
0A15
0CCF
0E89
0E84
0DB0
0D6D
0DED
0E30
0D8F
0CB4
0CA9
0D50
0D88
0CDD
0C37
0C85
0D5B
0D93
0CFD
0C9D
0D29
0DFE
0DFD
0D1B
0C5C
0C66
0CE3
0D47
0D8C
0DC7
0DCE
0DA9
0DCC
0E48
0E68
0DB6
0CE8
0CEE
0D61
0CF1
0BB2
0B8A
0D3F
0DE7
095C
FFA2
F61C
F225
F392
F5D6
F5C2
F45C
F423
F56A
F679
F651
F5B9
F5A9
F5E5
F5B8
F52C
F4CB
F4AF
F4A0
F4B8
F530
F5B2
F5AB
F535
F503
F560
F5B7
F576
F4EB
F4E7
F59B
F64D
F647
F5AF
F53A
F553
F5D4
F656
F686
F64E
F600
F615
F690
F6ED
F6D9
F6C3
F742
F82F
F8C3
F893
F810
F7E5
F821
F846
F819
F7ED
F810
F855
F86A
F845
F817
F806
F832
F8AB
F923
F913
F871
F7EB
F818
F8AC
F8E5
F89A
F856
F879
F8A1
F851
F7CE
F7CD
F862
F8E2
F8DA
F894
F86A
F84E
F841
F896
F93C
F96E
F8BC
F7CA
F75C
F700
F5D7
F4C7
F698
FCCF
04FF
0A8F
0B6A
09C0
08CC
0934
097F
08FC
08A0
092A
09EA
09D1
08E8
0823
0823
08B1
0950
09C3
09F3
09D5
09A3
09BC
0A11
0A10
0991
0937
0983
0A00
09EE
095E
090B
093F
0978
0935
0892
0804
07D3
082B
095B
0B6F
0DA6
0EE6
0EF6
0EC0
0F09
0F74
0F3D
0E71
0DD2
0DD4
0E37
0E8B
0E95
0E4C
0DCE
0D7A
0DB4
0E60
0ED1
0E86
0DCB
0D68
0D95
0DCB
0D9F
0D4D
0D35
0D40
0D36
0D39
0D78
0DBF
0DBC
0D8A
0D7B
0D8A
0D5B
0CD4
0C60
0C6F
0CEF
0D61
0D46
0C57
0A97
08A2
0796
07F3
08A9
0849
0738
0778
096E
0A1B
0604
FDAD
F5CC
F287
F375
F504
F4F7
F437
F463
F53F
F565
F485
F3AC
F3AE
F443
F4C9
F4FE
F4EC
F4A8
F46B
F48F
F522
F5B0
F5BC
F55A
F50F
F520
F550
F56D
F5A9
F627
F687
F660
F5E8
F5C7
F645
F708
F77E
F76E
F70C
F6C4
F6D6
F715
F719
F6C5
F67C
F6A7
F725
F769
F73F
F71D
F781
F81A
F825
F788
F70A
F73F
F7C4
F7EB
F7B3
F79C
F7CC
F7F5
F7F1
F7FF
F83A
F857
F81A
F7CD
F7DB
F814
F7EA
F75C
F721
F79C
F834
F82D
F7B8
F7A2
F822
F88B
F836
F74F
F680
F62D
F639
F686
F76F
F99F
FD62
0203
05D4
0735
0613
0471
04EE
084A
0CB0
0FA5
1054
0FC3
0F39
0F0A
0EE8
0EA5
0E53
0DF9
0DA0
0D8F
0E0C
0ECD
0F1F
0EBF
0E3E
0E36
0E78
0E62
0DE2
0D99
0DF9
0EA2
0EDB
0E64
0DA5
0D24
0CFC
0CF9
0D01
0D31
0DA6
0E47
0ED1
0EF7
0E93
0DCB
0D11
0CD3
0D25
0DAE
0DF6
0DCC
0D78
0D6D
0DA7
0D5E
0BA9
0890
0550
034F
02E0
0334
0363
0344
031C
02F2
0298
023B
025A
02FA
0373
0347
02D6
02D5
0348
0380
031F
0293
026E
029A
02A9
02A3
02FF
03C0
0424
0393
0281
01ED
0239
02DD
033A
033D
0330
0332
0334
033B
035D
0388
0399
03A9
03FB
0466
042F
02F5
0195
01BF
0453
0852
0BA6
0CF0
0C83
0BBD
0B8C
0BCB
0BF2
0BF5
0C42
0CF5
0D77
0D26
0C21
0B41
0B27
0B9C
0BF6
0BFE
0C07
0C43
0C6E
0C49
0C10
0C24
0C65
0C55
0BCE
0B4E
0B60
0BEB
0C53
0C34
0BCD
0BA2
0BE2
0C47
0C56
0BD4
0B0C
0AB4
0B3C
0C1F
0C54
0B8E
0AC6
0B0B
0BE3
0B88
08ED
0525
0258
0180
01B1
0197
0106
00AD
00D4
0114
0121
013A
01A0
020B
01FC
016E
00E0
00BB
00E7
0111
0124
014A
018E
01BD
01A3
014E
00FA
00DF
0110
0174
01D4
020A
0216
0209
01FC
01FE
01FE
01D1
016E
0126
015F
0203
0279
0249
01B4
0156
014E
012C
00F1
01A9
0451
0844
0B77
0C92
0C2F
0BB4
0B8A
0B23
0A67
0A1B
0AB4
0B7A
0B78
0ADE
0AAE
0B27
0B62
0ABC
09E2
09D0
0A5F
0A8F
0A16
09B7
0A12
0AB8
0ADB
0A72
0A21
0A33
0A41
09FC
09B2
09CB
0A12
0A0D
09C9
09C3
0A16
0A47
09FB
097F
0961
09AA
09E7
09EA
0A12
0A8A
0A86
08C8
052C
0154
FF4C
FF8E
00A5
00DF
000E
FF54
FF71
FFDE
FFBB
FF30
FF27
FFE1
007B
0030
FF6C
FF33
FFC0
005B
0069
0023
0010
0043
005C
002E
FFE7
FFB6
FF9B
FFA6
FFF4
0054
005E
0013
FFFC
0054
0086
FFFB
FF19
FEDA
FF6A
FFDE
FF8C
FF11
FF60
002C
0037
FF4E
FF26
016A
0587
091B
0A81
0A33
09B1
09A8
09B8
0976
0916
08F5
0905
08FD
08D6
08C5
08D6
08DD
08D0
08D4
08FB
0921
0924
0916
0919
0928
091D
08F4
08D7
08D9
08C4
085A
07C2
077C
07CA
0852
0880
0841
0810
083F
088B
0891
086E
0890
08EF
08EE
0854
07E8
0876
0955
08AA
0593
017D
FECA
FE5C
FF08
FF57
FF1E
FF0E
FF47
FF2C
FE78
FDCE
FDD1
FE45
FE77
FE4C
FE4A
FEBE
FF4C
FF88
FF7B
FF6C
FF5F
FF21
FEC0
FE93
FEBE
FEF6
FEF2
FEDB
FF0D
FF7A
FFAF
FF71
FF15
FF08
FF46
FF74
FF68
FF51
FF4A
FF20
FEA9
FE3D
FE61
FEFA
FF33
FE99
FE16
FF4A
02AE
06B4
092A
0956
0874
080D
085C
0887
0819
07A1
07CF
0870
08BF
0867
07E2
07C4
0818
0877
0891
0869
082B
07F9
07DC
07D2
07C9
07B6
07A8
07B9
07D3
07BC
0767
0723
073F
0797
07B3
075A
06E0
06B5
06DF
0700
06E4
06C4
06E3
0726
073B
072D
0763
07DC
07AE
05B5
0200
FE32
FC34
FC74
FD9E
FE23
FDBC
FD45
FD5F
FDB6
FDB4
FD61
FD45
FD96
FDF5
FDFF
FDC6
FD9B
FD91
FD7F
FD52
FD28
FD0E
FCEE
FCCD
FCE0
FD3E
FDB0
FDF1
FE08
FE21
FE2F
FDFA
FD88
FD34
FD42
FD7E
FD89
FD59
FD34
FD36
FD33
FD16
FD19
FD4F
FD4D
FCBE
FC3B
FD1A
0005
03FE
0713
081F
07A9
070A
06FE
0745
075F
0738
0712
0707
06F5
06CC
06A2
0685
0663
0633
0624
0665
06D5
071E
0716
06F6
06FB
0716
070A
06DC
06CD
06EC
06F0
06A4
063C
0614
0629
0628
05F8
05E7
062B
067C
067F
0663
06A3
0731
0767
06FC
069B
06F1
0759
0634
02DB
FEBB
FC14
FBB2
FC6A
FCBF
FC71
FC35
FC64
FC9E
FC97
FC8D
FCCC
FD1D
FD1D
FCEA
FD00
FD7D
FDE4
FDC9
FD6A
FD4C
FD78
FD7B
FD23
FCCC
FCD2
FD09
FD0B
FCD7
FCCB
FCFB
FD0B
FCC4
FC7E
FCAA
FD16
FD32
FCE9
FCCF
FD3C
FDAA
FD6C
FCB6
FC68
FCB9
FCCE
FC18
FBA4
FD36
0110
0532
074C
0713
0635
062B
06C7
06FE
068E
062F
0666
06D4
06DA
067B
063A
0649
0655
061A
05CE
05D2
061B
0649
062C
05FB
05F4
0602
05F2
05CC
05C6
05ED
060D
05FD
05D7
05C8
05CB
05B8
058E
0575
057E
058A
0588
059C
05CF
05D3
056D
0502
0549
061D
0616
03DB
FFE1
FC54
FB07
FBB1
FC90
FC7E
FBE3
FBA1
FBD1
FBE8
FBBD
FBB9
FC13
FC6B
FC60
FC22
FC26
FC69
FC82
FC4E
FC38
FC8C
FCF9
FCF1
FC76
FC0F
FC17
FC58
FC6F
FC4C
FC28
FC28
FC3B
FC44
FC3D
FC2A
FC10
FC05
FC20
FC46
FC29
FBB6
FB62
FBB1
FC6F
FCB7
FC08
FB2A
FBB6
FE78
026A
0582
068F
0625
05B3
05ED
065B
0649
05C1
0568
0593
05EA
05F0
05AA
057C
058F
05A4
058A
0564
056D
0597
05A9
0596
0585
0587
0582
0563
0546
054B
055E
0556
0532
0518
051B
052A
0542
0572
05AB
05B0
0577
0555
0588
05CC
05A9
053F
0547
05FF
0659
04CB
0117
FCF6
FA94
FA8C
FB95
FC10
FB9D
FB08
FB09
FB75
FBA1
FB44
FAC7
FAB8
FB24
FB95
FBA8
FB6D
FB41
FB54
FB75
FB61
FB22
FB07
FB3C
FB8E
FBA5
FB74
FB39
FB2C
FB3F
FB38
FB0B
FAEE
FB13
FB5C
FB75
FB3D
FB03
FB1E
FB72
FB8A
FB40
FB0E
FB6E
FC03
FBDE
FADA
FA5E
FC26
0033
0460
0668
0610
0507
04D5
0562
05A3
0531
04A6
04AB
051E
0572
0571
0556
054F
0540
0507
04BD
0493
0498
04C4
0508
0545
0543
04EA
0473
0441
046F
04B4
04C8
04B8
04BB
04C4
0497
043A
0413
0462
04D4
04E1
0486
044C
0488
04D7
04B6
045D
0487
0530
0508
02BD
FEC0
FB33
F9DE
FA72
FB2D
FAF9
FA5B
FA58
FAF6
FB5B
FB13
FA9D
FA92
FAD9
FAF2
FACA
FABE
FAED
FB05
FAC9
FA7F
FA8C
FADE
FB0D
FAFA
FAEF
FB13
FB26
FAEA
FA94
FA89
FAC4
FAE7
FAD1
FAC7
FAF8
FB2D
FB1E
FAF0
FAF7
FB2A
FB26
FADD
FAC8
FB29
FB74
FB08
FA6C
FB34
FE3F
0265
0554
05D5
04D2
0419
0465
04FD
04FB
046E
0410
043B
049B
04BE
04A0
0486
0489
0480
0452
041D
0406
0413
0430
044F
046A
046A
0445
0415
0401
040A
040D
0401
0404
0422
0436
0424
0414
043B
0474
0460
03FB
03C1
0409
0467
0432
0392
0380
0462
050A
03BB
002D
FC26
F9C6
F98B
FA3D
FA8A
FA45
F9FC
F9FE
FA1E
FA30
FA4B
FA7E
FAA7
FAAE
FAB9
FAE9
FB11
FAE3
FA69
FA08
FA0F
FA55
FA75
FA59
FA43
FA69
FAA6
FAB4
FA85
FA49
FA35
FA4A
FA6E
FA87
FA84
FA5D
FA1F
F9F9
FA10
FA4B
FA6B
FA65
FA7E
FAD7
FB09
FA8E
F9B4
F9D1
FC16
0015
03D6
058A
0525
0419
03AB
03E8
042A
0426
041A
0435
044F
0440
0428
0437
044F
042D
03D2
0390
0394
03AC
0394
035E
035F
03B3
0417
0433
03FE
03B3
038C
0389
0381
0369
036A
03A9
040B
043E
0415
03BC
037E
0374
0373
0361
035E
0385
03B9
03C7
03C1
03D2
03DD
039F
0348
0375
042F
0442
023D
FE44
FA66
F8BA
F94B
FA5B
FA7C
F9E9
F9A5
F9EE
FA21
F9D7
F971
F972
F9C5
F9F6
F9E0
F9C8
F9E7
FA1C
FA31
FA25
FA13
F9FA
F9CA
F9A1
F9AD
F9E3
F9FF
F9E5
F9CD
F9FD
FA64
FAA4
FA80
FA2B
FA0B
FA39
FA5B
FA1F
F9B4
F98D
F9C8
FA05
F9FA
F9E2
FA22
FA8D
FA81
F9E1
F979
FA00
FAE4
FAE6
FA01
F9F6
FC60
0089
03ED
04E1
041B
0371
03A6
040D
03F8
03AE
03BC
0403
040B
03D5
03CC
040E
043C
0417
03D7
03C0
03B7
0384
0343
034A
03A2
03E2
03BF
036E
034E
0362
0369
034A
032A
032A
0340
0359
0367
0362
0345
031F
0303
02FC
030F
0342
0384
03A6
037C
032D
031C
035F
0378
0301
027D
02CB
03B0
037C
00DD
FCA8
F94A
F852
F91A
F9EF
FA07
F9D7
F9D5
F9C3
F952
F8DA
F8E3
F95A
F9B0
F9A4
F97C
F978
F980
F96F
F95B
F978
F9C5
FA0C
FA28
FA1A
F9F4
F9BA
F97E
F95B
F950
F946
F943
F96A
F9B0
F9CC
F997
F94D
F93E
F966
F993
F9B6
F9DD
F9FF
FA02
F9F8
FA0C
FA2C
FA0A
F9A5
F985
F9F5
FA50
F9C0
F8D0
F95F
FC83
00E5
0400
04B5
0417
03B0
03D2
03D9
0390
0370
03B7
03EF
03B6
035C
035E
039C
039A
0353
0332
0362
038C
036C
0333
0337
0374
039F
0391
0373
0377
0395
03A8
039E
0376
0332
02EC
02D1
02D5
02C0
028D
0281
02BC
02F7
02EF
02D8
0303
0351
0351
02F8
02CB
0312
034C
02F7
028C
02F0
03CE
035E
006B
FC16
F8DD
F80A
F8C0
F967
F966
F927
F914
F915
F90A
F913
F93E
F954
F939
F930
F969
F9A0
F986
F94F
F969
F9D0
FA10
F9F2
F9C1
F9D4
FA14
FA21
F9E3
F99F
F995
F9B1
F9C3
F9C2
F9C2
F9C9
F9E3
FA17
FA3F
FA1B
F9BA
F981
F996
F9A2
F959
F911
F950
F9F7
FA3E
F9D4
F960
F992
F9FA
F9AC
F8F4
F990
FC97
00CB
03B5
0436
035C
02CA
0300
0368
0382
0367
0355
034B
0336
032E
0342
0345
0322
030F
0337
0365
0352
0318
0309
032F
034A
033A
0326
0334
0348
0339
0313
0302
0307
0301
02F4
030C
0343
035D
034A
0340
034C
0333
02F2
02EE
0350
038F
0326
0278
0272
0329
0394
0308
0264
02E5
03F4
034A
FFC4
FB2B
F866
F859
F967
F9C5
F957
F90B
F93A
F968
F947
F92A
F95F
F9A8
F9A9
F982
F980
F995
F977
F92C
F905
F921
F951
F976
F99C
F9BE
F9B7
F979
F938
F924
F929
F917
F8FB
F91F
F98D
F9E7
F9D9
F986
F94E
F963
F9AE
F9F4
F9EC
F978
F8ED
F8D8
F94A
F99F
F958
F8E9
F933
FA26
FA85
F993
F892
F9B0
FD63
0198
03E5
03F2
0338
02F1
0310
031C
0318
033E
036B
0350
0303
02E8
0312
0322
02F8
02EE
0342
0391
036B
02FE
02C8
02E3
02FE
02F4
02F3
0311
031C
02F7
02DB
0301
0332
0311
02B8
02AA
030C
0367
0356
0311
02FA
0301
02E6
02B9
02B7
02C9
02A8
0265
0260
029D
029B
022E
0209
02CA
0396
028E
FF14
FAE7
F86A
F833
F8E7
F92C
F8F7
F8ED
F937
F970
F95E
F932
F919
F8FB
F8D7
F8E5
F933
F969
F93F
F8F2
F8E9
F91E
F93D
F929
F913
F91E
F93C
F95E
F986
F99F
F980
F92C
F8F2
F910
F94E
F94E
F920
F92E
F980
F99D
F952
F916
F955
F9BF
F9C9
F982
F96A
F997
F99C
F960
F96B
F9FA
FA55
F9C8
F92C
FA61
FDEC
01E7
03F7
03C8
02F2
02BE
02FC
02F8
02B6
02B9
0318
0365
0370
037F
03B0
03A9
0336
02C3
02C8
031B
0335
02F8
02BF
02C6
02F1
0316
032E
0335
0322
0302
02FC
0315
0316
02DD
02AA
02C0
02EF
02CC
027B
0292
0327
0381
0327
0298
0284
02C1
02A9
023F
0238
02C0
030C
029B
023B
02DB
03A1
0263
FE7D
FA20
F7FD
F852
F930
F927
F8A2
F894
F8EE
F900
F8B2
F896
F8DB
F903
F8CC
F8B4
F921
F9A6
F99E
F92E
F904
F950
F996
F97F
F943
F936
F94E
F953
F943
F951
F987
F9B2
F9AA
F985
F962
F945
F939
F955
F97A
F96D
F941
F950
F99C
F9AD
F94D
F8FB
F92B
F97F
F953
F8D9
F8FB
F9DD
FA53
F989
F8BD
FA2F
FE30
0257
0426
03BB
030B
0336
03A2
0384
0316
02FB
0329
0326
02F3
0304
0355
0352
02CE
0272
02BC
0335
032A
02BE
0292
02C1
02D2
02A2
02A1
030A
0367
032F
0295
0242
026B
02A0
0294
0289
02BB
02ED
02DA
02B9
02D2
02FC
02E8
02AC
028F
0288
0260
023A
026F
02DD
02E0
0258
021D
02CA
0346
019D
FD97
F98B
F7EF
F8AF
F9BE
F9BC
F928
F906
F95B
F97D
F938
F8FB
F90A
F923
F916
F921
F96D
F9A6
F97A
F91F
F8F6
F8F7
F8ED
F8F3
F93B
F992
F98C
F92F
F8F7
F92F
F988
F99B
F97F
F98C
F9B2
F98C
F921
F8FC
F950
F99F
F982
F949
F962
F99A
F97F
F932
F930
F976
F980
F936
F934
F9B6
F9F1
F941
F8C2
FA7B
FEA7
02C9
044F
0362
024A
0277
033C
0363
02EF
02B8
02FB
0326
02E2
02A2
02D1
0328
0331
0303
0301
032B
0334
030D
02E9
02CD
029A
0261
025F
0295
02B5
028F
0256
024E
0265
025A
023B
0256
02AA
02D4
02B5
02AA
02E9
0316
02E3
0298
02A1
02D7
02CE
028F
0290
02CF
02BC
0236
020C
02C6
0338
0173
FD59
F95A
F7DB
F8A2
F987
F943
F890
F88E
F921
F962
F914
F8D9
F91A
F970
F95F
F913
F8FD
F91D
F920
F8F8
F8DD
F8E3
F8EE
F8FE
F928
F956
F958
F937
F938
F979
F9BD
F9C1
F994
F977
F970
F953
F92D
F943
F98C
F99E
F951
F911
F938
F983
F988
F95D
F95F
F980
F961
F910
F91A
F993
F9B2
F90D
F8D9
FAE5
FF20
030E
0462
037C
0295
02E1
0387
035C
029C
0256
02C9
0328
02E5
0280
02A7
0332
0370
0330
02DE
02CC
02D9
02D3
02CA
02DE
0301
030B
02ED
02B4
0273
0237
0213
021D
0259
02A7
02E5
02FB
02E3
02AF
0297
02CC
0329
0350
0326
02ED
02D5
02BF
02A0
02B2
0302
0316
0281
01C5
01EB
02EB
0310
00B2
FC7A
F908
F822
F8F0
F97E
F933
F8FB
F96C
F9D4
F968
F88F
F84E
F8D2
F945
F918
F8BE
F8CF
F91F
F920
F8DA
F8D2
F932
F98D
F992
F96F
F968
F965
F930
F8F3
F90F
F97D
F9C2
F98C
F929
F910
F93F
F95E
F951
F94D
F964
F95D
F91A
F8E7
F91C
F996
F9B9
F93C
F8D1
F9BC
FC8F
0056
033C
0419
0366
029E
02B4
0355
039D
034C
02EE
02F7
0330
032D
02FB
02F2
0321
0336
0306
02CF
02D4
02F9
02F2
02C1
02A7
02C0
02D9
02D5
02D4
02E7
02E5
02BE
02B5
02FE
034A
031F
028E
022E
0259
02B9
02D1
02B3
02C3
02EE
02BF
0244
0243
0307
0371
01EA
FE55
FA7B
F851
F82A
F8D7
F938
F933
F932
F94F
F955
F937
F923
F91A
F8F2
F8AE
F899
F8D9
F92C
F936
F8FA
F8D0
F8EE
F92F
F956
F962
F973
F981
F961
F91C
F8FB
F927
F963
F955
F901
F8CB
F8F5
F944
F953
F91E
F900
F92E
F971
F98C
F9AA
FA08
FA56
F9EF
F8F6
F8CA
FACA
FEA5
024B
03DD
036D
028E
0270
02E1
0324
0315
0316
0341
033F
02F4
02C0
02EF
0341
0346
030E
030B
0360
03A0
0370
0304
02C9
02CD
02D0
02C3
02DC
0327
0354
0332
0304
0323
0373
0380
032D
02E6
02FE
0334
031C
02CD
02B9
02E5
02CC
023E
01E7
027C
036D
030E
005E
FC61
F951
F875
F918
F9B2
F994
F932
F919
F92F
F91D
F8F2
F903
F952
F981
F965
F946
F96A
F99F
F98A
F93C
F925
F96D
F9B0
F991
F93E
F921
F944
F952
F92D
F91D
F94E
F973
F93C
F8DC
F8D2
F925
F954
F925
F904
F952
F9B3
F98F
F915
F917
F9C6
FA2E
F985
F8A6
F97E
FCBC
00C0
033B
0388
02F1
02D5
033D
036C
032C
02F5
030E
0322
02E3
02A0
02D1
0354
0391
034D
02FE
0319
036B
0364
02E6
026A
025B
0297
02B9
02A6
029D
02B9
02D1
02C8
02D0
0317
0369
0370
0331
030A
0323
0333
0305
02D7
02FF
0343
0315
028A
027E
0352
03D8
024B
FE80
FA7D
F87F
F8B0
F964
F953
F8DD
F8F6
F98F
F9C1
F93F
F8C9
F900
F97F
F988
F92A
F91B
F991
F9EA
F99E
F902
F8D0
F923
F977
F972
F955
F972
F9AD
F9C0
F9B2
F9BC
F9CE
F9AA
F95B
F93A
F965
F985
F951
F90B
F91C
F965
F960
F902
F8F5
F99D
FA3E
F9CD
F895
F86F
FAD9
FF1C
02CD
0430
03B9
0317
0332
038C
0375
0316
0314
037A
03A1
032C
0295
028C
0309
0367
0348
0307
031B
036A
0377
031E
02BD
02A9
02C9
02DE
02E7
02FD
0307
02E5
02BA
02D3
0328
034D
030E
02C1
02CD
0303
02E9
0294
029A
0316
034C
02C1
022C
0299
0395
0323
0000
FB85
F87A
F826
F939
F9B4
F93B
F8DD
F934
F99C
F960
F8CB
F8AB
F91C
F978
F94C
F8EF
F8E0
F919
F93C
F932
F933
F94D
F94A
F91E
F90E
F949
F99C
F9B7
F9A5
F9AC
F9D6
F9D8
F994
F95E
F98F
F9F7
FA17
F9D3
F99B
F9C4
FA03
F9E0
F97C
F96B
F9C7
F9E2
F945
F8CF
FA25
FDC3
0200
0476
045E
031F
0282
02DF
034E
033A
0310
035D
03E3
03F3
037C
031D
033D
038A
0393
0372
0384
03C2
03CA
0382
0342
0348
035D
0337
02FD
0304
0331
0313
02A2
026C
02C9
0348
0343
02CF
028F
02BB
02DD
029B
024D
0266
02A2
026C
01F3
0222
031F
037A
0192
FDB1
FA0D
F88F
F901
F9BE
F9B5
F93F
F91B
F94E
F961
F934
F923
F954
F979
F949
F8F3
F8CE
F8DC
F8DA
F8BA
F8B7
F8F6
F93C
F942
F923
F939
F999
F9ED
F9ED
F9BA
F99B
F995
F973
F932
F91E
F962
F9B9
F9CD
F9AC
F9B3
F9F8
FA21
FA01
F9F5
FA53
FAB1
FA4F
F96B
F98E
FBFF
000F
0377
049F
040D
036A
037D
03B3
0371
030D
032D
03AB
03D2
0371
0319
0343
039F
039A
033C
0307
0329
033D
02FB
02B2
02CC
032C
035F
0346
032C
033B
033F
0315
02F9
0327
035F
0334
02B9
0282
02D3
0336
032D
02E1
02D6
02FF
02CE
022E
01EB
029A
035E
0279
FF47
FB48
F8C0
F87A
F948
F9A2
F937
F8C4
F8CB
F902
F8FB
F8D2
F8ED
F955
F9A3
F999
F975
F98B
F9D1
F9FD
F9F6
F9EA
F9F7
F9FF
F9DD
F9A4
F97A
F960
F94A
F949
F977
F9AB
F997
F93D
F90F
F95D
F9D1
F9CE
F954
F915
F983
FA2D
FA61
FA2D
FA35
FA9A
FA9C
F9D8
F960
FAE4
FE92
0280
0483
045B
0395
0384
0400
0426
03BF
035B
0358
036B
033D
0300
031F
0389
03C1
0384
030F
02BD
02A6
02B6
02ED
0345
0381
036C
0330
0332
0382
03AF
0365
02F8
02FF
0381
03DE
03AD
0348
0346
0397
039A
0312
0281
026A
0293
0272
022F
0285
0373
0395
0176
FD71
F9BC
F83D
F8C1
F98C
F976
F8E6
F8CD
F948
F9A6
F97C
F921
F90C
F936
F94F
F94A
F95E
F995
F9BD
F9BD
F9B7
F9C4
F9C7
F9A7
F997
F9C8
FA04
F9DE
F94E
F8E0
F900
F971
F9A9
F997
F9A1
F9EF
FA1E
F9DE
F983
F99A
FA13
FA4B
F9FC
F9B1
F9EE
FA54
FA22
F992
FA0E
FCA5
0089
03A1
049C
0414
038A
03A9
03E5
039E
030B
02D8
033A
03C3
0405
03FD
03DC
03AF
0372
033F
0339
034E
0348
032A
0332
0372
039F
0372
031F
0318
036D
03B0
0393
0355
0357
0385
0379
0328
0302
0340
0376
0326
028C
0259
02B3
02FC
02CD
02AD
032E
03A9
028A
FF36
FB29
F8AC
F887
F979
F9E1
F971
F8FF
F91D
F97F
F9A7
F993
F989
F998
F999
F993
F9B3
F9F1
F9FD
F9AF
F955
F951
F994
F9BC
F99D
F976
F981
F9A6
F9AE
F9A2
F9B2
F9D6
F9D0
F99D
F999
F9FE
FA78
FA7D
FA04
F9A0
F9BF
FA20
FA49
FA44
FA78
FADF
FADB
FA36
F9F1
FB79
FEEE
029D
0496
0484
03B6
036F
03B1
03C5
0376
0334
0345
035C
0324
02D6
02E7
035C
03BE
03C1
0390
0371
035E
0340
033A
0379
03D4
03EB
03B5
038A
03A2
03BB
0381
0323
0312
0355
0373
0330
02F6
0330
0392
0379
02E2
027D
02B3
0308
02E8
02A3
02FC
03BB
035C
00B8
FCAD
F986
F8B0
F97E
FA3C
FA1B
F99B
F976
F9AA
F9C5
F9A9
F9A0
F9D2
FA0C
FA17
F9FF
F9E3
F9C1
F990
F974
F99C
F9E8
FA05
F9D9
F9AB
F9B9
F9E0
F9CE
F98F
F97D
F9B9
F9ED
F9D3
F9AB
F9E0
FA50
FA60
F9DE
F96F
F9B6
FA67
FAA7
FA44
FA01
FA67
FACC
FA3C
F934
F9A0
FCB1
012A
046F
051D
0421
0345
033E
0386
0398
039D
03DA
041F
0410
03C2
0391
0392
038E
0375
037C
03AC
03B8
0376
033D
0377
03FB
042D
03DB
0387
03A7
03F2
03D9
0365
032A
0360
038E
034E
0305
0348
03D9
03D7
0318
02A4
034B
0423
0336
FFDC
FBCC
F96D
F956
FA0F
FA0F
F965
F925
F9BA
FA73
FA89
FA0C
F994
F973
F988
F9AE
F9E7
FA24
FA34
FA12
F9FF
FA22
FA3A
F9FE
F99E
F992
F9F0
FA41
FA29
F9E6
F9E8
FA25
FA2F
F9F7
F9EE
FA48
FA8A
FA3F
F9CF
FA01
FABD
FAEA
FA07
F95C
FAD7
FEA7
02AC
0497
043E
0357
0343
03C2
03E7
038F
036A
03CF
0447
044E
0406
03E8
0407
0413
03E6
03B2
039A
0385
0368
0378
03D1
041E
03F7
0385
035D
03B2
0404
03D4
0361
0341
037E
039A
0363
0356
03C3
041A
03A2
02C1
02B3
03BA
042E
0230
FE0F
FA51
F90E
F9DF
FABE
FA86
F9DE
F9D0
FA4E
FA8B
FA4C
FA1E
FA58
FA94
FA55
F9C5
F96F
F97D
F99E
F9A3
F9B9
F9F8
FA17
F9E4
F9AD
F9D9
FA3F
FA51
F9F5
F9BD
FA14
FA94
FA9E
FA43
FA2E
FA89
FAB6
FA48
F9D2
FA13
FAAE
FA86
F990
F981
FC02
0065
0401
04F4
03F6
0323
036E
0407
03EF
035C
0327
0382
03DC
03D9
03C6
03F3
041E
03EE
0396
0393
03E8
0419
03E8
03BA
03EC
043A
041D
03A2
0365
03AA
03FC
03DF
038B
0387
03D3
03EA
039D
035D
037C
039B
0351
0307
037A
0450
03DE
00FE
FCC6
F9B4
F927
FA1A
FAAB
FA40
F9BC
F9E4
FA59
FA5D
F9F3
F9B6
F9E0
FA0C
F9EF
F9CC
F9F5
FA39
FA32
F9F5
F9FC
FA68
FABC
FA8B
FA13
F9E4
FA15
FA3E
FA1F
F9F6
FA11
FA5E
FA9B
FAB9
FAC7
FA9F
FA19
F98E
F9A7
FA67
FADC
FA50
F99E
FAA0
FE02
0221
048F
0492
0399
0347
03B5
03F2
039D
035B
03B4
044B
047C
0448
0434
0465
0462
03E5
035A
0350
03AF
03E2
03AD
036D
037E
03C3
03E4
03D3
03BC
03AC
0391
0386
03C3
0427
0432
03B9
0344
0362
03CB
03B8
0320
02FF
03E0
049C
0343
FF7E
FB5E
F951
F9A9
FAA0
FA9F
F9D5
F966
F9B0
FA08
F9E8
F9A4
F9C9
FA39
FA6B
FA37
F9FA
F9F5
F9F8
F9CA
F993
F99F
F9E2
FA15
FA22
FA35
FA54
FA48
FA0A
F9F7
FA51
FABE
FAB6
FA43
FA01
FA36
FA6E
FA3C
FA01
FA59
FAF8
FACE
F9B3
F949
FB62
FFAE
03A4
0515
0450
0360
038D
0448
0479
040F
03C4
03E7
040C
03E8
03CA
0402
044C
0438
03E3
03D7
0439
0490
0488
046A
0494
04C2
0467
0397
0314
0354
03DF
0400
03B7
0397
03D0
03ED
03AB
0375
03AF
03F6
03AE
0325
0354
0448
0464
020A
FDC9
FA2A
F910
F9E4
FAAE
FA82
FA24
FA6C
FAFF
FAFB
FA54
F9D7
F9F1
FA2D
FA0C
F9D1
FA05
FA8D
FABD
FA54
F9D8
F9D1
FA18
FA2D
FA06
FA08
FA51
FA80
FA52
FA18
FA3D
FAA8
FAE2
FAD0
FABF
FAD3
FAC9
FA87
FA74
FAD9
FB2A
FAA7
F9C3
FA3B
FD2F
0170
046B
04CF
03C2
0347
03F2
04B7
04A6
0414
03DA
0414
0435
0405
03EC
042C
0467
0432
03C7
03B3
03FF
0420
03C9
0366
037F
03F8
043E
0413
03C8
03AB
03A2
0381
036A
039B
03FA
042D
0423
0415
0404
039F
02F2
02C6
03AD
04BE
0408
00A3
FC17
F90B
F8AB
F9C1
FA6B
FA2B
F9DB
FA20
FA95
FA96
FA3E
FA1D
FA57
FA7D
FA4E
FA14
FA25
FA55
FA44
F9FB
F9E9
FA3D
FA9F
FAAF
FA7E
FA5F
FA68
FA67
FA4A
FA3F
FA64
FA94
FAA9
FAB3
FAC6
FAC0
FA85
FA5E
FAAB
FB35
FB36
FA75
FA15
FBA5
FF42
0319
051A
0500
043E
0421
048F
04B0
0452
040D
0444
0494
0479
0413
03EE
0434
0484
0482
044A
0422
040E
03EF
03D9
0402
045E
0497
0479
0436
0413
0404
03DB
03A5
03A6
03E6
0423
0433
0439
0444
040A
0363
02E9
037A
04DA
054C
0326
FEDA
FAD6
F931
F9B8
FA98
FA8E
F9F9
F9CF
FA34
FA80
FA58
FA17
FA26
FA63
FA6C
FA3A
FA1D
FA34
FA4B
FA3C
FA2D
FA42
FA57
FA36
FA01
FA07
FA55
FAA3
FABB
FABF
FADA
FAF1
FAD8
FAAE
FAB9
FAE1
FAC4
FA60
FA4E
FAE6
FB80
FB1E
F9FE
F9E5
FC52
0091
0429
054D
0481
039E
03AD
042F
0450
040D
03F5
0436
0470
0460
043D
044E
0472
0465
0439
0438
046E
048F
046D
0436
0423
042A
0422
041C
0446
0484
047E
0427
03EF
0428
048B
048F
0431
03F2
0409
040B
03AD
0372
0408
04EA
0467
0170
FD28
F9FD
F948
FA24
FACB
FA8A
FA0E
FA0C
FA51
FA52
FA0D
F9F6
FA34
FA6B
FA50
FA11
FA01
FA1F
FA30
FA2A
FA33
FA52
FA57
FA3D
FA48
FA99
FAE2
FAC2
FA5C
FA35
FA80
FAD0
FAB8
FA63
FA46
FA75
FA96
FA8D
FAB0
FB13
FB1F
FA60
F9A6
FA9D
FDE9
0210
04B3
04EE
03FF
039F
0427
04B3
049A
0438
0436
049C
04F0
04F7
04E5
04E4
04D4
049B
046D
047C
049F
048C
0450
0447
048F
04CD
04AC
0453
0428
043F
0449
0420
03FE
0413
0433
041A
03EA
03F3
041D
03F8
0386
037B
0442
04EF
03D7
007B
FC72
FA01
F9DA
FAAD
FAE2
FA43
F9BD
F9E9
FA6A
FAA3
FA89
FA6F
FA68
FA40
FA04
FA10
FA84
FAF4
FAE0
FA58
F9EC
F9F5
FA47
FA81
FA8B
FA80
FA6E
FA4B
FA2A
FA37
FA72
FAA8
FABB
FAC1
FACE
FABC
FA6D
FA25
FA49
FAB7
FAC7
FA46
FA28
FBC7
FF45
0304
0517
0510
042F
03D8
043C
04A9
04AF
048C
0490
0498
045B
03F3
03D4
0430
04B9
04F5
04C4
045F
040F
03F5
040E
0442
046B
0471
0469
0477
0490
047E
042B
03DA
03DE
042E
046D
0467
0446
0434
0412
03C3
03A3
042A
0505
04D7
0279
FE70
FAC0
F91F
F96D
FA2F
FA49
F9E8
F9C8
FA20
FA81
FA99
FA98
FAC5
FB09
FB1A
FAEF
FAC5
FABB
FAAB
FA6F
FA29
FA15
FA45
FA94
FADC
FB0C
FB0F
FAD3
FA73
FA38
FA4E
FA8D
FAAD
FAA5
FAA3
FABA
FAC8
FAC5
FAE7
FB3C
FB57
FAC6
F9FE
FA66
FD06
012C
04C6
0631
0599
0479
03FB
0421
0456
0454
0449
0458
0466
0460
0464
048A
04B1
04AA
0480
0467
046E
0468
043C
0409
0401
0421
0447
0460
0468
044A
03FA
03AB
03B3
0417
0460
0431
03D8
03F8
0496
04E6
0458
0384
0383
0443
0427
01C0
FDB1
FA50
F94B
FA15
FAE7
FAD3
FA6C
FA82
FAF4
FB0C
FA97
FA1B
FA08
FA36
FA4F
FA5D
FA98
FADD
FACA
FA5E
FA15
FA47
FAB0
FAD4
FAAF
FAAA
FAE8
FB14
FAED
FAC4
FAFF
FB72
FB8B
FB2C
FADD
FAF5
FB09
FAA4
FA61
FB98
FEB0
0241
045A
0485
0403
0415
0497
04A4
041A
03D6
046D
0544
0563
04BA
0423
042F
047B
0465
03F7
03C4
040C
046A
047E
0465
046F
0493
0489
0449
041E
0429
0431
040C
03EF
0415
044F
0441
040D
0439
04B3
045D
021D
FE67
FB21
F9D3
FA2E
FAB4
FA85
FA20
FA4D
FAF5
FB56
FB19
FAAD
FA8C
FAA5
FAAE
FAB2
FAEC
FB44
FB55
FB02
FAAE
FAA9
FAC1
FAA0
FA6B
FA93
FB15
FB5B
FB0A
FA97
FAA8
FB15
FB1B
FA8B
FA36
FAC2
FB88
FB62
FA78
FA94
FD24
0145
047A
0545
047D
03F0
0449
04C5
04B1
045A
0455
048F
047E
0417
03E0
041E
0464
0446
0403
041D
0484
04A3
044B
040B
0457
04C5
049A
03E4
0382
03E8
0481
0486
0420
0410
046A
046D
03C5
0355
0403
0509
0462
0130
FD18
FAA1
FA7B
FB0F
FABD
F9C5
F98B
FA7A
FB79
FB70
FAAB
FA41
FA97
FB0A
FAFD
FAA3
FA87
FABB
FAE3
FAD9
FAD8
FB02
FB20
FB03
FAD7
FAD8
FAE8
FACC
FAB4
FB05
FBA3
FBD0
FB1F
FA3F
FA39
FB02
FB65
FAB4
FA16
FB7D
FF41
036C
05A3
057D
0485
0436
0493
04C6
0487
0456
048D
04DE
04DA
0499
047F
049D
04A4
0474
044C
0465
0492
048E
0466
045E
0479
0475
0442
0429
0455
047F
0450
03FD
040B
0473
0476
03AE
02E7
0353
04C7
055F
035C
FF36
FB54
F9B3
FA1D
FAE7
FAF2
FA84
FA54
FA78
FA83
FA58
FA57
FABA
FB32
FB58
FB2D
FAFA
FAD9
FAA8
FA6E
FA6C
FAB8
FB06
FB09
FADE
FAD8
FAFE
FB03
FACE
FAB7
FAF8
FB36
FAF4
FA68
FA66
FB33
FBF2
FBA7
FAC4
FB16
FDC3
01BC
0494
04F9
03E5
034C
03F4
04F9
053B
04AF
0425
0421
0465
0486
047E
0484
0495
047F
0445
0431
046A
04B6
04C1
0485
0438
0402
03EB
03FB
043C
0480
047C
0430
0417
0488
0513
04EC
0410
038D
042E
051D
046B
0143
FD22
FA75
FA24
FAEF
FB2B
FAA3
FA5A
FADF
FB8E
FB83
FAD2
FA50
FA75
FAE4
FB12
FAFF
FB00
FB1F
FB0E
FAB7
FA70
FA8D
FAE6
FB16
FB08
FAF8
FB0D
FB22
FB1B
FB16
FB29
FB1E
FACC
FA89
FAD1
FB6F
FB7E
FAA2
FA0C
FB83
FF41
0342
0534
04D0
03DB
03E4
04A6
04E5
044B
03C2
0406
04A8
04CD
046A
0434
0482
04DD
04C3
0469
0455
048C
0497
0447
0409
0441
04AF
04CA
047A
042B
042E
045C
047B
0493
04B7
04AC
043C
03CA
03FE
04B4
049D
027A
FEBB
FB5F
FA05
FA69
FB05
FAEB
FA8C
FAAA
FB2C
FB5E
FB0A
FABB
FAE7
FB45
FB47
FAF0
FAC3
FAFF
FB40
FB22
FAD0
FABB
FAFB
FB3F
FB4F
FB46
FB37
FAFD
FA93
FA53
FA96
FB1B
FB4A
FB0F
FAFE
FB68
FBB6
FB42
FAA1
FB6E
FE6B
0249
04C9
0506
042A
03D3
0455
04DD
04DE
04AD
04C3
04F9
04E1
0487
045D
0488
04AA
047A
0434
0432
0455
0437
03DB
03BF
0429
04B1
04CC
0483
045B
0482
0492
0441
03E9
0406
0466
0453
03BA
0376
0421
04D3
03C8
0079
FC84
FA2C
FA14
FAF2
FB4E
FB08
FAE3
FB27
FB51
FB0E
FAC9
FAFE
FB6C
FB6C
FAED
FA91
FAC8
FB36
FB42
FAEB
FAB6
FAE2
FB23
FB30
FB2B
FB53
FB81
FB69
FB27
FB27
FB84
FBD1
FBBF
FB9E
FBD4
FC1D
FBC4
FADF
FAC2
FCBA
006D
03E4
056B
0520
0471
0462
04B3
04A5
0421
03BF
03E3
0443
046B
0459
0466
04AD
04E4
04D3
049F
0487
048B
0482
046D
0476
0497
0495
0458
0426
043B
0463
0443
03F8
03FD
0460
0486
0408
037C
03C1
048A
043A
01AC
FDCB
FAD6
FA18
FAD2
FB79
FB76
FB45
FB50
FB62
FB3F
FB22
FB54
FB94
FB68
FAE1
FA99
FADE
FB3D
FB2B
FACC
FAAC
FAEC
FB1A
FAF4
FAD5
FB20
FB95
FB9E
FB34
FAFB
FB54
FBBB
FB7D
FAD2
FAAF
FB63
FBFF
FB99
FAE0
FBAB
FEBF
029A
04E9
04F6
0423
0402
0496
04D7
0465
03F6
0426
0496
049A
0447
043F
04AB
04F9
04C2
0465
0474
04D6
04F5
04A8
0468
0487
04B9
04A6
0483
04AE
04EA
049F
03E4
039E
044F
052B
0507
0405
0394
0478
055B
0415
0046
FC0C
F9D9
FA0C
FB11
FB75
FB47
FB50
FBAF
FBC3
FB46
FAC6
FAD4
FB34
FB45
FAFB
FAE3
FB39
FB77
FB14
FA5B
FA17
FA8B
FB1E
FB32
FADD
FAA0
FAB1
FAE8
FB36
FBA5
FBEE
FB9B
FAD3
FA88
FB45
FC2E
FBE3
FA85
FA1D
FC70
00B8
0447
055A
04BD
045A
04DE
056A
0538
04AA
047C
04AA
049E
0437
0405
0461
04E2
04EE
0496
046D
04AF
04FE
04FE
04CD
04B6
04B1
0480
042A
0406
0437
0477
0485
0490
04DF
0537
0510
0477
0445
04FF
05C1
04D6
01AA
FDB8
FB2C
FAB9
FB32
FB38
FAB7
FA7C
FACE
FB12
FACE
FA68
FA7B
FAE5
FAFA
FA89
FA2A
FA61
FAE5
FB1D
FAF8
FAF3
FB3F
FB73
FB3B
FAEC
FB10
FB94
FBDD
FBA6
FB57
FB5B
FB84
FB72
FB44
FB6B
FBC9
FB9A
FA9C
F9FE
FB6E
FF1E
0330
056C
0555
0449
03C4
0402
045F
0482
04AA
0501
053B
0519
04E5
0515
0590
05B6
0533
046B
03F3
03E6
03F4
0401
043C
04A9
04EB
04BF
0469
045A
0494
04AD
0482
0468
048D
048F
0417
03A8
0423
055F
05BA
03AB
FFA7
FBF6
FA7F
FB0F
FBF5
FBFC
FB57
FAD1
FAB4
FABB
FABF
FAE2
FB2E
FB59
FB32
FAF5
FB07
FB64
FBA9
FB96
FB5E
FB51
FB73
FB91
FB97
FB9E
FBA9
FB91
FB52
FB2D
FB50
FB81
FB62
FB06
FAF0
FB4A
FB82
FAFF
FA4C
FAED
FDCE
01F7
053D
0648
05A5
04D7
04AE
04D3
04B5
0460
0437
044D
045B
0447
044B
0484
04AD
047F
0424
040A
044A
048C
048C
0470
047B
049C
048B
0450
043F
0478
04A8
0487
0458
0485
04E4
04CD
041E
03AC
0436
0510
0474
0178
FD5A
FA6B
F9CE
FAA0
FB4A
FB35
FAE5
FAE3
FB1D
FB51
FB85
FBD3
FC08
FBDB
FB6C
FB33
FB62
FBA4
FB95
FB45
FB0B
FB03
FB04
FB0A
FB41
FBA7
FBDF
FBA4
FB3C
FB24
FB61
FB83
FB60
FB68
FBF3
FC76
FC0C
FAD3
FA52
FC11
FFD7
03B3
05C6
05D6
050E
048B
0484
04B2
04F8
055A
059A
055C
04B2
0434
0454
04CC
04F1
0492
042A
043C
04A7
04EB
04DD
04CB
04F6
052B
0519
04C4
047B
0467
0470
0489
04C6
0509
04F0
0458
03D9
0439
053C
0565
035B
FF81
FBDD
FA39
FA8B
FB5F
FB84
FB1A
FAEF
FB4D
FBB3
FB9E
FB38
FB0B
FB43
FB84
FB6F
FB1E
FAEF
FB04
FB1D
FB03
FAD0
FAC4
FADD
FAEA
FADE
FAED
FB2B
FB61
FB5A
FB38
FB3B
FB44
FAEE
FA53
FA64
FC29
FF84
030B
0537
05B2
0548
04DE
04B3
049D
048D
04A5
04E4
050D
04F0
04B8
04BD
0514
056A
0568
051B
04E3
04FD
0536
0533
04EB
04BB
04EC
0546
0558
0512
04CE
04C2
04BA
048D
048D
050D
057E
0496
01A9
FDC2
FADA
FA04
FA8E
FB19
FB12
FAE6
FB02
FB3F
FB4C
FB3D
FB62
FBC0
FC02
FBE7
FB98
FB5C
FB36
FAFA
FAA7
FA78
FA8E
FAB7
FAAD
FA77
FA71
FADA
FB71
FBB0
FB69
FB0C
FB0B
FB32
FAE8
FA4F
FAA3
FD0B
010F
04A9
0629
05CA
0529
054F
05C7
05AB
0503
049B
04D2
052B
0511
04A9
047D
04B5
04ED
04CC
0479
0450
0467
0491
04B8
04F1
0535
054C
051D
04E3
04E8
0519
050C
0491
0417
0449
0510
0539
037C
FFEE
FC3B
FA33
FA25
FAD8
FAFD
FA72
F9FB
FA14
FA78
FAB5
FACD
FB02
FB52
FB78
FB61
FB48
FB5F
FB86
FB87
FB64
FB52
FB6D
FB90
FB8D
FB70
FB6D
FB96
FBBB
FBA7
FB5F
FB27
FB24
FB22
FADD
FABC
FBDE
FEF5
0314
061B
06C2
05E4
0560
05EC
0683
060B
04E4
0450
04B5
0534
050E
04A6
04B9
0527
0533
04B6
0463
04B1
0527
0508
0459
03CF
03D2
0410
0423
0429
0465
04A4
047C
0415
042D
0514
05E8
052E
024E
FE59
FB46
FA3C
FAAD
FB22
FACA
FA16
F9DA
FA38
FA99
FA99
FA87
FAD4
FB51
FB74
FB2F
FB0B
FB58
FBAE
FB94
FB41
FB4C
FBC1
FC0E
FBDE
FB98
FBC0
FC27
FC32
FBCA
FB98
FC07
FC84
FC27
FB1C
FAD3
FC9F
0035
03C0
057B
053B
045F
044F
0516
05AF
0571
04D7
04B9
0527
056B
051D
04B3
04CE
0543
055B
04E3
0472
0478
0498
0440
039C
0358
03AC
0422
0455
046F
04AA
04C0
0451
03B9
03DF
04E5
0575
03F4
0058
FC7E
FA6F
FA92
FB98
FC08
FBA8
FB55
FBB5
FC5A
FC64
FBBB
FB35
FB7D
FC2C
FC58
FBCD
FB47
FB69
FBE4
FBF9
FB8C
FB3B
FB64
FBB3
FBD1
FBF5
FC6B
FCE0
FCD1
FC64
FC46
FC96
FC84
FB85
FA82
FB41
FE6A
028B
056B
060F
054A
048B
048E
0514
0579
055E
04F0
049D
04A3
04DB
04FE
04F4
04CB
0494
0460
0458
0494
04EB
0500
04C4
04A2
04EF
054A
0510
045B
0404
046A
04CD
046E
03C8
03F7
04DD
04C2
0247
FE49
FB27
FA48
FAE4
FB6B
FB60
FB54
FBA6
FBF5
FBD8
FB71
FB24
FB13
FB19
FB20
FB33
FB50
FB64
FB67
FB7A
FBAD
FBDF
FBE4
FBBA
FB8F
FB88
FBA2
FBB2
FB83
FB1C
FAE5
FB41
FBE5
FC03
FB62
FB13
FC8B
FFF9
03C6
0605
063F
0592
0542
057A
05A3
056A
0518
0503
0511
04F4
0495
043D
044A
04C9
0557
0582
053E
04ED
04E0
0505
0518
0506
04EF
04E0
04BB
0481
0467
047A
0466
03FC
03BA
0438
04F5
045D
0190
FDBD
FB24
FAC7
FB9E
FC0A
FB96
FAF9
FAD5
FB05
FB28
FB39
FB59
FB73
FB75
FB92
FBF1
FC45
FC1E
FB95
FB41
FB78
FBF0
FC25
FBF5
FBA9
FB85
FB81
FB6A
FB36
FB12
FB32
FB92
FBDC
FBA7
FB2C
FB89
FDD8
01B0
0514
0649
058C
048D
046F
04D2
04D1
045A
0411
0436
0454
0419
03DF
0416
048E
04C6
04BA
04D5
052E
0557
04F9
045F
0416
0435
044D
0412
03CC
03FB
0494
04FA
04C8
0469
04A0
0566
057D
0381
FF94
FBB3
F9F6
FA88
FBA6
FBBA
FAEA
FA70
FAD5
FB84
FBD3
FBE1
FC1E
FC71
FC66
FC01
FBDC
FC44
FCB4
FC8E
FBF3
FB8D
FB99
FBB6
FB9A
FB8A
FBDE
FC59
FC61
FBD7
FB63
FBAD
FC6E
FCA5
FBE7
FB33
FC23
FF32
0302
0583
05D9
04FA
046A
04A5
0505
04F5
04B3
04BF
050B
0524
04E9
04AE
04AA
04AE
048B
046C
0488
04A6
045E
03CA
038F
03FE
0490
0498
043A
0438
04DD
0580
055B
049B
043E
04D4
0591
04E4
020C
FE0A
FADC
F9D0
FA81
FB77
FBA1
FB2B
FAE3
FB20
FB7B
FB8A
FB67
FB5F
FB72
FB71
FB62
FB70
FB89
FB68
FB12
FAFC
FB6F
FBFB
FBEA
FB3C
FAC3
FB0D
FBA8
FBC6
FB68
FB51
FBDC
FC4F
FBCE
FAB3
FA8F
FC97
003A
0384
04EA
0498
03F4
0419
04E2
0572
054F
04D6
049E
04B7
04C2
0494
0466
0461
0455
041E
0408
046D
0513
054D
04DD
0453
045D
04D3
04FA
049A
044D
048B
04D9
0482
03CD
03D2
04D9
057E
03FA
003F
FC4B
FA42
FA70
FB6A
FBD4
FB90
FB4C
FB63
FB97
FBA7
FBAB
FBCD
FBE7
FBB0
FB30
FAC8
FABB
FAE7
FB08
FB27
FB78
FBED
FC2D
FC13
FBF8
FC3B
FCA4
FC96
FBEC
FB5E
FBA9
FC82
FCC6
FBE6
FAEF
FBB1
FECC
02D6
059E
062C
0568
04D8
0504
054B
0509
047F
0459
04B6
0504
04E1
049E
04B5
050B
051E
04DA
04C9
0544
05C6
0590
04BC
042D
0457
04A6
046F
03FC
0415
04B3
04E6
0433
037B
03E0
04FA
04E3
024F
FE36
FAEE
F9E8
FA91
FB63
FB84
FB3A
FB2A
FB83
FBEC
FC05
FBD2
FBA4
FBB0
FBD7
FBD4
FB98
FB63
FB72
FBA9
FBBF
FBAD
FBC0
FC23
FC92
FCA5
FC53
FBE7
FBA3
FB94
FBBB
FC13
FC55
FC14
FB66
FB56
FD21
00C1
047D
065B
0602
04E2
0485
0500
054D
04D1
0419
03FF
048A
0501
04ED
04A3
04AA
04FA
0527
050D
04F6
0508
04F9
0493
042C
043F
04BB
0510
04FA
04D8
0502
0520
04AE
03FB
0403
04FB
0589
0404
0065
FC8B
FA72
FA63
FB0C
FB14
FA60
F9D0
FA16
FAF4
FBA3
FBAB
FB4D
FB1B
FB4E
FB9B
FBB1
FBB2
FBF2
FC5A
FC6D
FBFE
FB82
FB75
FBC0
FBF7
FBF6
FBE7
FBCB
FB79
FB1C
FB39
FBE5
FC43
FB8B
FA81
FB1F
FE54
02B1
05C6
069C
0640
061D
0676
06A6
0648
05AA
053C
0510
04FC
04F6
0506
0521
0537
0555
0580
059C
0592
0572
0545
04EB
045D
03E1
03C4
0404
0468
04CE
052A
054D
0505
0499
04AE
0550
054F
033F
FF5A
FBBA
FA53
FAF4
FBC9
FB94
FACE
FA93
FB14
FB86
FB4F
FABC
FA73
FA9B
FAD5
FAE5
FAF4
FB2F
FB74
FB8F
FBA0
FBF1
FC79
FCC1
FC69
FBBA
FB5C
FB84
FBA7
FB49
FAC9
FAE1
FB75
FB98
FAFF
FAE1
FCBA
0061
03FD
05DB
05EC
052A
042F
02E5
0172
0087
007E
00CA
00C0
0073
0058
0072
005D
0002
FFBB
FFC6
0004
0044
0088
00C4
00B9
0058
0024
00D1
026B
043D
0580
05D3
052E
0420
03FD
059A
0753
0589
FE66
F4D0
EE3C
ED4B
EF6B
F067
EF33
EE0A
EE79
EF47
EECF
EDAE
EDA3
EEC2
EF6B
EED6
EE21
EE75
EF4E
EF76
EEF3
EEED
EFC1
F053
EFB7
EE9B
EE4E
EEE0
EF32
EEA3
EDDA
EDB4
EE22
EE75
EE63
EE44
EE71
EEC3
EEDE
EEC6
EED6
EF3A
EFA7
EFC1
EF92
EF75
EF99
EFCA
EFB9
EF73
EF5F
EFB7
F027
F031
EFD9
EFA2
EFD4
F020
F037
F050
F0C8
F172
F1AD
F137
F09C
F0A0
F163
F23C
F273
F1FE
F173
F167
F1D9
F23E
F208
F14A
F0BA
F0EE
F19B
F201
F1F1
F1E3
F20E
F210
F1C2
F1AF
F232
F2A2
F232
F15D
F175
F280
F2AB
F10B
F00D
F35C
FB0D
0292
0588
045C
02E0
034D
0463
045A
03AA
03DE
04E9
053C
044C
0369
03A6
0443
0410
0351
0327
03AD
03F0
039A
0374
0411
04E5
0521
04D8
04A5
0495
042E
03A0
03F9
05BC
07E5
08FF
08C8
0834
0818
0872
08D1
08E2
0893
0820
0804
0883
0932
094C
08B4
0849
08DA
09F2
0A45
0965
085F
0847
08CD
08D6
081E
0774
0774
07BD
07B9
079A
0805
08E6
0921
07C7
0556
0360
02EA
036F
03BA
0352
02D2
02E1
0355
038C
035A
0333
0360
0381
0333
02DC
0315
0389
034E
0269
0211
02DD
03B6
0366
029D
02FC
040F
02B8
FCD3
F4A4
EF15
EE6A
F036
F0FB
F053
F03A
F17A
F29C
F25B
F17A
F17E
F27D
F32F
F2D5
F219
F1E8
F249
F2AA
F2C3
F2A1
F255
F214
F242
F2DA
F331
F2DD
F266
F289
F316
F337
F2BA
F263
F2C2
F35E
F375
F32C
F335
F382
F339
F235
F187
F1F1
F2B4
F2BD
F244
F257
F30F
F35A
F2A0
F1BD
F1C6
F288
F2DF
F261
F1CD
F1C4
F1EC
F1BC
F17D
F1BB
F23D
F254
F1F2
F1BF
F20B
F263
F24E
F205
F21C
F2A2
F311
F30C
F2ED
F34B
F41A
F4A7
F476
F3DC
F393
F3E3
F455
F451
F3EC
F3D6
F451
F4AE
F450
F3DF
F468
F574
F539
F38C
F371
F84A
016A
09DF
0D4D
0C43
0AC4
0B48
0C9D
0CB8
0BCC
0B74
0C02
0C26
0AFA
0912
077A
068A
0614
0600
0634
0651
0604
059B
05A5
061A
0658
062E
062C
069D
06EC
0699
0623
0646
06CB
06DF
065D
05F9
0621
0666
063C
05D5
05C2
0604
0611
05C3
0587
0594
05AB
05EC
0716
0958
0B73
0BFC
0B22
0A6D
0AC5
0B7D
0B7C
0ABE
0A1F
0A12
0A2A
09F9
09CD
0A2B
0AEC
0B62
0B34
0AAF
0A53
0A54
0A90
0AB3
0A92
0A67
0A7D
0AB2
0A98
0A2E
0A0C
0A80
0AEB
0A6D
08F8
0761
0655
05BE
055D
0550
0581
052C
03F8
033D
048C
069E
057D
FF01
F632
F08F
F043
F274
F35B
F27E
F1E4
F266
F2C2
F220
F18B
F210
F2DB
F298
F1B1
F1AC
F2BD
F373
F2F2
F237
F299
F3E0
F4B4
F484
F412
F416
F43F
F3FC
F38F
F395
F400
F444
F43D
F44F
F4B2
F535
F5A7
F604
F638
F616
F5AD
F550
F53B
F552
F55A
F55D
F583
F5AD
F58D
F537
F52A
F589
F5BF
F54A
F485
F437
F494
F50A
F503
F478
F3CD
F369
F366
F391
F3A4
F390
F383
F3A1
F3D3
F3E9
F3F7
F452
F502
F578
F539
F4A4
F48B
F502
F54D
F512
F4D5
F4ED
F4DC
F446
F3D8
F458
F53C
F53E
F464
F442
F58A
F698
F5E3
F550
F8E5
017F
0A9D
0EEC
0DFE
0BE2
0BCB
0D0C
0D7A
0CE1
0CC5
0DA7
0E4C
0DD2
0D10
0D27
0DC6
0DD3
0D2C
0CAD
0CBE
0CE3
0CB2
0C65
0C4E
0C60
0C74
0C9D
0CD8
0CB5
0BB1
09FF
0888
07F4
0803
0807
07C5
0783
0785
07CF
0833
0862
081A
0786
0729
0731
072E
06B5
0615
05F8
0676
06EC
06E1
06AF
06E8
076A
0780
0702
06AC
0713
07BE
07C7
071C
06A0
072F
08C9
0AAA
0BE0
0C03
0B87
0B4C
0BAF
0C2C
0C0D
0B59
0ACB
0AE4
0B4E
0B75
0B5C
0B72
0BBD
0BD0
0B9E
0B95
0BBE
0B9D
0B33
0B4C
0C23
0C9D
0BD5
0AD9
0B73
0CEF
0BA4
04F5
FB39
F401
F252
F3ED
F4CD
F3D7
F2E2
F341
F427
F465
F429
F444
F4AC
F4A3
F40B
F39E
F3D0
F42B
F42C
F410
F453
F4C9
F4EF
F4C3
F4B8
F4EF
F513
F4E9
F495
F44C
F418
F3FA
F403
F430
F45A
F470
F4A9
F537
F5DE
F624
F5F5
F5C3
F5E2
F620
F63A
F654
F6A9
F70F
F730
F71C
F727
F753
F740
F6BD
F623
F5F0
F62E
F67B
F69B
F6B2
F6E9
F711
F6E6
F681
F641
F669
F6DD
F743
F746
F6DD
F668
F642
F643
F5F7
F562
F513
F548
F584
F547
F4F6
F554
F63D
F696
F5DF
F529
F5AA
F6E0
F73A
F686
F64B
F72D
F791
F62B
F4FE
F7D3
FF59
076F
0B3D
0A4B
0844
082C
0960
09B2
08DF
088B
09B4
0B94
0D07
0DD7
0E59
0E9C
0E88
0E59
0E73
0EC9
0EDD
0E78
0DF6
0DC8
0DE5
0E01
0DFD
0DD5
0D78
0D02
0CE3
0D63
0E20
0E6F
0E20
0D9D
0D57
0D55
0D5A
0D48
0D2A
0D19
0D1E
0D33
0D1D
0C68
0ADC
0904
07E4
07E8
086A
0879
07F2
0776
0787
07F8
084C
083D
07F3
07C1
07CD
07F1
07F4
07D6
07D5
0814
085A
084F
07EF
07A0
07A9
07C1
0783
071D
0723
079D
07E9
07B6
07A2
086A
09ED
0B6B
0C6B
0CF6
0D14
0CB9
0C3A
0C27
0C6A
0C23
0B1E
0AD0
0C85
0E90
0CE8
05A6
FBFC
F55D
F40D
F594
F666
F5B5
F513
F57F
F638
F654
F61B
F637
F680
F663
F605
F60B
F67F
F6BB
F65A
F5B4
F539
F4E7
F493
F45E
F491
F520
F59C
F5B7
F588
F552
F53A
F552
F5A0
F5E3
F5B8
F539
F518
F5B7
F682
F68F
F5D4
F53B
F574
F621
F669
F60C
F58F
F573
F5A3
F5CE
F5F5
F654
F6D7
F726
F723
F71C
F757
F7AD
F7B9
F75D
F6F1
F6DE
F71E
F74E
F745
F75E
F7F0
F89A
F8A4
F804
F78F
F7E5
F897
F8C3
F854
F810
F855
F871
F7BA
F6CF
F6D4
F7B9
F839
F7D5
F7A5
F892
F9B2
F979
F80E
F71F
F754
F755
F63A
F5ED
F96C
00AB
07BC
0AD2
0A1C
08B8
08B5
0982
09E0
09DA
0A31
0AD5
0B00
0A83
0A1F
0A68
0AF6
0B10
0AA8
0A35
09F1
09CA
09D2
0A24
0A6D
0A29
097D
0962
0AA1
0CD0
0E9C
0F17
0E8B
0DF1
0DDB
0E13
0E31
0E2E
0E45
0E84
0EAA
0E6F
0DDA
0D3E
0CF6
0D20
0D90
0DFB
0E21
0DED
0D8B
0D55
0D7B
0DC4
0DCC
0D7E
0D1C
0CD5
0CA3
0C95
0CE1
0D5A
0D42
0C13
0A66
098C
09EF
0A6E
09D3
0890
082C
0910
09DF
0962
083C
07E1
0887
0906
08B1
0832
0849
089A
0866
07F3
0833
0920
0990
0905
0887
0907
09D3
09BB
091F
0962
0A42
091C
03EE
FC66
F6BD
F562
F6C3
F7A4
F6CC
F587
F53D
F5C1
F622
F618
F61A
F66D
F6BA
F6A0
F63E
F60D
F64E
F6D3
F73B
F74E
F720
F6FC
F71A
F75B
F750
F6BC
F5F5
F5A0
F5F0
F65F
F645
F590
F4E5
F4E4
F587
F62E
F650
F605
F5D5
F61E
F6C4
F755
F76B
F6F3
F64D
F61B
F6B3
F7AC
F824
F7A9
F6CC
F67D
F6E7
F73E
F6EC
F682
F6EF
F7E7
F7E5
F652
F51F
F76D
FE42
070A
0DB0
101F
0F9F
0EE5
0F42
0FE9
0F90
0E44
0D4F
0DA1
0EBE
0F69
0F20
0E95
0E9B
0EFE
0EDB
0DFD
0D43
0D6D
0E1A
0E57
0DF0
0D9D
0DD7
0E26
0DE9
0D60
0D65
0E19
0E72
0D71
0B63
099B
08FB
0939
0978
093C
08B7
085C
085E
0892
08C3
08F1
092D
0955
0928
08B3
0869
08A6
091D
0922
08A6
0876
0922
09F1
09BF
08CD
08C0
0A1C
0A9B
0737
FFEE
F889
F507
F5B5
F78A
F7E5
F709
F6B5
F76F
F820
F7EC
F751
F737
F79D
F7C7
F760
F6DA
F6C1
F709
F74B
F75F
F77A
F7C7
F829
F872
F88A
F85D
F7D4
F713
F694
F6C2
F773
F7FB
F7D9
F732
F68D
F62F
F5ED
F59F
F577
F5AE
F615
F643
F62F
F63E
F6AA
F721
F73F
F719
F707
F714
F6F5
F6A0
F67C
F6C4
F710
F6E2
F681
F6A0
F72E
F731
F66F
F6A1
FA24
0131
08F9
0E03
0F42
0E8F
0E43
0EED
0F82
0F40
0EA9
0E98
0F04
0F20
0E8C
0DE7
0DF6
0E8B
0EB1
0DF3
0D16
0D27
0E11
0EAF
0E55
0DBC
0DEF
0ED2
0F43
0EB9
0E12
0E65
0F63
0F82
0DD9
0B47
096F
08F0
08FE
089E
07D2
0768
07E0
08C7
0937
08DE
0856
0850
08B4
08DE
08A5
08AA
0954
0A0A
09EC
0938
091C
09E8
0A3C
08FF
0781
0821
0A77
0A76
04DA
FBAC
F4D6
F3E8
F6A7
F85B
F75B
F5F7
F668
F7E3
F85B
F7AF
F786
F891
F985
F923
F801
F79A
F837
F8C4
F87D
F7E6
F7CB
F80C
F7F9
F784
F745
F770
F77B
F708
F6A9
F71E
F82B
F8AE
F805
F6D5
F639
F680
F70D
F75C
F792
F7EB
F822
F7DB
F75E
F748
F791
F783
F6CE
F61A
F625
F6B0
F6EE
F6B8
F6AF
F717
F74F
F6F5
F6D0
F7B2
F8CC
F885
F745
F818
FD5E
0594
0C8A
0FB2
1022
103D
10AD
108F
0FB7
0F3A
0F9B
0FE3
0F3B
0E6C
0EBA
0FE7
1079
0FCF
0EE1
0EBD
0F26
0F35
0EBE
0E5E
0E6A
0E96
0EB5
0F06
0F76
0F5A
0E81
0DD6
0E31
0EDD
0E47
0C17
09CA
08DB
0908
0907
086F
0811
086A
08C1
0853
07B3
080F
0956
0A1E
098C
0885
085E
08FD
0924
086C
07F0
0897
0974
08F9
077E
073D
0928
0AA2
07DF
007D
F89F
F4CF
F582
F772
F7D3
F6F7
F6A0
F72A
F765
F6CE
F66B
F728
F866
F8E5
F885
F83B
F887
F8CE
F86F
F7B5
F75B
F783
F7A4
F775
F75F
F7DE
F8B8
F933
F8EA
F833
F7C0
F801
F8CA
F965
F932
F847
F761
F70B
F71B
F71D
F6F7
F6E0
F6DD
F6AC
F63D
F5E5
F5F2
F634
F63F
F611
F61B
F690
F718
F752
F75F
F79F
F829
F8AC
F89E
F7A0
F62F
F616
F95C
0012
077E
0C49
0DAB
0DC6
0EB2
1004
1007
0EBD
0E17
0F1B
106A
1064
0F90
0F8B
1062
1088
0F5A
0E3D
0E88
0F8D
0FB8
0F17
0F26
1040
10C9
0FA2
0E0A
0DDF
0EEF
0F7F
0F0C
0EE5
0FB7
100A
0E3D
0B24
0952
09C8
0ABB
0A24
0866
077A
082A
0955
09D1
09C0
09CB
09FA
09F5
09D3
09ED
0A01
096A
085B
07FD
08E7
09FD
09D9
08ED
0918
0AA2
0ACB
068A
FE8E
F753
F4BF
F663
F8A6
F8FF
F80C
F79B
F805
F847
F7F6
F7CB
F841
F8BF
F89D
F831
F819
F828
F7CC
F73F
F760
F848
F8E5
F877
F7CB
F81B
F92A
F96C
F842
F6EC
F6C3
F77A
F7E3
F7D0
F80A
F8BA
F8F3
F829
F72F
F707
F75C
F701
F5DC
F534
F5DB
F6E6
F703
F64F
F5FD
F67D
F705
F6F7
F6C6
F70C
F76A
F72F
F6B3
F71F
F88A
F942
F7E5
F5EF
F6EF
FCAE
04B8
0A98
0C5B
0C22
0D1F
0FC3
11AA
1113
0F38
0E92
0FA9
10B8
1061
0F6A
0F44
0FF2
104E
0FFB
0FCA
1037
1080
0FDE
0EF1
0EF2
0FCA
1021
0F67
0EB4
0F07
0FBC
0FA2
0EE4
0EA7
0F06
0EB4
0CEA
0AC0
09CD
0A0D
0A1F
096A
08E6
0972
0A70
0ABC
0A4E
09F4
09E7
09A8
0919
08D5
0922
0961
08FE
086D
087B
08EB
08BC
07E5
07CC
0930
0A3F
07F7
0198
F9EE
F4CF
F3B5
F50F
F67C
F70D
F742
F79C
F7D3
F779
F6CF
F677
F6A8
F6FC
F71B
F725
F75B
F79F
F790
F726
F6D0
F6EC
F749
F77F
F78C
F7C3
F824
F847
F7F9
F791
F76D
F78C
F7D9
F883
F980
FA16
F975
F7E6
F6C0
F6D5
F760
F717
F605
F577
F618
F70A
F751
F73F
F7A8
F852
F835
F73A
F69D
F72D
F80F
F809
F774
F7BA
F8F8
F971
F83C
F77E
FA77
0165
089C
0C3F
0C3C
0BBC
0D22
0F94
10BA
1001
0F24
0FAA
10F4
114B
103C
0EFE
0EAD
0EF9
0EED
0E6B
0E22
0E57
0E7B
0E33
0E1A
0ED9
0FE2
0FFB
0F11
0E84
0F41
105A
103F
0EE0
0DB4
0DAF
0E0E
0D78
0BC7
0A19
0952
094D
0977
0984
095E
08EF
0871
0870
0905
0980
0955
08F5
0924
09B4
09B2
08EC
086E
0901
09D3
098C
087D
0876
09F7
0A8E
0733
FFFD
F897
F4D0
F55B
F7EB
F9D0
F9FB
F8FD
F7DF
F74A
F757
F7AE
F7D0
F794
F75B
F7A7
F86D
F914
F918
F899
F824
F81F
F86C
F899
F86A
F816
F7F6
F80E
F814
F7ED
F7C9
F7CD
F7E9
F811
F865
F8DC
F902
F86E
F767
F6CB
F709
F797
F7B3
F770
F76F
F7B9
F7A4
F706
F6B3
F750
F83A
F86F
F801
F7E9
F85E
F866
F768
F654
F658
F6EB
F677
F52F
F5E5
FAF2
02E4
097D
0BFC
0B88
0B37
0C90
0E87
0F74
0F32
0EED
0F75
104E
1077
0FB0
0EAD
0E36
0E46
0E37
0DB2
0D37
0D6F
0E1E
0E5E
0DDF
0D6B
0DC3
0E8C
0ECA
0E3F
0DA8
0DAE
0E1F
0E54
0E12
0D93
0CF0
0C0B
0B10
0A74
0A44
09F3
0931
0889
08B3
0990
0A58
0A97
0A8B
0A8E
0A94
0A61
09EC
0961
08F1
08D1
093B
0A04
0A70
09FC
094D
097A
0A0E
08A5
0379
FC00
F613
F437
F56D
F6F3
F76D
F798
F840
F8D3
F86E
F782
F768
F86F
F942
F8A3
F70C
F611
F66E
F744
F763
F6DE
F6DA
F80A
F9C7
FAC1
FA5C
F91F
F808
F7AD
F7F4
F855
F85A
F817
F827
F8E9
F9BC
F975
F7D1
F60C
F5A4
F6A2
F797
F775
F6BC
F686
F6EA
F724
F711
F76C
F858
F8CF
F816
F703
F6D5
F760
F770
F6E4
F702
F844
F902
F7C2
F647
F86B
FF5F
07A0
0CAA
0DB9
0D99
0E81
0FD4
0FFE
0F01
0E38
0E60
0EFD
0F77
0FE0
104A
1040
0F83
0EAA
0E6F
0ECE
0F54
0FCB
1011
0FCF
0F01
0E68
0EB0
0F55
0F35
0E4D
0DFF
0F02
0FDC
0E94
0BA0
09B3
0A3D
0B97
0B7C
0A20
096A
09E4
0A36
09AB
0982
0AA8
0B4B
0850
0154
F9D3
F5A6
F53C
F60C
F606
F55B
F541
F61F
F750
F7FB
F7B6
F6B1
F5A9
F57D
F65D
F773
F7AF
F706
F685
F706
F830
F90B
F926
F8CB
F866
F82B
F836
F877
F87C
F7CE
F6D3
F6B6
F7F7
F95B
F91F
F73C
F5AD
F603
F776
F822
F7AE
F787
F854
F8A3
F730
F5CF
F836
FF74
07E2
0C97
0C61
0A42
0981
0A71
0B52
0B20
0A69
09F3
09C9
09D1
0A3D
0AE7
0B12
0A73
09D1
09FB
0A90
0A97
0A05
09B5
09F3
0A03
0986
0986
0B2E
0DD2
0F74
0F4E
0EB0
0EEC
0F97
0F9D
0F0B
0EB2
0EA7
0E59
0DE4
0E05
0EA1
0E9D
0DCC
0DDB
0FB9
10BD
0CAC
033A
F9AE
F59C
F721
F9C7
FA26
F8D3
F7F1
F7F7
F7DD
F736
F6A9
F694
F694
F689
F6ED
F7A5
F7B1
F6BA
F5EB
F64C
F719
F6EF
F5F9
F5A9
F662
F6DB
F62E
F556
F5B3
F6D0
F6FB
F5F0
F558
F63E
F779
F793
F6F9
F70B
F7D5
F840
F82B
F890
F95F
F8F5
F6F5
F683
FB86
0578
0EBD
1238
1078
0E2D
0E6F
1031
1103
106F
0FCE
0FE7
1017
0F9B
0EAC
0DF9
0DCC
0E23
0F00
1009
1045
0EFA
0CAA
0AAE
09BD
0975
093F
092A
097C
09EE
09F4
099E
0991
0A0A
0A80
0A7B
0A37
0A11
09E1
0979
094E
09D7
0A71
09F5
08AC
0885
0A36
0AEB
06B5
FDB5
F53A
F287
F548
F88D
F8B3
F6BE
F5AF
F64D
F6FD
F6CA
F6B1
F7A0
F8BE
F8BC
F7CB
F726
F73A
F769
F762
F79C
F853
F8EE
F8D4
F847
F7F4
F7FE
F816
F850
F90A
F9E5
F9D3
F884
F6FD
F644
F633
F638
F663
F6ED
F75F
F736
F70E
F7DB
F8F2
F84C
F5C6
F4F6
F9B8
02F3
0AC7
0CD5
0AB9
092D
0A1E
0B8F
0B82
0AA8
0A90
0B02
0A94
0935
0891
09C7
0C00
0DCB
0ED3
0F7A
0FA4
0F0A
0E1E
0DAC
0DD4
0E20
0E69
0EE0
0F42
0EF6
0E1D
0DC9
0E99
0FA4
0F9B
0EAB
0E3D
0EC4
0F20
0EA6
0E56
0F1E
0FEF
0F20
0D2C
0C37
0C8A
0B26
0541
FC73
F5CA
F475
F6AD
F86D
F800
F6BC
F62C
F62A
F5EC
F57F
F580
F601
F66F
F671
F641
F61E
F5EF
F5AB
F5AF
F647
F729
F7B8
F7B1
F745
F6D0
F6B3
F746
F867
F948
F912
F7F7
F71F
F74C
F7E9
F7F8
F792
F7B2
F883
F8E9
F843
F7B0
F87F
F9D9
F983
F787
F7A0
FD77
07AC
1034
1262
0F90
0CEC
0D8B
0FDD
10B7
0F37
0D03
0BAA
0B1A
0A9F
0A28
0A16
0A51
0A58
09F6
0965
08ED
08B8
08D3
090F
0911
08D5
08E0
099A
0A8E
0AC9
0A0A
091E
08D9
0912
0926
0918
095E
09CB
09CC
09DA
0B43
0DE1
0F54
0DF4
0B9D
0BB2
0E19
0E2A
0800
FDDC
F656
F531
F7CD
F945
F82E
F6C9
F6D7
F77A
F748
F68A
F691
F7AC
F8C7
F8E7
F838
F791
F786
F821
F8EA
F909
F806
F69C
F62B
F6ED
F783
F6E8
F5EC
F5F7
F6E7
F752
F6C0
F656
F6E8
F77B
F6C5
F574
F573
F701
F82A
F7B4
F6F3
F77B
F856
F78D
F5F1
F726
FD1B
04F6
09F9
0AD3
0A88
0C05
0EA3
0FE7
0F43
0E84
0EFB
0FE5
0FEB
0F11
0E68
0E87
0EFE
0F36
0F28
0F12
0EF5
0EB0
0E41
0DC1
0D50
0D3A
0DCB
0EB2
0F0D
0E78
0DAE
0D8C
0DA9
0CC0
0A92
08A3
0863
0938
0956
084B
0786
0808
08D6
08AB
082F
08F5
0A4D
08E8
02B9
FA42
F493
F401
F61F
F731
F640
F4FB
F4B1
F501
F535
F570
F5F9
F669
F650
F62F
F6E5
F837
F8E6
F86F
F7C2
F7DB
F863
F878
F80F
F7CB
F7D0
F7B1
F770
F7A3
F870
F916
F8FF
F8AE
F8EA
F95B
F90A
F825
F7FC
F8E0
F966
F89D
F7B4
F817
F8D8
F7DA
F5B8
F66A
FCB9
0605
0C6C
0D13
0AB4
098C
0A89
0B9F
0B74
0AC0
0A78
0A60
09F6
097E
097C
09B7
0994
0925
0908
0953
096E
0936
0945
09CB
0A12
09CB
09FD
0B99
0DCC
0ED3
0E46
0D85
0DB1
0E4F
0E64
0E1C
0E45
0EAA
0E4B
0D42
0CF4
0DC7
0E3A
0D4D
0C86
0DB8
0F44
0CD5
04A8
FAAD
F4D8
F4E2
F72C
F7A9
F628
F503
F556
F621
F671
F68B
F6C4
F69F
F5B8
F4C4
F4C9
F5B2
F673
F689
F680
F6D9
F744
F758
F75D
F7B8
F81C
F808
F7BF
F7EA
F876
F8A1
F83C
F814
F8A2
F90A
F843
F6DF
F683
F796
F8B2
F8CD
F89D
F8F2
F8E6
F76B
F647
F95C
01E7
0BC2
1116
107A
0DE5
0D74
0F0A
0FF0
0F20
0E0B
0DDA
0DE3
0D57
0CE3
0D94
0EF4
0F7B
0EB8
0DCB
0D80
0D13
0B9C
09BA
08D5
0926
0991
093E
087A
07F4
07D5
07E8
081C
086D
089D
087D
085C
089C
08F9
08EE
08C9
0952
0A34
0A0C
08AD
0812
099C
0B18
086E
00CD
F8A1
F523
F6B8
F926
F908
F72B
F616
F648
F671
F634
F68D
F7B6
F856
F779
F627
F608
F71D
F7E1
F781
F6C5
F694
F6B1
F697
F698
F731
F7E7
F7D9
F730
F6FC
F7AB
F86D
F864
F7B3
F70D
F6B3
F675
F663
F6A7
F6D1
F649
F58B
F5CB
F6ED
F719
F594
F4F9
F8E7
014B
098A
0D1A
0C15
0A45
0A4B
0B58
0B96
0B0D
0AEE
0B3D
0AE3
09C9
0968
0AC9
0D02
0E47
0E03
0D30
0CDA
0D1D
0D98
0E3C
0F10
0FC3
0FE8
0F81
0ED6
0E0C
0D47
0CDF
0D05
0D4F
0D24
0CA2
0C8F
0D3E
0E01
0E16
0DB4
0D93
0D90
0CDB
0B8A
0AE5
0B43
0A7F
0602
FE4B
F742
F45F
F52B
F65C
F5DF
F4AD
F4A3
F5D2
F6D3
F6EC
F6B6
F6D0
F6EB
F680
F5C3
F55A
F570
F59B
F5A2
F5D4
F669
F702
F714
F6A1
F63A
F667
F746
F86F
F91C
F8B0
F76F
F676
F6A1
F78B
F810
F7CC
F781
F7D1
F82F
F7C4
F705
F731
F82D
F83D
F6CE
F688
FAED
03D4
0C8C
1066
0F5F
0D7D
0DD8
0F96
0FF5
0DFD
0B2C
092D
083B
07DB
0802
08EB
0A3C
0B11
0AF5
0A67
0A26
0A42
0A1E
0950
0841
07D3
086E
0975
09C0
08CC
076A
06F1
07B4
08AA
08BE
0800
0742
06FA
071A
07DD
09CE
0CA2
0EBB
0EC1
0D78
0CF2
0D86
0CA6
07B9
FFAA
F88F
F59A
F61F
F714
F6B0
F5D0
F5F3
F6FD
F793
F717
F663
F667
F6E2
F6E3
F65C
F6A0
F914
FD7D
01E8
046E
04EE
04CA
0524
05B9
05A2
04C7
040D
0422
0497
0498
041F
03F6
0479
0506
04E1
0440
03E6
03F6
03D6
033E
02D9
035A
044F
048C
03D9
03AA
05A0
0989
0D53
0F1C
0EEE
0E3D
0E16
0E38
0DEF
0D45
0CF7
0D56
0DC1
0D7A
0CB9
0C75
0D27
0E19
0E3F
0D7A
0CA5
0C73
0CA2
0C9D
0C79
0CD3
0D96
0D83
0B66
07A7
0438
02B2
02DD
033C
02E1
0244
0259
033F
042A
046B
042A
03EA
03CA
0384
0313
02DC
0315
0348
02CC
01C3
0127
01B1
02E3
038C
034E
0341
04CC
07F1
0B19
0CA1
0C75
0BDB
0BD8
0C2A
0BE5
0ACB
09AD
0975
0A2C
0B15
0B8A
0B87
0B64
0B5F
0B88
0BE4
0C5E
0CA5
0C68
0BDA
0BAB
0C4B
0D18
0CB2
0A48
0698
036B
01FC
01FE
0235
01DF
0154
0156
01FA
0291
0296
0255
0274
02FD
0347
02E1
022A
01CA
01C0
0172
00B6
0041
00B8
019E
01D3
014B
0194
042D
0882
0C2A
0D4B
0C4D
0B10
0ACD
0B2E
0B59
0B2C
0B27
0B77
0BAC
0B6A
0AF3
0AC6
0AF0
0B0B
0AE2
0AD1
0B49
0C1E
0C9A
0C52
0BB7
0B87
0BAA
0AFC
087F
04B8
0189
0075
012F
021E
022B
01B0
0196
020C
0277
0275
0263
02B3
0333
0352
02F1
0284
0252
020A
0159
0090
004E
0096
00BC
0064
0054
01C4
04E9
0871
0A9C
0ADE
0A2E
09DD
0A4A
0AD3
0AD1
0A57
09F2
09D7
09B0
093A
08D0
0902
09B3
0A13
099C
08D6
08B7
095B
09D3
096F
08BA
08BA
094F
08FE
06B1
0347
00DF
0093
016A
019D
009B
FF69
FF35
0006
00EC
012C
00E3
00A0
00B3
00FB
012C
011D
00D9
0087
0056
006E
00D8
015B
018F
014B
010B
01BC
03DC
06C7
0919
09F3
09C4
09A4
0A07
0A67
0A3D
09DA
09E5
0A5D
0A90
0A2B
09B9
09D6
0A31
09EA
08E0
080F
0841
08EA
08CF
07C1
0703
07A9
08F9
08E8
064F
0253
FF56
FEB1
FFA6
006F
0019
FF31
FED1
FF5D
0030
0076
0014
FF97
FF6A
FF75
FF77
FF7F
FFBD
000D
0007
FF96
FF2F
FF29
FF2C
FEB3
FE2A
FEEE
01BD
057A
0802
085F
07B3
07BA
08C7
0999
0930
081D
07BF
088E
09AC
0A1C
09DD
099E
09A4
098A
0914
08B5
08F8
0994
0995
089E
078D
076B
07DF
0746
0491
00C4
FE15
FDA0
FE66
FEBC
FE44
FDFA
FE7A
FF09
FEA6
FD8E
FCFC
FD8E
FE8D
FF09
FF16
FF74
002E
006A
FFB9
FEF4
FF29
FFFF
0003
FEAF
FD98
FEF0
02FD
0784
09F7
09DC
08D5
0889
08FD
0915
083B
071B
06B5
0727
079E
0774
06F2
06D7
0753
07CF
07CA
0785
079B
081C
0882
088C
08B9
0976
09FD
08C2
0549
012A
FEBC
FEBE
FFB9
FFD5
FEDD
FE11
FE4D
FEFC
FF05
FE43
FD82
FD51
FD65
FD58
FD6B
FE10
FEF1
FF09
FDFE
FCD2
FCC7
FDBF
FE4E
FDAE
FD0E
FE5F
01E8
05B7
07AD
07B8
077E
081B
08E2
089F
0775
06CB
0774
0899
08DD
0810
0731
06F5
06F0
067B
05E1
0611
073B
084B
082C
072B
0699
071C
07B8
06D2
0405
00A3
FE76
FE19
FEB2
FF16
FEE9
FE90
FE5A
FE0A
FD58
FC92
FC67
FD0E
FDEB
FE4B
FE36
FE49
FEAF
FED2
FE3B
FD62
FD29
FD8D
FD87
FC8C
FBC7
FD25
010D
0588
0812
07FD
06B9
05F7
0606
0632
0617
060C
065C
06B7
06BB
06A9
0718
07F9
0872
07E5
06D2
064B
0695
06D1
0633
0540
0546
0683
075D
05F4
0255
FEAE
FD12
FD6A
FDE5
FD49
FC32
FBF2
FCB6
FD66
FD29
FC73
FC3E
FCB5
FD2E
FD3E
FD3C
FD89
FDC7
FD5B
FC73
FC11
FCC8
FDD6
FDFE
FD27
FCBC
FE3C
018B
04F0
06AA
067D
05A4
056F
0614
06D2
06FF
06B8
0693
06D9
073D
0757
071E
06CE
0683
062F
05F7
062B
06BB
070C
06AD
061B
0646
0728
0743
0517
010E
FD72
FC2E
FCF3
FDDB
FDA7
FCCF
FC6E
FCB4
FCE6
FC93
FC2B
FC36
FC80
FC6F
FBFC
FBD7
FC76
FD5D
FDB4
FD4E
FCDD
FCF2
FD33
FCDF
FC09
FBE7
FDAC
0116
0473
062B
0622
058E
0589
060C
065B
0614
0598
0569
0591
05C4
05E6
0615
0646
062D
05B7
055C
05A0
0654
06A0
0614
055C
058E
06B6
0763
0600
028B
FEC0
FC7C
FC14
FC59
FC1B
FB59
FAF4
FB69
FC3C
FC9F
FC64
FC0D
FC13
FC51
FC62
FC38
FC2C
FC6C
FCB1
FCAC
FC79
FC6C
FC79
FC40
FBD3
FC18
FE00
014B
0470
0600
05FF
059F
05C8
063C
063C
05A8
0513
04EB
04F5
04D7
04BB
050F
05B0
05E0
0534
0450
0443
0539
0639
065E
05F2
05F5
0689
065E
041E
0032
FCBB
FB8B
FC5B
FD4C
FD03
FBF8
FB98
FC71
FD92
FDBB
FCCC
FBC5
FB89
FBFD
FC69
FC69
FC3B
FC2E
FC2E
FBFF
FBB8
FBAE
FBE4
FBFA
FBD0
FC0F
FDA3
0096
03B2
058D
05D3
055C
050C
04EE
0494
040A
03E7
0477
0531
0554
04E0
0484
04AD
04F6
04D7
0481
04A5
055F
05DD
056F
04A0
04AD
05C5
0651
0481
0076
FC7D
FAD0
FB77
FC8E
FC8F
FBCA
FB92
FC53
FD20
FCFA
FC14
FB63
FB57
FB64
FB02
FA80
FA8D
FB29
FB8C
FB35
FAA4
FAA3
FB1E
FB49
FAEF
FB2C
FD49
00FE
0461
05BD
0540
0485
04AD
055B
0589
04F6
0453
043F
0494
04D4
04F8
0550
05D0
05E4
053A
0465
0451
0514
05AE
053C
0424
03A3
042C
0491
032F
FFE6
FC78
FAD4
FB37
FC2F
FC64
FBE7
FBAF
FC18
FC73
FC01
FB00
FA5A
FA84
FB0A
FB45
FB2B
FB1E
FB2E
FB09
FAA7
FA9F
FB57
FC2B
FBFE
FAD0
FA53
FC47
0060
0441
05CA
0523
041E
03F8
043F
0411
03A1
03EC
0521
0621
05EE
0503
04B3
0553
05CF
052D
03F9
0392
0454
0528
0509
046E
048D
056C
0574
0326
FF07
FB4D
F9C9
FA57
FB6F
FBD6
FB86
FB26
FB18
FB35
FB35
FB04
FAB4
FA52
F9FB
F9E6
FA3F
FAD6
FB34
FB19
FAC9
FABE
FAF9
FAEA
FA3B
F993
FA43
FCF4
00B5
03A3
049B
0423
03A6
03EB
0484
04A9
0444
03F2
0425
0498
04C4
049A
048D
04DA
0529
050C
04AF
04AB
052D
058E
0522
0437
03CD
0426
040B
020B
FE66
FB31
FA3D
FB35
FC32
FBF7
FB0F
FAA0
FAC5
FAAA
FA02
F987
F9E2
FAAE
FB16
FB09
FB2B
FBA2
FBAB
FAC2
F9A0
F979
FA56
FAED
FA68
F9B3
FA8F
FD7C
0120
03B9
04B0
049F
044C
040F
0402
043E
04A4
04CD
047F
0409
03EF
043B
0471
043B
03D8
03C8
0422
0484
0488
0441
041D
046E
0505
0537
043B
01C7
FE7F
FBAD
FA4A
FA39
FA80
FA54
F9CD
F98B
F9D6
FA50
FA77
FA47
FA17
FA11
FA04
F9CF
F9B1
F9F4
FA6B
FA91
FA3D
F9E8
FA0B
FA64
FA4F
F9F4
FA9E
FD66
0194
04EC
05D4
04D7
03D7
03E5
0480
04B8
0482
046D
0496
0482
040C
03C2
0407
0467
0441
03C6
03B1
0415
042E
039E
0338
03CF
0491
037D
FFCE
FB56
F8BF
F8D5
FA18
FAC5
FA96
FA45
FA29
F9F6
F99D
F99C
FA30
FAC7
FAB3
FA12
F9A1
F9B8
F9FF
FA16
FA0D
FA08
F9D5
F959
F93E
FA9E
FDBD
016F
040F
0502
04F0
04B9
0491
0445
03E9
03D2
0409
041E
03BA
032A
0308
0386
043E
04BB
04E6
04DD
04A3
0445
041A
0464
0498
0379
005F
FC52
F965
F8B4
F95B
F9AC
F925
F8B5
F929
FA08
FA55
F9F9
F9C3
FA27
FAA4
FA9D
FA3F
FA17
FA1F
F9E3
F975
F985
FA38
FAAA
FA4B
FA2D
FC14
0015
03F5
0573
04B2
03B4
03C4
0444
0421
0385
035A
03BF
03E8
0374
0309
0343
03BE
03B5
0343
0332
03B5
040A
03B1
034E
03A0
03FC
02BF
FF66
FB84
F938
F90E
F9CF
FA3C
FA35
FA32
FA3C
F9FB
F988
F974
F9EC
FA5D
FA30
F9A0
F966
F9C5
FA41
FA67
FA5F
FA7A
FA7C
F9E9
F926
F9A9
FC79
00B0
03F0
04B0
03A2
02B8
02F8
03C5
041A
03E6
03C4
03E0
03C9
0356
0311
0362
03DC
03D1
0349
02E6
02E2
02D8
02AC
02FF
0407
0475
0275
FE24
FA09
F895
F991
FAB1
FA6D
F966
F8EF
F933
F96F
F963
F99B
FA39
FA86
FA10
F97F
F9A3
FA30
FA36
F9A7
F979
FA08
FA50
F975
F888
F9B5
FD81
01CC
0407
03E6
0328
032E
03B0
03D5
039F
03A5
03E9
03CD
0324
0299
02BE
0335
033F
02E5
02E1
0375
03F7
03CD
0365
0397
042E
03AD
00F6
FCDA
F993
F893
F938
F9D5
F9A0
F931
F947
F9B6
F9CA
F962
F91A
F961
F9DF
F9FF
F9C1
F993
F991
F975
F939
F940
F992
F98C
F8E6
F8BB
FAA7
FEB3
02B3
045C
03B0
02AB
02BF
036A
0384
0306
02D4
033A
0394
036B
032A
034B
0382
034C
02F2
0326
03C0
03BF
02E5
0263
032B
041A
02EC
FF1E
FAE1
F8C9
F914
F9E9
F9E6
F973
F97C
F9DD
F9CC
F93E
F8F5
F943
F98A
F93F
F8CD
F8F4
F996
F9D9
F96F
F910
F967
F9FF
F9E4
F944
F9A5
FC27
FFF6
02F4
03DF
035E
02E9
0311
0343
02FD
02A7
02E4
038E
03E0
0393
033C
0369
03CB
03AF
030D
0298
02BE
0312
0315
02FF
0336
0325
0185
FE1A
FA7E
F89F
F8B3
F94F
F952
F90B
F93B
F9B7
F9B2
F918
F8B9
F901
F94F
F8FE
F872
F886
F938
F9B5
F99D
F978
F9AB
F9AE
F902
F886
F9E9
FD83
0182
03BF
03E7
0356
0326
0333
0306
02D5
0314
0389
0388
0307
02D3
0367
0425
041F
0361
02D8
02FB
033D
030A
02C6
032F
03EF
0371
0099
FC57
F901
F80E
F8CD
F983
F95E
F8EA
F8DD
F91A
F91E
F8EB
F8F9
F95A
F97F
F90D
F884
F899
F92A
F96A
F917
F8D7
F923
F977
F936
F90F
FA9C
FE45
0234
0418
03A6
02B1
02D0
03AF
040C
039D
0334
0358
0396
0362
02FD
02F6
033F
0351
0313
0302
034A
036B
0314
02D3
0336
038E
0255
FF1A
FB64
F937
F901
F97C
F96F
F8EC
F8A4
F8B5
F8AD
F876
F887
F90F
F987
F96C
F901
F8F2
F95A
F9A7
F982
F952
F982
F9B4
F947
F8A4
F94F
FC35
0044
033C
03E6
0324
02A2
02F7
0374
0382
036E
03B8
0419
03DD
030C
028C
02F2
03AD
03C7
0322
0284
0271
029F
02B4
02FA
03A6
03C4
01CD
FDB0
F98C
F7C6
F882
F9BD
F9C3
F8F4
F8B0
F940
F999
F911
F859
F86E
F930
F9A3
F957
F8D9
F8D1
F937
F9AE
FA17
FA5B
FA0D
F905
F84C
F998
FD56
01B0
0430
0437
0359
0333
03B2
03B5
02F1
0250
029C
0370
03E4
03BB
0379
0373
0379
035E
034C
0354
0320
028C
0239
02D4
03D1
036A
008E
FC61
F94C
F87D
F8E6
F8E7
F851
F83B
F924
FA1F
FA1D
F958
F8E7
F92F
F978
F92B
F8BA
F8E2
F97D
F9B5
F951
F904
F946
F98D
F946
F931
FAD1
FE63
0217
03E7
03C6
035B
03BB
043E
03DB
02D8
0269
02F4
0391
0363
02C4
02A2
0322
0389
0360
030A
0303
0328
0324
032D
0391
03B6
024C
FEF4
FB2C
F8FE
F8E0
F96B
F941
F899
F88B
F94E
F9E7
F995
F8D9
F8BD
F967
FA0E
FA13
F9AF
F963
F943
F928
F934
F98F
F9CE
F958
F899
F92D
FC2D
0077
037A
03E8
02F9
02B6
0380
0405
036D
028E
02A1
037E
03E5
0358
02AB
02AA
0305
0308
02D4
0306
037E
0362
0298
0245
031B
03C4
0211
FDD6
F9A5
F81A
F90B
FA21
F9D9
F8EF
F8C9
F975
F9DF
F98A
F91C
F930
F97B
F972
F934
F944
F990
F993
F947
F955
F9EF
FA3D
F986
F8B4
F9C3
FD5E
01A6
03FE
03C2
02AE
0289
0339
037D
02EF
0276
02C8
0360
035E
02D6
02AC
032C
03A3
0367
02CA
0276
026D
023F
021B
02AD
03A1
0340
004F
FBF5
F8E5
F870
F946
F971
F8C9
F8A4
F97F
FA2E
F9B1
F8C0
F8B1
F97D
F9DF
F949
F8B6
F922
FA11
FA58
F9E2
F9A5
F9F3
F9E0
F8F8
F896
FA8B
FE9F
0267
03E2
0378
02FA
0346
03A9
0361
02CF
02BE
032D
0373
034E
0324
0325
02EB
0240
01B6
01F7
02B4
02F2
0271
022A
02E6
03B5
02A3
FF16
FAE1
F87F
F882
F957
F963
F8B6
F867
F8E1
F974
F981
F940
F934
F951
F93C
F910
F945
F9D3
FA12
F9BA
F96D
F9C0
FA26
F9A6
F89F
F8F5
FBEE
004F
0361
03D1
02E1
028D
0339
03C8
037A
02D2
029B
02CB
02D9
02B4
02CC
0335
036B
030F
0280
024B
0260
0251
0235
029F
037D
0388
016F
FD88
F9DD
F848
F8B8
F995
F9A1
F913
F8CE
F90C
F94A
F92D
F905
F937
F999
F9B5
F97C
F956
F97C
F9AB
F9A9
F9A7
F9CE
F9B4
F8F8
F85D
F98B
FD1A
0165
03E8
03D4
02B1
0258
02EE
0359
031D
02E4
032F
037B
0323
027F
0261
02D0
0306
02B4
0275
02BF
0310
02C8
0269
02F9
0415
03B7
0089
FBE9
F8B6
F844
F946
F9C9
F95F
F8FA
F92C
F97A
F959
F90A
F912
F95C
F973
F948
F93E
F973
F994
F975
F966
F99B
F9A8
F905
F824
F874
FAF6
FEF3
0270
03F3
03A3
02CB
0275
02B4
0308
031B
030A
030D
031E
0318
0306
0312
0332
032C
02EF
02BA
02C7
02F8
0316
033D
03A0
03C7
0285
FF43
FB31
F884
F83F
F94D
F9F1
F9B2
F955
F965
F989
F95C
F922
F940
F969
F91B
F89F
F8C5
F986
F9DF
F956
F8D1
F930
F9C7
F952
F842
F8CA
FC27
00A7
0355
034F
025F
0255
02FC
032E
02CE
02AD
0307
0345
031F
0310
0364
03A3
035D
0303
0337
03A2
0366
02AC
0292
0335
02DA
000B
FBE1
F90C
F8C6
F9B7
F9FF
F966
F904
F962
F9E1
F9E1
F994
F965
F94A
F920
F91B
F951
F95C
F901
F8C6
F934
F9D0
F9B4
F92F
F9E7
FCE2
00E4
0386
03CA
02E8
0280
02D3
032F
0337
0318
02EE
02BB
02B6
0304
0349
0313
02A2
02B4
0359
03B1
032E
0293
02DA
0351
0212
FE97
FAD9
F910
F932
F98F
F93F
F8E5
F92C
F9AE
F9B9
F967
F94A
F968
F952
F91B
F943
F9B1
F9A2
F904
F8D2
F97F
F9FB
F95C
F8C7
FA63
FE5C
023E
03B2
0318
0293
031E
03BA
0372
02CC
02B5
0303
0309
02D8
02F9
0352
034F
02F7
02EC
0346
0353
02CB
0285
031D
036B
018B
FD81
F9C1
F871
F911
F99C
F939
F8B5
F8D0
F93F
F96E
F95D
F958
F959
F93F
F939
F979
F9A3
F944
F8C5
F8FF
F9BC
F9BA
F8B8
F88F
FB1A
FF90
031D
0406
033F
02B8
030B
0370
0368
034F
0366
034D
02E2
02B5
030E
034E
02EA
026E
029E
0329
032D
02C0
02E2
039C
0339
0049
FBEA
F8E1
F876
F945
F97B
F912
F906
F96A
F96B
F8DF
F890
F8E7
F94D
F934
F8F8
F935
F9AF
F9B7
F962
F961
F9A4
F94E
F882
F915
FC61
010C
041D
0442
02F7
0258
02C5
0329
02EC
029E
02CF
0338
035C
034E
034F
0341
0302
02D9
02F0
02DF
0262
021E
02CE
03BA
02EB
FF74
FAFD
F839
F80E
F8FF
F964
F936
F94D
F9BB
F9DD
F989
F93A
F935
F93D
F929
F92A
F94E
F949
F90C
F913
F9A2
FA07
F980
F8D3
F9F7
FD95
01C2
03F7
03CB
02EA
02C3
0325
033F
02F1
02B3
02AA
029C
028E
02C8
0323
031A
02B1
0291
02F2
0327
02D1
02B1
0361
03CB
0206
FDEC
F9D6
F827
F8C8
F9AF
F98A
F8F2
F8DE
F933
F954
F94B
F97D
F9C6
F9B3
F95E
F947
F974
F97A
F957
F984
F9F7
F9D2
F8CE
F86D
FA9D
FF06
02E1
0406
0333
0293
02F4
036D
034C
0302
0312
032F
02E7
028E
02B9
0333
0342
02E2
02C7
0315
030E
0280
0267
0335
036E
0132
FCF3
F95E
F85F
F92D
F9BF
F95E
F8F0
F91D
F968
F949
F920
F965
F9BC
F99E
F94C
F951
F986
F96F
F936
F972
F9F3
F9D2
F912
F953
FC04
0035
0345
03D5
0319
02D7
0339
035B
0312
0303
035A
0383
0337
02EC
02FE
0318
02DE
02A0
02D4
0324
02F0
028D
02F1
03C4
0315
FFC9
FB7B
F8DB
F8AB
F95E
F977
F925
F938
F99D
F99E
F939
F920
F97E
F9AE
F969
F94B
F9B1
FA00
F9B4
F962
F9B2
FA11
F980
F89E
F983
FD19
0183
03FA
03E3
0308
02FC
036A
0358
02E7
02D8
032D
0346
0310
0309
0343
0344
02ED
02C9
031A
0348
02DD
0281
0312
03CE
02B0
FF0E
FAE7
F8BC
F8D6
F985
F991
F94D
F95E
F99F
F99B
F96B
F975
F9A3
F989
F93C
F945
F9A4
F9B3
F94B
F92B
F9AE
F9FF
F96D
F903
FA9D
FE5D
0221
03D2
0392
0310
0332
0367
031E
02CA
02FE
0367
0369
0326
0324
035A
0357
0325
0339
0388
0379
02F3
02CD
036D
0394
0181
FD71
F9D5
F8A6
F94B
F9CF
F978
F91E
F96B
F9E3
F9D5
F967
F932
F953
F96E
F968
F97D
F999
F968
F911
F92F
F9BB
F9CD
F928
F93B
FBA2
FFD4
034E
0447
037A
02DD
0336
03AE
0380
030C
02FB
033B
0358
034E
0355
0355
0323
0303
0348
03A0
037B
0307
0319
03AE
0349
008C
FC51
F926
F880
F952
F9BD
F958
F909
F947
F994
F986
F95E
F970
F98F
F977
F95B
F985
F9BB
F999
F957
F985
F9E6
F9A6
F8F6
F991
FCAB
00FB
03DB
0432
0357
0311
0388
03C5
036F
032B
035E
0392
0365
0331
0354
037E
0352
031E
0345
036B
0312
02A4
02FD
03BC
030C
FFD5
FB87
F8D9
F8C7
F9BD
F9E9
F950
F908
F957
F991
F966
F93F
F965
F991
F986
F977
F990
F997
F962
F956
F9C6
FA2A
F9C6
F93B
FA58
FDCC
01D3
03FE
03DB
02FD
02CE
033A
0385
0387
0393
03B1
03A0
036B
0365
0385
0367
031C
0331
03A6
03AF
0309
02A8
0344
03C0
022B
FE58
FA79
F8C6
F930
F9F1
F9F1
F99C
F98F
F98E
F941
F902
F938
F98D
F987
F962
F998
F9EA
F9B8
F931
F936
F9E7
FA2D
F96A
F8FA
FAE3
FF0B
02DE
0434
0394
02EF
0312
0353
033D
0335
0387
03CC
03A3
0354
0353
0374
0351
031F
0362
03D8
03AB
02F3
02E0
03C5
03EE
0184
FD32
F9AE
F8BC
F984
FA22
F9F6
F9B7
F9D8
F9ED
F9A5
F962
F978
F993
F971
F96D
F9CB
FA06
F9A2
F92A
F96D
FA0A
F9D1
F8CD
F8EF
FBD7
006D
03C0
0442
033A
02B1
0308
0358
033D
032E
0361
037C
0357
0352
039A
03C6
0383
0334
0353
038E
034D
02E5
034D
0443
03DB
00C1
FC48
F93D
F8DE
F9E6
FA7C
FA32
F9C5
F9AE
F9AE
F994
F991
F9B9
F9C4
F999
F988
F9B1
F9B1
F966
F959
F9D6
FA26
F98A
F8C8
F9BE
FD1D
013A
03B3
03EC
0342
0309
0337
0347
034A
0389
03C3
0393
0334
032B
0362
0359
0319
0334
03B7
03DC
0345
02DC
0390
046E
033E
FF6A
FB29
F915
F94F
FA00
F9F7
F9A6
F9B7
F9E5
F9AA
F94E
F96F
F9EC
FA14
F9D6
F9D6
FA36
FA3E
F9AA
F94F
F9C1
FA2B
F99E
F8FE
FA5C
FE2F
0254
0451
0404
0342
0346
0397
037C
0345
037B
03C9
0398
032A
032B
0388
0391
0325
02E5
031C
034D
0328
033E
03F4
042A
022A
FE1C
FA67
F910
F98E
FA03
F9BE
F97F
F9BD
F9EE
F9A3
F958
F99E
FA26
FA34
F9D4
F9B3
F9F5
FA10
F9E4
FA08
FA85
FA65
F961
F91F
FB78
FFD5
036A
0453
037B
0305
038F
0403
03A6
0326
0346
03AC
03A5
034F
0336
0355
0347
0327
0354
039C
0370
02FE
0323
03E6
03B0
0104
FCB6
F974
F8D0
F9AE
FA17
F9A6
F95A
F9B0
FA1A
FA17
F9E6
F9E5
F9FD
F9F6
F9F0
FA16
FA2B
F9F1
F9C1
FA16
FA89
FA29
F93D
F9A1
FC9F
00FA
0411
04B2
03F8
0385
03B0
03D0
038F
034D
034D
035D
0353
035B
037A
036A
032B
0334
039F
03C3
0341
02D3
034D
03FC
0307
FFC2
FBD2
F985
F959
F9DC
F9CD
F968
F964
F9AC
F9BC
F9A3
F9C9
FA19
FA1F
F9E2
F9E2
FA3A
FA66
FA1F
F9DE
FA0F
FA38
F9BA
F951
FAB3
FE55
0253
0459
0419
0335
030C
0382
03E1
0405
042F
044D
040F
0396
0361
0385
038E
0352
033C
037F
0394
0321
02CE
0361
0420
0321
FF97
FB34
F89A
F89F
F9C3
FA4B
FA09
F9D0
F9E8
F9D4
F964
F916
F947
F9A7
F9C6
F9C3
F9FE
FA5B
FA61
FA0C
F9F4
FA59
FA87
F9D1
F8F4
F9C5
FD19
0175
0455
04A4
0397
030A
0386
0433
0449
0401
03EE
0414
0406
03B7
038D
03B4
03CF
0391
0341
034F
0393
0389
033F
0367
0416
03FC
01A2
FD6F
F9C4
F8A1
F997
FA97
FA64
F99D
F95E
F9B4
F9E0
F9AE
F9AA
FA10
FA51
F9F5
F971
F980
FA08
FA41
F9F6
F9D3
FA3C
FA88
FA13
F9AE
FB1A
FEC0
02B6
04A5
0442
0348
0333
03C5
03FB
03B2
0391
03CD
03D3
035E
030D
0377
042C
0443
03B6
0364
03B3
03EF
0376
02EA
034F
042E
038C
004F
FBF9
F942
F932
FA4E
FAB1
FA21
F9B0
F9EA
FA42
FA2D
F9F1
F9FE
FA23
F9EF
F991
F9A5
FA2E
FA75
FA23
F9E0
FA4E
FADE
FA78
F95A
F96E
FC2C
008C
03E2
04A2
03C0
0321
036D
03DF
03CC
0383
038E
03D2
03D8
03A2
0397
03C9
03D7
039B
037F
03C4
03F6
0388
02D8
02EC
03E9
045C
0299
FEC7
FAF7
F920
F955
FA29
FA76
FA3E
FA07
F9F7
F9E2
F9D9
FA1B
FA8B
FAA4
FA38
F9C6
F9DD
FA49
FA67
FA24
FA26
FAB8
FB1E
FA8F
F9B1
FA64
FD93
01C4
0468
0489
0387
0326
0398
03E6
03A0
0362
03A3
03EC
03A9
033A
0367
0415
044C
03B3
0322
0357
03C5
0377
02BA
02D5
03E3
03F8
0150
FCDF
F99E
F949
FA9A
FB3D
FA9C
F9F4
FA1F
FA83
FA4D
F9CC
F9D6
FA62
FA93
FA1D
F9BE
FA14
FAA4
FAA3
FA3F
FA4F
FADF
FAF2
FA1D
F9AD
FB76
FF75
0364
04F6
0425
02E2
02C5
039C
043C
0422
03C7
03B0
03CA
03C6
03A9
03AF
03CE
03BD
037A
0362
0396
03AD
035A
0312
0378
0414
034C
0030
FBFC
F928
F8E2
F9FB
FA8B
FA21
F9C1
FA19
FA93
FA6B
F9E2
F9C7
FA33
FA7E
FA55
FA26
FA52
FA88
FA62
FA32
FA85
FB0D
FADF
FA10
FA42
FCD1
00E4
0410
04EB
0452
03EC
0429
0444
03D1
036E
03B3
043B
0441
03C8
037F
03B4
03EB
03BA
0368
0370
03AC
0394
032B
031E
03A9
03C6
0214
FE99
FB1B
F972
F9B9
FA77
FA69
F9BC
F960
F9AF
FA1B
FA24
FA06
FA3A
FAA4
FAC0
FA7A
FA51
FA91
FADC
FACA
FA92
FAA6
FAD6
FA8F
FA13
FAD2
FDC6
01D5
048F
04C7
03BD
0367
0424
04CC
0495
040D
03FC
0432
03F9
035F
032B
039F
0403
03C2
0342
0330
0362
033A
02DD
032C
0431
045A
0211
FDE6
FA51
F91E
F9B9
FA4C
FA0A
F9A1
F9C5
FA25
FA22
F9E1
F9FD
FA7F
FAC8
FA87
FA3D
FA6A
FACB
FAD0
FA9F
FADF
FB82
FB87
FA75
F995
FAE6
FEB5
02EB
051C
04F8
0426
040F
047E
048A
0417
03D6
0416
0455
041D
03B3
0398
03BC
03B1
0376
036F
03A2
0389
0303
02D4
03A5
0497
03BC
0051
FBFE
F956
F931
FA25
FA75
F9F7
F9AC
FA11
FA89
FA71
FA08
F9F8
FA58
FAA7
FAA3
FA93
FAB7
FAD8
FABD
FAA1
FAD3
FAFF
FA89
F9BF
FA1D
FCC8
00F2
044A
0542
047F
03C5
03E8
044E
0441
03F8
040A
0462
0463
03E8
0382
039B
03DA
03BF
0377
038B
03EB
03F6
038F
037C
042D
048E
02E9
FF0B
FAF0
F8D9
F915
FA1B
FA85
FA54
FA31
FA3D
FA21
F9E5
FA00
FA83
FAE4
FAC3
FA7B
FA93
FADE
FAC4
FA49
FA29
FAAF
FB08
FA63
F981
FA51
FDB4
021F
0501
0551
0453
03D2
0438
04AA
048A
0427
0408
041A
03FA
03AE
039B
03D3
03F8
03DC
03CE
0407
042A
03C7
0345
038D
0484
0485
0204
FDB0
FA2C
F95A
FA70
FB27
FA72
F95B
F941
FA0D
FAA5
FA91
FA67
FAA0
FADF
FAA3
FA2F
FA1D
FA67
FA7D
FA4A
FA61
FAEF
FB2D
FA8C
FA0B
FB78
FF21
02FD
04B4
0424
0338
0377
047D
0503
04A8
0423
0401
0407
03DD
03B7
03E5
0433
0436
040A
0428
0484
0476
03C1
0332
039A
0453
0398
0096
FCAF
FA31
F9F5
FAC4
FB0C
FA8D
FA17
FA28
FA63
FA58
FA2B
FA37
FA6C
FA7B
FA6B
FA86
FABE
FAA0
FA1B
F9DC
FA6A
FB26
FAF9
FA08
FA1A
FCAB
00E5
0437
0505
042F
039E
03F8
0456
0402
038A
03C1
0472
04B3
044B
03F2
0424
0469
042C
03B9
03C6
0444
0464
03F2
03CE
047D
04DA
031A
FF25
FB26
F957
F9BE
FA9F
FABD
FA76
FA95
FAF6
FAE6
FA64
FA29
FA86
FAE4
FAAF
FA38
FA33
FAA9
FAF1
FABA
FA81
FAAC
FACE
FA57
F9D6
FACF
FDF6
0204
04CC
0551
0477
03B9
03A6
03D6
03EA
03FB
0426
0432
03F6
03C6
0403
047E
049D
0437
03D8
03EA
0410
03BC
033B
0375
0469
0485
023F
FE24
FAA7
F99A
FA67
FB22
FADE
FA53
FA5D
FAC3
FACD
FA7F
FA73
FAC0
FAC7
FA4F
F9FF
FA61
FAF4
FAED
FA87
FAB9
FB91
FBD4
FAD0
F9EF
FB66
FF57
0342
04C1
0416
0368
03E6
04BC
04B6
03FF
039E
03E3
0436
0437
0445
04A1
04CF
045B
03BF
03C7
044B
044E
0385
02FC
03A0
0491
03CE
00A0
FCB8
FA71
FA62
FB1F
FB33
FA95
FA25
FA50
FAB9
FAEF
FAE5
FAB5
FA5C
F9FC
F9FD
FA8E
FB30
FB28
FA84
FA26
FAA0
FB57
FB47
FA96
FACB
FD1A
00CF
03D9
04DA
0454
03BA
03C8
041F
0438
0428
0442
0480
0495
0477
0465
046A
0447
03F1
03D1
042F
049B
046B
03C1
038E
0430
047D
02D4
FF27
FB6F
F9BF
FA37
FB3B
FB76
FB10
FADA
FAF5
FAD7
FA53
F9EE
FA12
FA6A
FA76
FA53
FA7D
FAEB
FB08
FAA3
FA5E
FAB5
FB1C
FAC2
FA1E
FAF0
FE28
025C
04FB
0502
03D8
035D
03D5
0435
03F1
03A7
03FF
04AC
04FC
04E6
04E0
04F4
04AE
040A
03B7
0414
047D
043A
03BC
040F
0506
04CE
0207
FDC2
FAA4
FA07
FAC9
FB16
FAA4
FA75
FAFD
FB77
FB2F
FA8A
FA4E
FA6E
FA49
F9DA
F9DD
FA99
FB3A
FAF6
FA47
FA49
FB03
FB3E
FA66
F9DB
FB8F
FF83
0368
0512
04A4
03F5
0425
04A4
047E
03DA
0398
03FE
046C
0465
043F
0473
04CB
04B1
0433
0408
047C
04ED
04B3
0434
0448
04AF
03DB
00CD
FCAC
F9DF
F999
FAC6
FB86
FB3C
FAA8
FA81
FA9F
FA9E
FA9A
FAD6
FB1E
FB04
FA98
FA5A
FA76
FA8E
FA6D
FA78
FAF1
FB39
FA8B
F982
FA01
FD17
016C
046C
04EC
0413
0399
03EE
045E
0483
04B5
051C
0537
04A2
03DC
03AB
0406
043A
0406
03F4
045E
04B9
045E
03B5
03DC
04F3
056A
0392
FFAF
FBE3
FA15
FA38
FAD8
FADE
FA6E
FA38
FA66
FA91
FA69
FA21
FA19
FA61
FAB8
FAED
FB0C
FB33
FB48
FB15
FAA0
FA48
FA5D
FAA5
FA9A
FA37
FA61
FC23
FF6A
02CB
04B5
04E1
0461
044D
04B5
04F6
04C7
048C
04AE
04FF
04FB
047D
03E3
0391
038F
03BF
0424
04BE
0533
0502
043E
03B9
042C
0524
0517
02E0
FF0D
FB8E
F9EF
FA14
FAAE
FAC3
FA73
FA54
FA7F
FA87
FA41
FA1B
FA7F
FB27
FB67
FB0C
FA9A
FA8D
FAB8
FA9F
FA4F
FA5F
FB07
FB8C
FB1A
FA0D
F9FE
FC30
0012
03A4
054B
0520
0471
0446
0496
04CD
04AC
0478
047B
04A0
04AA
0488
0467
0469
047B
0480
047E
0486
0480
043A
03CD
03BB
0467
0551
0526
02E6
FF12
FB7A
F9BA
F9DE
FAA7
FAF4
FABB
FA95
FAC0
FAEA
FAD2
FAB0
FAD4
FB14
FB05
FAA5
FA7D
FAE4
FB78
FB8D
FB1B
FAC9
FAFF
FB3C
FAC3
F9E1
FA18
FC97
00BD
045F
05BF
0514
0406
03E2
0481
04F4
04C9
0461
0439
0448
043D
041B
042D
0473
0485
0428
03BF
03D5
0454
0497
0457
042A
04B0
0563
04C2
01EA
FDD4
FA9B
F991
FA35
FB0A
FB2A
FAD5
FAAE
FADA
FAFE
FADF
FAAD
FAAC
FACD
FAD0
FAA6
FA98
FADF
FB49
FB65
FB13
FABD
FACA
FAFC
FAC2
FA35
FA7D
FCBD
0094
0415
0586
050A
0442
045A
04F0
04FF
0465
03FA
0450
04EB
0503
0496
0449
0463
0470
040E
03A7
03E3
04A5
050F
04AF
042B
0463
0516
04D1
027E
FEBE
FB77
FA08
FA34
FAB8
FAC5
FA8D
FA9C
FAF5
FB1F
FADF
FA89
FA8E
FADD
FB0D
FAFE
FAFE
FB41
FB72
FB23
FA86
FA58
FAE0
FB6B
FB20
FA58
FA9D
FD11
00F9
0448
0595
0543
04BC
04CB
0516
0506
04B1
04A6
0506
0550
0509
046B
0419
045A
04CD
04FA
04DE
04CB
04D6
04BC
0465
0441
04B7
054B
04B3
021B
FE46
FB20
F9FF
FA7C
FB1B
FAED
FA51
FA1C
FA73
FABF
FA96
FA41
FA41
FA9C
FADE
FAC8
FA98
FA9E
FABF
FAAD
FA78
FA8E
FB0E
FB62
FAF3
FA2D
FA80
FCFB
00EF
0451
058E
04F6
0428
0442
04F1
053B
04D5
045E
0469
04BF
04D0
0486
0450
0473
04A4
0489
044B
0455
04A2
04B1
044C
03FF
0461
0505
0484
01F0
FE0F
FAD7
F9A4
FA19
FAC8
FAC3
FA4C
FA23
FA79
FAD4
FAD1
FAA1
FAAE
FAF7
FB17
FAD8
FA8B
FA96
FAE6
FB0B
FADE
FAC1
FB03
FB47
FAFE
FA7C
FB1B
FDD5
01DB
0501
05CD
04E2
041B
047D
055D
0595
0504
0482
049A
04EB
04D8
047C
0468
04BB
04F0
04AB
0450
0473
04EA
04F5
045F
03F7
0483
0565
04DD
01E9
FDA8
FA7A
F9BF
FAAA
FB64
FB02
FA31
FA08
FAB1
FB63
FB7A
FB24
FAEE
FB03
FB18
FB08
FB06
FB37
FB4F
FAFB
FA7B
FA76
FB11
FB83
FB14
FA52
FADF
FDAB
01AA
04AF
058D
050B
04AF
0503
0552
04F8
0447
0400
044F
04B1
04C7
04C3
04EA
0509
04C0
0431
03F5
045A
04DC
04CB
043B
0404
04A7
055E
04A8
01CF
FDD9
FAC6
F9CC
FA5A
FAF1
FABB
FA2F
FA28
FABB
FB32
FB12
FAB2
FA99
FAB3
FA81
FA08
F9F0
FA8F
FB3F
FB2E
FA8E
FA68
FB15
FB92
FADF
F9C0
FA50
FD9A
0218
051E
0586
0482
03E5
0440
04DA
0509
04EE
04EB
04FC
04E6
04BC
04CA
050C
051F
04CB
0464
0465
04C9
0502
04B1
0434
044E
0528
05C7
04BD
0197
FD93
FABD
FA27
FB07
FBB5
FB6B
FACA
FAB7
FB21
FB3E
FAC1
FA42
FA5F
FAE2
FB1C
FAEC
FAD6
FB1E
FB4D
FAEC
FA60
FA72
FB1C
FB62
FAAF
F9FB
FAFD
FE37
0227
04B7
052D
048B
042B
0469
04C2
04C8
04AC
04C9
0519
0543
0520
04EE
04EE
0506
04E5
0489
0456
049A
050C
051A
04B7
048F
0517
0595
048A
0160
FD65
FABF
FA56
FB1C
FB76
FAF8
FA79
FAAB
FB35
FB5A
FB06
FAC4
FADA
FAEB
FAAC
FA71
FAB7
FB51
FB80
FAF9
FA68
FA9F
FB74
FBD6
FB33
FA74
FB42
FE41
022B
04E6
0568
0483
03D8
042F
04F5
053F
04E8
0489
0492
04C2
04AF
0473
047B
04CF
04F3
04A4
044D
046E
04D0
04CD
045D
0454
0527
05CE
048B
00F8
FCD1
FA58
FA25
FAEF
FB42
FAED
FA9E
FAB4
FAEA
FB06
FB3A
FBA4
FBE5
FB88
FAC5
FA55
FA91
FB00
FB00
FAA6
FA9A
FB23
FBA8
FB5E
FA69
FA09
FB85
FEE1
02AC
0523
059B
04E2
0458
049E
0534
0549
04BD
0435
0442
04BB
0509
04E4
0497
0481
04A1
04BE
04CD
04EC
0506
04DB
047E
0474
04FF
0557
0413
00BB
FCAF
FA1E
F9ED
FAF7
FB75
FAEA
FA51
FA91
FB54
FBA4
FB41
FAD8
FAF3
FB3A
FB19
FAB3
FAB5
FB45
FBB4
FB73
FAEF
FAF2
FB6D
FB72
FAAB
FA3F
FBCA
FF61
0333
0542
0542
048C
046C
04F4
0561
053F
04CC
047C
0469
046C
046D
047F
04A6
04C8
04D6
04E5
0503
0508
04B7
041C
03B7
0413
0504
0566
03F7
009F
FCD8
FA82
FA4A
FB31
FBBC
FB66
FAC6
FA8D
FABA
FAED
FB0A
FB45
FB92
FB93
FB2B
FACC
FAF4
FB6F
FB90
FB25
FAD8
FB50
FC29
FC46
FB55
FA9B
FBD4
FF4C
034D
05AF
05CF
04E3
046F
04C9
052D
0504
04A0
049E
04F7
0514
04B7
0465
04AE
054A
0565
04C1
0412
0415
048C
04AA
044C
043F
04F8
0576
0416
008E
FC9E
FA6F
FA73
FB47
FB7B
FB03
FABD
FB13
FB87
FB80
FB16
FAC5
FAC2
FADF
FAFF
FB3C
FB8D
FB93
FB19
FA8D
FAA3
FB65
FBE3
FB3F
F9EE
F9A9
FBCF
FFDE
03B8
0587
0541
045C
0421
048F
04D9
049D
0447
045D
04C8
050F
050F
0513
0537
0522
0497
040C
043F
052F
05DF
0586
04A8
048A
0572
05EA
0428
0030
FC1D
FA24
FA8E
FBBF
FC22
FB9E
FB20
FB38
FB8B
FB8F
FB54
FB43
FB69
FB5A
FAEB
FA93
FAD8
FB80
FBC3
FB55
FAD5
FAF3
FB6A
FB4E
FA7B
FA38
FC04
FFC6
039B
059A
058A
04B5
044C
046C
048F
0482
0481
04A9
04B8
0482
044B
0472
04DC
050A
04C7
0477
0495
04FD
0508
0469
03BB
03E3
04E2
0567
03ED
005A
FC53
F9DE
F99C
FA75
FAF9
FAC7
FA89
FAC5
FB32
FB45
FAF9
FAC4
FADE
FB09
FB0B
FB09
FB2E
FB43
FAFF
FA9C
FABB
FB6F
FBE8
FB6B
FA82
FAAF
FCDE
0051
0354
04D9
0529
0525
0546
0566
054A
0505
04CF
04C1
04C1
04B4
049C
049A
04B9
04D9
04CD
04A5
04A7
04E7
050C
04B7
0430
043D
050B
056B
03D1
002B
FC59
FA63
FA7D
FB2E
FB30
FAB2
FA90
FAF5
FB44
FB27
FB03
FB3F
FB91
FB77
FB08
FADA
FB2D
FB97
FBA1
FB56
FB20
FB38
FB75
FB84
FB34
FA9A
FA3F
FB0C
FD91
0126
0429
056E
0546
04EA
04FE
0524
04E4
0478
046A
04C0
0500
04EF
04D9
04FD
0526
0519
04FC
050E
0522
04EA
0483
0461
049E
04D2
04CB
04E7
0546
04FA
02CC
FEF8
FB7B
FA27
FACA
FBB7
FBD0
FB67
FB3C
FB5F
FB66
FB45
FB52
FB8D
FB81
FB05
FA95
FAAC
FB20
FB77
FB8E
FB8C
FB78
FB45
FB33
FB87
FBE1
FB78
FA72
FA6C
FCED
0144
04D0
05B3
04BF
0424
04C7
05A4
0596
04D7
0474
04CE
0559
0589
0566
0533
04FF
04CE
04C7
04E7
04E2
049D
0479
04BE
0509
04E2
04A8
052D
0633
05F8
0316
FE8D
FB15
FA49
FB22
FBA0
FB30
FAC3
FAFE
FB61
FB42
FAD4
FAB1
FAE0
FAF2
FADA
FB0A
FB9C
FBFF
FBD0
FB6E
FB5C
FB76
FB52
FB07
FAF5
FAF1
FA6D
F9BE
FA6C
FD8C
01FF
0539
05E2
0517
04B7
0535
05A5
0569
04F9
04F2
0534
0545
0513
04E7
04CE
049B
0465
047D
04D3
04EC
04B0
04A8
051C
0572
0509
0460
0484
0542
04D7
01FD
FDCF
FAD9
FA48
FAE3
FAF2
FA53
FA18
FAAE
FB55
FB5B
FB00
FAE5
FB25
FB69
FB8B
FBA5
FBA6
FB56
FAE1
FAC8
FB1B
FB4B
FB10
FAF8
FB7C
FC04
FB9E
FAB3
FB1E
FE0C
0248
0556
0617
059E
0567
058E
0555
04AF
045D
04B0
0515
04F9
049A
0489
04C6
04DA
04A5
048A
04BA
04E7
04D7
04C0
04C7
04A0
042B
040B
04D3
05B6
04D0
014D
FCC2
F9CC
F972
FA6E
FB14
FB17
FB25
FB7F
FBAF
FB76
FB2F
FB30
FB4E
FB41
FB2C
FB51
FB87
FB6C
FB13
FAF2
FB27
FB45
FB1E
FB24
FB9E
FBEB
FB65
FACD
FBEB
FF6B
03A4
0624
063F
0568
0524
056C
0568
04F9
04BF
04ED
0501
04AF
0471
04C2
054E
055D
04E0
048C
04D9
0572
05C1
05A3
0539
0497
0401
040C
04DD
0554
03CC
0012
FC10
FA00
FA24
FAD4
FAB7
FA39
FA75
FB6F
FC1E
FBDE
FB2A
FACD
FAF1
FB3E
FB6E
FB75
FB43
FADD
FA93
FABC
FB2A
FB56
FB32
FB48
FBBB
FBCC
FB04
FA86
FC38
005B
04B8
06BC
0631
0517
050B
059D
0588
04AB
040E
044F
04EC
0527
04FC
04DE
04FC
052B
054E
0563
053F
04BB
042E
0432
04C0
0510
04B7
0460
04C3
052A
03E7
006F
FC61
F9FD
F9D2
FA95
FAFC
FB05
FB34
FB74
FB4F
FAEB
FAE5
FB5B
FBB1
FB76
FB08
FB00
FB5E
FBB1
FBCF
FBEE
FC10
FBEB
FB8D
FB81
FBE6
FBFC
FB48
FAD3
FC5F
0030
0445
0641
05DA
04C9
049B
0531
0594
056A
0517
04E2
04B6
049B
04CB
053A
057C
054C
04E8
04A8
0482
044A
0434
0488
04ED
04AF
03F4
03D8
04CF
0568
03A5
FF89
FB87
F9F3
FAA4
FB94
FB77
FAE1
FAD7
FB46
FB75
FB4A
FB50
FBA8
FBBE
FB38
FA96
FA94
FB37
FBDF
FC17
FBF3
FBBB
FB9B
FBBC
FC21
FC4E
FBA2
FA79
FA7F
FD1C
019C
057F
06DE
062A
053F
052F
0588
0586
052C
04EA
04CD
049F
047A
04AD
0518
053B
04E3
0472
0443
043A
0422
0421
0464
0491
0432
03BB
0441
05B1
0608
0346
FE12
F994
F859
F9DA
FB76
FB79
FA7C
F9F6
FA54
FAE4
FB0E
FAED
FADB
FAFB
FB41
FB9D
FBE9
FBFB
FBE5
FBE5
FC00
FBEA
FB86
FB40
FB79
FBBF
FB43
FA59
FABA
FDAE
0230
05A8
068E
05C6
053A
05A0
0634
0637
05E4
05BD
05AC
0556
04E3
04C8
04FF
04F7
046C
03D1
03B3
040F
0474
04A5
04AF
048D
0440
0438
04F8
05FE
0598
0293
FDF1
FA51
F969
FA80
FB87
FB63
FAA1
FA44
FA83
FAEC
FB33
FB59
FB5C
FB29
FAE1
FACC
FB0E
FB8C
FC1D
FC8C
FC82
FBCE
FAED
FACE
FBAC
FC63
FBB7
FA52
FAAE
FE4F
0395
0717
0729
055D
0465
051B
062F
0647
0583
04CF
0494
049D
04CD
0531
0591
057C
04F6
0494
04C9
0551
0592
0557
04DD
045F
0404
0421
04F2
05B6
04D6
0187
FD23
FA26
F9C5
FADB
FB6E
FAD2
F9F7
F9F2
FAC6
FBB2
FC15
FBD0
FB26
FAA2
FAC7
FB81
FC09
FBBC
FAF2
FA9C
FB0A
FB8D
FB85
FB3F
FB54
FB8A
FB2E
FAA2
FB90
FEF3
0367
0655
06B1
05D2
0579
05CF
05C8
0501
0451
047F
0535
059F
057C
0524
04CB
0466
041F
0444
04BE
0509
04E2
04A3
04B4
04E4
04D4
04B5
04F5
0521
03EA
00C9
FD0F
FABA
FA60
FAEA
FB39
FB4E
FB9C
FBEB
FB9D
FAD3
FA6E
FAD4
FB57
FB3F
FAD7
FAE4
FB7A
FBF1
FBEC
FBC1
FBC7
FBD8
FBC4
FBCD
FC24
FC4A
FBB1
FB04
FBF2
FF2B
032A
05A6
05EF
053A
04CA
04A5
0446
03DD
0418
04FA
05AA
058C
0505
04CE
050E
056E
05A9
05A2
053B
0498
0451
04CC
0562
04F2
0386
02C1
03DC
0591
0513
0168
FCD6
FA6A
FAB2
FBB9
FBD6
FB57
FB57
FBE1
FC16
FB9D
FB11
FAF3
FB01
FAE1
FACE
FB19
FB72
FB55
FAE5
FABC
FB04
FB57
FB8D
FC05
FCC3
FCED
FBE8
FAC7
FBAA
FF49
03BD
065B
064E
04F8
0408
03F9
0455
04A6
04CC
04CA
04CA
0524
05EC
0682
061B
04E1
03F5
0411
04B2
0500
04FD
0533
0581
0530
0445
03D9
048C
051E
039F
FFF9
FC5D
FAD2
FB0F
FB66
FB13
FACB
FB2A
FBB3
FBA6
FB23
FADC
FAFB
FB1B
FB2A
FB94
FC53
FC92
FBCF
FABF
FA7A
FB11
FBA0
FBB7
FBD2
FC4A
FC8B
FC04
FB81
FC9F
FFBE
033E
0538
057A
0549
058A
05EC
05CF
053C
04C2
04B2
04E8
0525
0539
04F8
046D
0408
0443
04DE
050B
048C
0425
0492
056D
05B8
0553
0516
0552
04F3
02C0
FF31
FC20
FABC
FA76
FA4F
FA50
FB05
FC1A
FC74
FBB3
FAC6
FAA7
FB1C
FB4B
FB25
FB66
FC4A
FD0B
FD03
FC95
FC62
FC2F
FB55
FA15
F98F
FA35
FB0F
FB28
FB2E
FCDA
009F
04CB
073E
077D
06A6
05CB
0527
04AC
0489
04D7
053A
0533
04BD
0442
040C
0418
0457
04BD
04FF
04C3
044A
045C
0543
062E
0632
0596
0566
05C2
053F
029B
FE8B
FB34
F9E1
FA00
FA67
FAC3
FB3F
FB8C
FB2E
FA90
FACE
FC2C
FD6C
FD43
FC01
FB21
FB5A
FBDC
FBA7
FAD7
FA30
FA07
FA37
FABF
FBA9
FC64
FC2B
FB55
FB93
FE2E
023D
0562
064B
05CE
0568
055C
04FA
0419
0369
036C
03E1
045D
04DE
056E
05B7
0564
04D6
04C6
0542
0599
0577
0555
0586
0582
04DC
0448
04A2
04EB
0276
FBDC
F349
ECE9
EAF3
EBF4
ED1F
ED57
ED73
EE4F
EF8D
F038
EFD1
EE90
ED2B
EC81
ED0E
EE50
EF08
EE8A
EDA1
EDA2
EEAF
EF92
EF7D
EF1F
EF7E
F067
F0DD
F0AE
F0AD
F139
F17D
F0A4
EF44
EEAD
EF21
EF90
EF43
EECB
EEE0
EF37
EF30
EF0E
EF66
EFC1
EF1B
EE16
EF73
F52A
FD62
0397
0514
0359
01B5
0186
01BB
014A
00A7
00AC
0132
016C
012F
0117
0185
021F
0270
0282
0297
02B9
02DA
030E
0344
0324
028F
01FC
01D6
01DF
01AC
0197
0288
0486
0639
066B
05AF
059D
069F
077A
074B
06DA
0736
07FC
0824
07EF
0876
0911
06BD
FF7C
F5A9
EE78
ECBF
EE79
EFDF
EFB2
EF6E
F035
F140
F16F
F105
F0F7
F156
F14C
F07F
EF99
EF41
EF4E
EF49
EF34
EF3E
EF36
EEDB
EE75
EE80
EEE7
EF26
EF1B
EF2E
EFA0
F021
F05C
F083
F0DE
F11C
F0BC
F009
EFDB
F047
F06A
EFEF
EFC2
F075
F0D8
EF9B
EE3D
F0A2
F8AE
031B
0A22
0B3E
0933
081F
08FA
09D5
094C
081F
0790
07AE
07D3
07E8
0848
08D7
08FC
0898
0837
081E
07F1
078B
0782
0838
08F5
08C6
07F2
07BA
0889
0939
0875
065F
044D
032F
02D1
02A3
0281
0277
026D
0277
02DD
0370
0367
029B
0249
0387
0503
0379
FD49
F4FE
EF3C
EE25
EFB5
F0B7
F03E
EF8C
EFA2
F02A
F07E
F09A
F0BA
F0CF
F0C4
F0E7
F17C
F230
F280
F28F
F2E8
F36D
F34B
F252
F17C
F18E
F1F2
F1A7
F0EA
F0F2
F214
F32F
F342
F2CE
F2EF
F399
F3BC
F310
F293
F2F1
F381
F37D
F338
F33C
F2F3
F1A8
F0A5
F2C5
F911
00B8
0589
0636
0519
04D8
0590
05D7
054A
04D5
050B
056E
056F
0522
04C4
0447
03AC
035C
03A0
0415
0429
0412
0478
0545
0598
052E
04E2
0542
057C
04AB
039E
041C
066D
08C0
096B
08E4
08BB
0942
096D
08D4
0868
08C2
0921
0901
0974
0B52
0C85
0936
0067
F62B
F010
EFAB
F1CA
F2CD
F24D
F20F
F2CC
F37F
F35F
F2FD
F32A
F3BB
F3EE
F392
F328
F30B
F2F8
F281
F19E
F0BB
F05C
F0D8
F1F9
F2E1
F2BB
F1D2
F15F
F206
F303
F346
F2ED
F2E4
F35D
F389
F300
F28B
F2D6
F320
F259
F13A
F19D
F36D
F3FE
F1DC
EFFD
F33D
FC73
06BF
0C74
0CAC
0AF7
0A6F
0AEC
0B00
0A9E
0A95
0AB7
0A31
093D
0912
09FB
0AC5
0A6B
0983
0957
0A1F
0AF4
0B3F
0B42
0B2E
0AB1
09EA
09BB
0A89
0B6E
0B6D
0ABC
0A11
093A
0793
05A8
0505
05FB
06C8
05EC
047E
04A6
062D
069F
053C
0486
0653
0801
0500
FCD5
F455
F04F
F0A1
F1C2
F1BB
F197
F255
F2EF
F261
F1A6
F21A
F308
F2A9
F11B
F078
F1E5
F3F8
F4C5
F453
F3FB
F423
F3F3
F33F
F323
F427
F51B
F4CE
F3E7
F3DC
F4BA
F53F
F4E9
F492
F4E0
F535
F4E9
F490
F51D
F624
F655
F5A5
F57B
F643
F671
F52C
F4BD
F860
FFD4
06C6
0954
07FA
062F
0615
06DC
0722
070B
0753
07A2
0726
0625
05B2
060D
0668
0645
0621
066D
06B7
067D
062A
0670
06E5
0669
0516
047D
056C
0696
066A
056F
0594
0773
099E
0AB5
0B0F
0B9E
0C29
0BD1
0ADF
0A8F
0AFF
0AF9
0A45
0A7D
0C39
0CA4
080F
FEED
F654
F2D6
F3EF
F5A0
F58C
F4C6
F4E8
F57B
F54C
F4AD
F4D3
F5BF
F642
F5D4
F515
F482
F3D1
F2EF
F2A5
F374
F47C
F481
F3CA
F3C0
F4A7
F517
F440
F359
F3BF
F4D3
F4FE
F428
F39F
F3D3
F3B3
F2BE
F23D
F356
F4E8
F4E9
F398
F337
F456
F4B0
F31E
F2C5
F7E0
01D9
0AF9
0E7E
0D4A
0B96
0B8D
0BEF
0B69
0AE1
0B91
0CBE
0CDC
0C01
0BA4
0C4B
0CF4
0CDD
0C8F
0CB7
0CFE
0CAC
0BFE
0BE7
0C97
0D2B
0CF9
0C67
0C1A
0BFA
0BA5
0B2F
0ABB
09F8
08B6
07AD
07B2
0857
0843
071D
062D
067D
0726
06B1
05A6
0600
07A2
072C
01E0
F9B9
F3DF
F306
F4E6
F5AA
F472
F33F
F35C
F3CF
F383
F32F
F3FC
F560
F5C1
F4CB
F3DA
F3F7
F4A2
F4F4
F514
F5B4
F6A7
F6F6
F65C
F5C3
F5E4
F64B
F63E
F5E7
F5DC
F604
F5CD
F53A
F4F5
F54F
F5DE
F63A
F684
F6DD
F6E8
F67D
F654
F6F1
F747
F5F3
F432
F5C4
FC89
0542
0A6D
0A21
0797
06C1
07EA
08C1
084F
07EA
0877
08DF
0826
075A
07F2
095A
09BA
08BC
07D8
07F6
0834
079A
06DC
0749
0897
0927
0873
07B5
07D1
07EB
071A
0644
0702
0946
0B6D
0C6B
0CAC
0CD6
0CD5
0C91
0C94
0D1E
0D3F
0C2D
0B19
0BF2
0DE1
0CE2
0655
FCD0
F5C7
F3D8
F4EC
F5C0
F58F
F586
F618
F676
F655
F688
F761
F7D5
F710
F5EA
F5B1
F635
F639
F576
F4ED
F52F
F571
F4D9
F3F2
F3EA
F4D0
F572
F51E
F482
F483
F500
F555
F56C
F584
F576
F50F
F4D7
F57A
F67D
F674
F508
F3D3
F45C
F5B9
F5B7
F477
F550
FB07
03FC
0B80
0EB1
0EC0
0E6C
0E9D
0E69
0D6D
0CAD
0CEB
0D7F
0D75
0D12
0D41
0E0E
0E9A
0E6F
0E07
0DDC
0DB4
0D38
0CBE
0CE1
0D7E
0DBE
0D43
0CA8
0CAE
0D4C
0DE8
0DF5
0D1D
0B59
0958
084B
089C
0936
08B9
0756
0697
0730
07EF
07A2
072A
0811
094E
076B
00E4
F8EF
F453
F430
F571
F531
F3F3
F3D9
F532
F646
F61C
F5A7
F5E9
F650
F5EE
F527
F504
F586
F5C4
F585
F590
F656
F743
F799
F76F
F751
F75F
F755
F73D
F762
F78D
F744
F6CB
F700
F7C9
F7DE
F6BD
F5C9
F669
F7D9
F835
F751
F6F3
F7D3
F817
F64A
F4CB
F7F4
0073
0969
0D6E
0C2C
0996
08B1
090E
0916
08BA
08D8
094A
0920
085B
0819
08C7
094D
08B5
07AD
077F
0837
08D1
08DF
08F9
097D
09E3
099B
08FA
08BD
08FA
0923
08F3
08C2
08EC
0985
0ABC
0CBC
0ECD
0F71
0E2A
0C94
0CB4
0E61
0F77
0EE0
0E21
0EE6
0FB3
0CD0
04EC
FB86
F59F
F4C6
F65A
F73F
F6E8
F685
F697
F685
F614
F5FF
F6C9
F7DA
F84C
F7FD
F754
F672
F55B
F48A
F48D
F510
F509
F423
F365
F3FE
F5A3
F6D4
F69C
F583
F4A5
F495
F549
F66A
F739
F6E0
F587
F4A2
F55D
F6F5
F791
F6B2
F5CF
F60F
F67C
F5BE
F531
F83C
FFF6
08E3
0E4C
0F1B
0E26
0E35
0F40
0FCD
0F7B
0F43
0FB3
1033
100E
0F61
0EA6
0E15
0DD4
0E1F
0EA8
0E96
0DAF
0D01
0D89
0EB6
0F18
0E53
0D78
0D55
0D68
0D06
0CBF
0D82
0EA7
0E46
0BCE
090F
07EC
0814
0804
076D
0733
0775
073C
0673
06B3
08C9
0A4F
077C
FFD2
F78B
F37C
F440
F67E
F72F
F658
F58A
F557
F50C
F456
F3FD
F4CC
F653
F740
F6DB
F5CC
F570
F679
F847
F973
F920
F7DA
F70D
F773
F852
F871
F7A5
F6EE
F71F
F7D1
F7F9
F749
F692
F6B4
F79B
F874
F8B4
F885
F84E
F83F
F86D
F904
F9DD
FA34
F943
F75E
F606
F664
F7EA
F8DB
F853
F736
F6E5
F76D
F7BB
F761
F747
F817
F8D1
F7F6
F61D
F64A
FAE1
02A2
095B
0BDD
0AC5
092A
091E
0A11
0A79
0A0D
09D5
0A75
0B39
0B0F
0A00
0921
0937
09D5
0A09
0998
0917
0912
0987
0A51
0B88
0D26
0EAD
0F8A
0FB7
0F9D
0F6A
0EEF
0E36
0DE4
0E79
0F83
1000
0F9E
0F06
0ED6
0EDD
0EA7
0E42
0DFA
0DDC
0DDE
0E4F
0F5A
1046
0FED
0E45
0CD6
0CFB
0E2E
0ED6
0E81
0E18
0DD5
0C8D
09DA
07B6
0830
09F7
08EB
02E6
FAB1
F541
F478
F5E8
F681
F5E2
F57F
F5D8
F604
F576
F4D7
F4ED
F59F
F65D
F6DE
F714
F6DE
F645
F5CE
F60D
F6C7
F729
F6EF
F6D4
F777
F84A
F845
F75E
F6AC
F70C
F829
F906
F912
F88A
F801
F7D1
F7FE
F84C
F861
F814
F7BE
F807
F918
FA22
FA15
F8E3
F7B2
F79D
F873
F8FF
F87F
F799
F77C
F84C
F8E2
F85E
F77C
F7A3
F8C8
F929
F7B3
F628
F7D8
FDEE
05A2
0AB3
0B6B
09D1
08EC
09AC
0ACB
0AF3
0A3E
09AC
09D0
0A65
0AD3
0ABD
0A31
0995
096A
09EA
0ABC
0B26
0AB8
09D5
0952
0993
0A2A
0A72
0A5F
0A65
0AB4
0ADB
0A6D
09DA
0A35
0BEF
0E18
0F45
0F1D
0E95
0EA0
0F16
0F30
0EA3
0DE1
0D79
0DA7
0E5A
0F4B
0FEB
0FB1
0EC1
0E00
0E17
0E95
0E8C
0DEF
0D85
0D8E
0D5F
0CC6
0CD1
0E08
0E80
0B1D
0360
FAE3
F61A
F5E6
F74F
F766
F635
F583
F5F2
F689
F674
F5F8
F5A1
F574
F560
F5B2
F685
F733
F6FA
F62D
F5EA
F68B
F70F
F695
F5C7
F60C
F77C
F896
F82C
F6E4
F644
F6C1
F75F
F73B
F6B3
F6AA
F737
F79E
F781
F768
F7DB
F893
F8F3
F8FB
F923
F963
F926
F862
F803
F8B9
F9CD
F9E3
F8E6
F843
F8F2
F9FE
F9DD
F8B1
F808
F85C
F85B
F774
F7DD
FC7E
04F4
0D0E
10DF
107A
0F15
0F11
1006
105D
0F87
0DF9
0C2B
0A7E
09AA
0A1F
0B1B
0B42
0A3C
0915
08D4
093B
0970
095F
09C1
0ACC
0BB4
0BB9
0B26
0AB8
0A88
0A30
09BD
09C1
0A5D
0AE8
0AC4
0A32
09EE
0A25
0A44
09D3
0937
093D
0A13
0B19
0BCF
0C73
0D8A
0EF1
0FD4
0FA7
0ED7
0E52
0E60
0E63
0DD8
0D2D
0D1F
0D9F
0E0B
0E6B
0F5D
1049
0EAB
0877
FF48
F7E0
F5BD
F7A0
F953
F87A
F691
F615
F733
F829
F801
F790
F7C8
F848
F822
F73F
F660
F603
F60A
F65C
F715
F7E3
F7F2
F6FE
F5F7
F5F3
F6B6
F709
F670
F5D5
F621
F6EF
F72F
F6C4
F697
F718
F786
F72E
F6B0
F722
F852
F8D3
F7FD
F6F7
F719
F804
F84A
F7B7
F793
F874
F911
F833
F6DC
F713
F8DC
F9FB
F93A
F865
F996
FB9B
FB4D
F8B3
F86E
FE68
087A
1049
1223
1031
0EBA
0F1A
0FA9
0F49
0EE1
0F52
0FE3
0FA2
0F05
0EFB
0F43
0EF9
0E47
0E31
0EB8
0E92
0D09
0B23
0A32
0A00
0978
08AC
08E8
0A6C
0B8D
0AE7
0965
08F5
09CF
0A73
0A13
09A1
0A17
0ADB
0AA9
0992
08E4
093C
09B4
0975
0918
09AC
0AD8
0B2E
0A24
08D4
0873
08E0
0940
0989
0A9D
0CB5
0E81
0E88
0D38
0CBC
0E35
0FA9
0D8A
0685
FD78
F718
F5B3
F783
F91A
F8EC
F810
F7FA
F882
F86D
F747
F5FB
F5C0
F6E1
F89F
F9E5
FA0D
F943
F857
F7FF
F839
F868
F833
F801
F850
F8CE
F89E
F7A9
F6FD
F778
F887
F8C8
F7CC
F695
F63A
F6A6
F700
F6EB
F6DB
F730
F796
F793
F752
F756
F796
F76A
F68D
F5B0
F5B6
F68E
F751
F76D
F74A
F78C
F80D
F821
F7C3
F7C5
F87A
F8E5
F836
F7DD
FAC8
01EA
0A54
0FAB
1076
0F22
0EBE
0FB9
1077
1030
0FD8
1043
10C7
1068
0F68
0EBD
0E8D
0E37
0DA8
0D9D
0E6F
0F63
0FB0
0F8C
0FA2
0FD5
0F76
0EAD
0E87
0F3C
0F70
0DFB
0BC4
0ABB
0B47
0BD7
0B1E
09BF
092B
098E
09C1
091C
086B
08A6
098D
0A22
0A22
0A2D
0A9A
0AED
0A9E
09E0
0956
093B
0939
08FB
0894
083F
0804
07E5
083B
095C
0A88
09BE
0562
FE59
F7FD
F560
F67E
F87A
F8B3
F748
F639
F69F
F78C
F7AE
F709
F690
F6BE
F748
F7D5
F854
F8A4
F894
F84B
F845
F88E
F889
F7DF
F759
F7F0
F932
F991
F88A
F780
F7D1
F8F2
F95D
F8C3
F835
F84A
F848
F78B
F6CA
F70B
F7EB
F80B
F730
F6B0
F756
F809
F776
F63A
F613
F750
F852
F7DB
F6BB
F67F
F74C
F7EB
F7C7
F7AA
F823
F83E
F6F2
F56F
F6BA
FC6B
0464
0A68
0BF9
0A6A
0922
0A2E
0CAF
0E89
0EEB
0EC8
0F2B
0FEC
103C
0FEC
0F90
0F8F
0FA9
0F86
0F53
0F69
0FA8
0FAF
0F96
0FD5
1055
104B
0F6C
0E9E
0EE5
0FF1
106B
0FAE
0E8A
0E35
0EE0
0FB8
0FF8
0F95
0ED9
0DE6
0CC9
0BA6
0A9A
09BD
0959
09C1
0AA0
0AF9
0A48
0955
0946
0A05
0A4A
0964
0850
086A
097F
09FE
0946
08B1
0998
0ACF
0933
032D
FAF9
F4F0
F390
F592
F7AD
F7D4
F68C
F57B
F567
F5DC
F632
F64E
F65C
F66F
F69D
F710
F7B1
F7FD
F79C
F701
F70C
F7EA
F8BD
F8C7
F87B
F8CB
F994
F9A7
F88C
F76B
F797
F8CD
F9A1
F957
F892
F83F
F879
F8D6
F91B
F938
F8F1
F83E
F7D2
F860
F94C
F914
F773
F612
F671
F7D2
F84C
F773
F6BA
F723
F7D5
F79D
F6ED
F721
F80C
F7DF
F60F
F526
F858
FFA0
075E
0BCC
0C39
0ACF
0A01
0A83
0B57
0B4A
0A36
0919
0906
0A10
0B37
0B7F
0B05
0ACE
0B84
0CD4
0E18
0F1D
0FF4
1071
105E
0FED
0F8C
0F5D
0F3C
0F26
0F49
0F8B
0F79
0EE1
0E49
0E6D
0F4A
1009
1002
0F6F
0EEE
0EBB
0EA8
0E8A
0E60
0E38
0E40
0EA9
0F4E
0FA7
0F60
0EC3
0E27
0D2D
0B23
0870
06D6
078D
097E
0A5D
099F
091B
0A06
0A75
0732
FFF2
F862
F47E
F4A6
F5FD
F60A
F4FF
F46E
F4ED
F5CF
F670
F6D3
F705
F6CB
F63A
F609
F6C4
F7EE
F86D
F7D8
F6F0
F6A6
F707
F75E
F744
F718
F750
F7D7
F84C
F8AD
F941
F9F4
FA24
F96D
F84C
F7B4
F804
F8A9
F8E8
F8AB
F868
F86D
F895
F8A8
F8A0
F890
F886
F8AD
F923
F99E
F984
F8BC
F80F
F840
F8F7
F916
F83F
F76A
F785
F7F9
F791
F6C2
F7FC
FCFA
0450
0A6E
0CF9
0C8F
0B65
0AEF
0B27
0B72
0B78
0B3B
0AEC
0AED
0B7B
0C2E
0C1F
0AF7
097E
08C7
0904
0997
0A18
0AAB
0B5B
0BA7
0B25
0A48
0A15
0B07
0C91
0DDD
0EBF
0F97
1082
1111
10D3
0FE0
0ED2
0E41
0E55
0EB8
0EEA
0EBB
0E59
0E06
0DD4
0DC0
0DD0
0DFF
0E28
0E24
0E0D
0E20
0E4B
0E1D
0D70
0CE7
0D4D
0E66
0F00
0E77
0D96
0D75
0DE0
0D82
0BB7
0985
087F
08F5
09C2
09C9
091C
088B
088F
08EA
091D
08DE
0847
07CA
07D5
084F
08B3
08C4
08DD
094A
099F
092F
0823
077B
07CE
0883
08D2
0903
09A7
09C3
0710
00D7
F9A7
F51B
F442
F529
F5BE
F60C
F70A
F872
F8E4
F80C
F73B
F783
F834
F805
F71C
F6CB
F792
F864
F82B
F743
F6E6
F780
F848
F864
F7F9
F7C9
F829
F8B6
F8DF
F87B
F7D2
F763
F788
F817
F869
F7FA
F70B
F66F
F6AA
F76D
F7FD
F80B
F7EA
F809
F855
F85A
F7DB
F71C
F691
F663
F668
F675
F68A
F6BA
F6FC
F72C
F73A
F738
F72C
F6FD
F6A1
F65E
F687
F707
F771
F781
F75F
F740
F71B
F6E0
F6C0
F6E8
F71D
F6F5
F68C
F68B
F740
F800
F7F4
F74E
F71A
F7C3
F888
F8A1
F84E
F834
F85F
F886
F8E5
F9CF
FA88
F9B0
F7A8
F79B
FC96
0597
0DC4
113A
10B3
0FAF
1009
10AA
1038
0F46
0F2E
0FDB
0FF4
0EF6
0E08
0E55
0F6A
0FEE
0F77
0EED
0F25
0FCA
0FD2
0EA1
0C97
0ABA
09DB
09F0
0A33
09FA
096D
0945
09CB
0A67
0A46
0973
08D7
0926
0A07
0A8E
0A5B
09E2
09BD
09FD
0A3C
0A21
09B5
094B
0921
0927
0927
0911
090B
092A
0951
0959
0932
08D5
0856
0819
08BB
0A7F
0CAF
0DFD
0DCA
0CE3
0C89
0CEF
0D2E
0CC2
0C52
0C9F
0D5A
0DA5
0D59
0D1D
0D50
0D83
0D3E
0CB8
0C7F
0CA6
0CD7
0CF9
0D25
0D1C
0C98
0C30
0CD8
0E2A
0E5B
0CC7
0B74
0C92
0EBD
0D7E
0666
FC8B
F5B1
F453
F5E4
F6CE
F671
F64E
F6D3
F6D6
F5C9
F4C6
F4EB
F5CD
F633
F5C5
F54F
F57E
F612
F663
F632
F5AF
F529
F506
F597
F693
F705
F65F
F53F
F4BC
F516
F5A1
F5DA
F604
F684
F728
F75C
F6FD
F688
F674
F6B1
F6F4
F72C
F76C
F79E
F7A2
F79A
F7D0
F841
F890
F856
F786
F68D
F61F
F6A3
F7B3
F86C
F85B
F7EF
F7D9
F819
F819
F7A4
F75D
F7E4
F8D2
F922
F897
F819
F86A
F913
F91F
F871
F7DC
F7FA
F876
F88B
F7EE
F715
F6AF
F6F7
F77A
F79D
F75E
F763
F821
F8F4
F89F
F70A
F5E8
F6BC
F86A
F842
F5E0
F4C0
F8A7
00EF
08D1
0C4D
0BC5
0A4F
09BF
098B
090C
08F9
0A0A
0B5D
0B77
0A4F
0946
0938
09A4
09D5
0A07
0AF6
0CB1
0E62
0F35
0F12
0E77
0DF2
0DE0
0E57
0F08
0F61
0F18
0E7D
0E0C
0DE3
0DCD
0DB7
0DC1
0DFB
0E51
0EA1
0EC1
0E96
0E3A
0E04
0E27
0E6E
0E73
0E25
0DE7
0E13
0E85
0EDF
0F0F
0F31
0F09
0E1B
0C80
0B03
0A2D
09A4
08E8
083F
084E
0902
097D
0934
0898
0876
08EC
096C
098D
0974
094C
08FB
087A
0810
07E8
07D7
07CA
0803
0895
090F
090B
08B0
0840
07AC
0705
0710
086A
0A1B
0A16
0801
068D
086A
0BFF
0C19
05CA
FC4E
F5BD
F4A0
F64F
F731
F6BC
F695
F746
F790
F6AC
F5A2
F5B9
F6A6
F731
F6FA
F6B4
F6DD
F72F
F74C
F73D
F734
F73C
F758
F785
F792
F73A
F69C
F655
F6CA
F782
F79F
F713
F6C5
F753
F826
F83C
F77D
F6B7
F685
F6C1
F700
F728
F74E
F76B
F758
F715
F6DD
F6DD
F6EE
F6C5
F653
F5E6
F5DD
F645
F6CC
F710
F708
F70C
F751
F781
F731
F6A1
F695
F739
F7CB
F797
F6E1
F66A
F669
F681
F695
F710
F81D
F921
F961
F8F8
F8A0
F8A9
F8C9
F8E8
F94A
F9CB
F9BF
F911
F8AA
F91E
F9AC
F967
F8E2
F964
FA86
FA26
F7BA
F68A
FABA
0400
0D02
10DE
1001
0E85
0EDC
0FDB
0F9B
0E5F
0DCF
0E6A
0F06
0E90
0D48
0C0E
0B35
0A92
0A1F
09F2
09E2
09BC
099A
09A0
099A
0954
0920
0980
0A56
0AF4
0AEE
0A89
0A37
09F2
0983
0921
094D
09FE
0A6E
0A13
0964
092F
097C
0994
090A
084F
081C
089B
094A
0996
098D
09DD
0B13
0CD5
0E1F
0E4A
0DAC
0D21
0D14
0D46
0D77
0DD9
0E8F
0F0D
0EA3
0DA7
0D47
0DFA
0EBB
0E68
0D50
0CBD
0D39
0DFA
0E0E
0D7C
0D05
0D0F
0D58
0D7B
0D5E
0D07
0C8A
0C38
0C60
0CCD
0CED
0CA1
0C3B
0B8F
09EB
07A4
06A6
0837
0A67
0929
02BA
FA30
F495
F3CC
F55E
F62B
F5CE
F5BC
F677
F70A
F6CE
F643
F609
F610
F60D
F622
F67C
F6CE
F6B3
F66A
F690
F717
F737
F6A9
F63C
F69C
F73A
F70A
F60D
F54A
F576
F638
F6EA
F763
F7CD
F811
F7F6
F79E
F77F
F7BD
F7E2
F785
F6E7
F6A8
F707
F7B9
F84B
F86C
F809
F76A
F718
F752
F7B3
F79F
F6FA
F64B
F62A
F6AD
F765
F7D7
F7D5
F78C
F74F
F765
F7C9
F81F
F813
F7BC
F779
F75B
F721
F6C5
F6A7
F6E6
F710
F6BB
F626
F5D7
F5EC
F62B
F68C
F736
F7E7
F7F5
F739
F680
F690
F70C
F72C
F740
F839
F986
F918
F687
F51A
F8CF
015C
09B0
0D07
0B9E
097F
0971
0AA0
0B1D
0AE6
0B6B
0D1A
0EDF
0FB8
0FB4
0F5E
0F07
0EDC
0F00
0F41
0F2A
0E9E
0E31
0E6E
0F01
0F0B
0E61
0DDD
0E27
0ECA
0EF1
0E83
0E0F
0DD8
0DAF
0D7D
0D7A
0DC3
0E20
0E52
0E58
0E49
0E2A
0E06
0DFF
0DFF
0D75
0BEE
09E6
088F
0871
08CF
08BA
084D
084D
08DA
0929
08A0
079F
0704
0724
0796
07DF
0802
0845
08A6
08CD
088E
0828
07FF
082E
086D
086B
082C
080B
0838
0866
0849
082B
087D
08E9
0899
07AE
0791
0937
0B9F
0CF2
0CDF
0CE0
0DC1
0E3A
0D04
0B7B
0C25
0E63
0DC9
072E
FD32
F5F1
F486
F66C
F773
F695
F5DC
F69A
F7A3
F762
F61F
F555
F59A
F63F
F697
F696
F661
F610
F5E1
F615
F67F
F6A9
F68A
F695
F704
F755
F6F4
F617
F58A
F593
F5AF
F580
F56D
F5D8
F659
F64A
F5CA
F585
F5A5
F5A4
F52A
F49E
F492
F500
F56C
F59A
F5CA
F627
F66C
F647
F5E5
F5C0
F5F9
F63A
F633
F5F2
F5CE
F609
F691
F704
F71C
F70C
F744
F7CA
F830
F838
F838
F893
F915
F928
F8B5
F858
F89A
F937
F988
F970
F950
F940
F8F4
F884
F87A
F8E3
F900
F86D
F7E8
F840
F8FC
F907
F86D
F863
F93E
F98F
F877
F810
FBC2
03C0
0BD6
0FA8
0F2D
0DC1
0DAF
0E43
0E21
0DB6
0E4D
0FC5
1080
0FA9
0E4B
0DCF
0E33
0E80
0E54
0E24
0E35
0E29
0DBD
0D3A
0D12
0D4F
0DAA
0DE2
0DEF
0DEF
0E03
0E36
0E6E
0E73
0E25
0DAF
0D62
0D56
0D5A
0D48
0D34
0D28
0D08
0CE6
0D11
0D9E
0E0F
0DE1
0D34
0CA6
0C97
0CDD
0D1F
0D39
0D2F
0CFF
0CB3
0C7E
0C8A
0CB1
0CA7
0C7F
0C99
0D07
0D63
0D6D
0D63
0D78
0D68
0CED
0C5E
0C42
0C7C
0C5C
0B9C
0AD9
0ACD
0B63
0BEB
0C1A
0C41
0C87
0C8C
0C13
0B7C
0B3D
0B4E
0B77
0BBF
0C11
0BF5
0B40
0ACD
0BAC
0D5D
0DA0
0AD0
0613
026E
019E
029D
0365
034D
02F6
02C5
0278
020B
020D
02BE
037F
0394
0315
02B6
02CD
0300
02F2
02CE
02DA
02F2
02D3
02A1
02B7
0300
0301
0289
0208
0210
02AA
0352
0385
0351
0330
035D
037C
0333
02F8
03F3
06B9
0A51
0CD9
0D4E
0C74
0BC2
0BB8
0BC2
0B8A
0B87
0BFF
0C40
0B93
0A74
0A22
0AF0
0BCF
0BBE
0B1C
0B11
0BE8
0CAC
0C7E
0BA7
0B06
0AEE
0B0A
0B0B
0AEE
0AB7
0A62
0A18
0A1C
0A6C
0AB5
0AD5
0B15
0BA9
0C0F
0B43
08C4
0544
0237
00AF
00B9
0181
01FC
019F
00C2
003E
0085
0130
0188
014F
00E1
00B0
00D7
011E
013B
0108
00A5
0063
0081
00D2
00D4
0058
FFE8
0029
00F0
0168
0135
00E7
0104
0132
00D1
001B
FFDF
0037
004D
FFCC
FFF0
023B
063A
0981
0A45
0949
08B5
0970
0A78
0A9F
0A0C
09AA
09CE
09FE
09E2
09C6
09FC
0A39
09FB
0959
08FE
0946
09C4
09D8
0974
0915
0915
093F
0931
08EC
08D7
092F
09A2
09B4
0959
08F5
08D7
0902
096A
09FC
0A33
0909
05F2
01E6
FEEB
FE42
FF35
000D
FFFF
FFA5
FFAE
FFE3
FFCD
FFA8
0005
00C9
0131
00EB
0085
007E
007E
FFF8
FF37
FF16
FFA6
FFE6
FF3A
FE74
FEBF
FFEB
009F
0031
FF87
FFBC
0099
00FB
007D
FFF6
0017
0057
FFE2
FF48
0042
0399
07CB
0A59
0A4A
08F6
0851
08E3
09AB
09B0
092A
08E0
08FD
0903
08BC
08A2
091E
09CE
09FA
098C
0920
0928
0957
092F
08CC
08B1
08F4
0916
08C8
085C
083B
084B
0835
07FF
07F0
0812
0835
0881
0959
0A67
0A42
07B5
0370
FFC1
FE62
FEE5
FF93
FF73
FEE1
FE84
FE6E
FE70
FEA6
FF3A
FFCD
FFB9
FEF1
FE3C
FE42
FEC1
FEF4
FEB1
FE94
FF0A
FFA2
FFA3
FF0A
FE8E
FEAD
FF07
FEEF
FE61
FE10
FE71
FF23
FF7C
FF69
FF4C
FF30
FEBA
FE23
FEA9
0150
0549
0844
08B2
0763
0679
06FD
080E
0862
07DF
0752
0728
071E
06FF
0707
075D
07A9
0794
075C
078A
081C
0873
0827
0798
076D
07C5
083D
0887
08A4
0892
083D
07C3
077D
0783
0772
06F2
066B
06B0
07CC
086B
06FF
0388
FFDB
FDF1
FE17
FEE9
FF06
FE59
FDC2
FDC1
FDF6
FDDA
FD82
FD5C
FD75
FD69
FD11
FCD0
FCF6
FD42
FD42
FD08
FD0E
FD7B
FDE0
FDE0
FDBC
FDF3
FE76
FEB5
FE74
FE19
FE02
FE03
FDE0
FDE2
FE64
FEFE
FEC6
FDAF
FD24
FEB8
0249
05F2
07E3
0808
079A
077C
0784
073D
06CD
06BD
0731
07B5
07D1
0793
075F
0768
0788
0795
07A4
07CC
07DE
0799
070F
06A4
0692
06AA
06A7
0694
06AD
06F0
0715
0704
0700
0724
0706
064F
058C
05B6
06A3
0697
0400
FF95
FBF7
FB14
FC48
FD65
FD2E
FC49
FBE1
FC23
FC64
FC50
FC35
FC54
FC70
FC41
FBEF
FBDE
FC22
FC6C
FC7E
FC69
FC55
FC42
FC26
FC28
FC81
FD23
FDAD
FDD7
FDB7
FD88
FD54
FD15
FD01
FD69
FE21
FE50
FD5C
FC1C
FC91
FFE1
04A8
07F3
0820
066A
055B
05FC
0725
0759
06A6
063E
06B4
075B
076A
0708
06DA
06FE
06FB
0691
0618
05FF
0643
0690
06AD
0695
065D
062A
0639
06A7
0722
0725
0699
0608
05F0
0623
062E
0625
068C
074C
0730
04F7
00EF
FD17
FB58
FBBB
FC9E
FC9A
FBDD
FB89
FC15
FCD1
FCE9
FC78
FC3A
FC7C
FCB5
FC5B
FBB3
FB7A
FBEB
FC7A
FC91
FC45
FC17
FC4F
FCC3
FD2D
FD6E
FD84
FD7E
FD80
FD99
FD93
FD1A
FC51
FBF2
FC7B
FD51
FD4A
FC55
FC0C
FE18
021F
05DA
0758
06CB
05E2
05CC
0648
0690
067E
0675
0696
0694
0648
05FB
05FD
0635
0654
064D
0657
0688
069D
0657
05D2
0568
0542
0539
052D
0538
0576
05BC
05C3
058F
0573
0596
05B3
057D
052A
0531
055B
0488
01D3
FDFD
FB1C
FAA2
FBE0
FCDD
FC71
FB40
FA98
FADA
FB50
FB53
FB06
FAE4
FB07
FB2C
FB32
FB39
FB51
FB62
FB5D
FB60
FB81
FBB1
FBE3
FC2C
FC84
FC9F
FC3A
FBA2
FB81
FC01
FC7C
FC4A
FBC0
FBC6
FC88
FD07
FC73
FB9B
FC68
FFA7
03C6
0642
062C
04E9
0462
04EE
056E
051E
0495
04DD
05F5
06CC
06A1
05DC
0569
0588
05B4
0584
0535
0537
0586
05C3
05B1
056A
0519
04D9
04CB
050E
0574
0595
054C
0504
0529
057B
055A
04D2
04BD
0579
05E6
0463
00CC
FCF8
FAED
FAE9
FB95
FBD6
FBCA
FBFC
FC51
FC49
FBED
FBCB
FC0E
FC25
FB97
FAC8
FA8E
FB1C
FBCF
FC07
FBDA
FBB9
FBBA
FB99
FB47
FB0E
FB1A
FB37
FB37
FB52
FBCD
FC64
FC83
FC1D
FBE2
FC4A
FCB8
FC2C
FADB
FA86
FCB0
00C1
0461
05CC
0565
04C6
04CE
050D
04E7
0495
04B4
0543
05A2
0572
0512
050A
0568
05D7
0622
063F
0617
0594
04FC
04CF
0524
056C
0523
048D
046E
04FE
059E
05AD
055A
0535
0540
04EF
0431
03D8
0488
0576
04DB
01E3
FDCB
FAC4
F9DB
FA48
FAB7
FABA
FABB
FAFC
FB24
FAE2
FA84
FA92
FB09
FB58
FB27
FACA
FABC
FAEB
FADA
FA5D
F9EB
FA03
FA8F
FB0C
FB31
FB2A
FB3B
FB64
FB88
FBA2
FBAC
FB75
FAE0
FA44
FA34
FAB3
FB05
FAA4
FA42
FB5D
FE8C
028D
0555
0603
0577
0503
0504
04FD
04B9
04AF
0538
05DB
05D0
0505
043B
041E
0488
04E2
04F2
04FB
052C
0550
0535
050D
0527
056F
057D
052D
04D1
04B6
04B7
0485
0434
041D
044A
045A
0424
0410
0468
047D
0315
FFDF
FC38
F9F7
F9A8
FA46
FAA0
FA96
FAA9
FAE3
FAB5
F9FA
F96D
F9CB
FACA
FB67
FB1F
FA79
FA37
FA66
FA88
FA75
FA7E
FACA
FAF4
FA9F
FA17
F9FD
FA60
FA9E
FA43
F9A6
F970
F9BB
FA11
FA25
FA29
FA50
FA74
FA98
FB63
FD89
00AA
034C
0448
03FB
03AE
03FF
045F
0425
0399
0386
0411
0492
048B
0442
0439
046B
0475
0445
043E
0487
04BD
0488
0436
0450
04CF
0510
04C0
0452
045C
04C1
04E9
04A7
0477
04AB
04E2
049C
041B
0406
042E
034C
0073
FC87
F9A5
F906
F9DD
FA8A
FA6A
FA26
FA5D
FACA
FACC
FA64
FA24
FA58
FAB5
FAE8
FB03
FB29
FB30
FADA
FA50
F9F9
F9F5
FA06
FA15
FA5A
FADF
FB21
FAA4
F9B7
F937
F970
F9B6
F95B
F8A7
F868
F8C9
F929
F921
F921
F9A4
FA48
FA50
FA0F
FAF9
FDF2
01DB
0481
04D8
03EF
0380
0414
04D5
04E7
0460
03F0
03EF
0424
0434
0404
03AB
034D
0314
031A
0346
0350
0325
030B
0346
03AD
03C9
0379
0327
0338
0384
039F
0381
0395
03FA
0430
03C1
030B
02E1
036A
03E6
03BF
035A
0351
033E
01EC
FF01
FBCC
F9FB
F9BF
F9DA
F95F
F8BF
F8D3
F974
F9B5
F937
F89C
F894
F8F9
F935
F925
F926
F968
F9A7
F9B1
F9B7
F9E9
FA0E
F9DF
F98D
F983
F9BF
F9CF
F990
F96F
F9C7
FA3C
FA29
F98D
F91D
F947
F9A4
F9AB
F988
F9BC
FA28
FA1A
F993
F9DC
FC44
004F
03DB
0538
04CC
0446
0488
04F7
04C3
0430
0425
04C0
051C
048D
038E
0326
039B
0434
0434
03AE
033C
033A
038F
03FF
045D
0473
041F
039F
0372
03C4
042C
0438
0400
03F1
0420
043C
0429
0438
0490
04C0
0461
03ED
0434
04E4
0450
0151
FD00
F9E4
F952
FA36
FAA4
FA0E
F973
F9AC
FA54
FA88
FA21
F9BB
F9C0
F9FB
FA19
FA1E
FA30
FA4B
FA59
FA6C
FAA1
FAD0
FAAB
FA2D
F9B8
F998
F9AC
F9A5
F986
F98B
F9AD
F999
F933
F8E8
F924
F9AD
F9E9
F9B4
F99A
F9F5
FA45
F9E5
F958
FA34
FD52
0169
0411
0439
0318
0287
02FF
038E
0383
034A
038E
0429
0467
041B
03CF
03DE
03F5
03BC
0373
038A
03DD
03DF
037F
0349
039A
0415
042A
03EA
03D3
03FE
03FC
03A6
0377
03D4
0452
0445
03BE
0372
03A8
03D2
0384
0344
03B9
044A
0350
0011
FC00
F974
F947
FA34
FA93
FA15
F98F
F986
F99A
F958
F8FB
F90F
F98F
F9EA
F9CA
F97C
F976
F9B9
F9F3
FA03
FA0D
FA16
F9EF
F997
F965
F99E
FA0B
FA40
FA32
FA31
FA59
FA53
F9EE
F997
F9D6
FA78
FABC
FA62
FA03
FA13
FA22
F9A3
F944
FA91
FDFC
01D6
03E1
03B9
02FE
032E
0401
044C
03D2
0373
03C4
0449
0444
03BF
0351
0334
031A
02D7
02AE
02C8
02DE
02AD
0278
02A3
0303
0313
02C7
02B3
0329
03A2
036F
02BC
025B
02A1
02F6
02C2
0258
026C
02EA
0319
02CF
02D5
0398
03F4
022D
FE38
FA41
F882
F8F4
F9B3
F976
F8D4
F8F1
F9B2
F9F7
F94B
F891
F8BF
F999
FA24
FA00
F9B1
F9B2
F9DA
F9DC
F9DE
FA24
FA7F
FA82
FA39
FA2D
FA80
FAA0
FA18
F957
F920
F97C
F9C1
F9A0
F98E
F9E9
FA40
F9F8
F95F
F94C
F9CC
F9EA
F94F
F955
FB9F
FFC8
035B
046E
0396
02DB
032B
03A4
034D
028F
027C
0334
03C1
0377
02BF
0255
0251
024E
023B
0270
0306
0388
0386
0321
02C6
029B
027D
0269
0281
02AC
0290
0226
01FA
0274
032A
0350
02D1
0284
02F9
03A6
03A9
031B
02D9
02FC
0235
FF61
FB50
F844
F784
F81E
F85E
F7EA
F7B8
F85B
F920
F928
F8AB
F890
F90E
F97B
F961
F92A
F960
F9C2
F9B0
F924
F8C7
F8F6
F951
F960
F93F
F94D
F974
F94F
F8E9
F8CD
F931
F98E
F96C
F928
F96C
FA16
FA47
F9A5
F8F4
F906
F987
F98A
F927
F9C3
FC54
FFF0
02A8
03A6
03BA
03EE
042E
03D5
0302
029F
0318
03B6
0393
02C9
022F
0231
026A
0272
0279
02CE
0339
0337
02CC
0292
02DE
0345
0339
02D2
02A1
02D9
0315
0307
02E6
0303
033D
033A
0308
0307
033A
032D
02C5
029E
0320
0372
0212
FEAC
FAD6
F88A
F828
F876
F865
F82D
F87B
F92B
F980
F945
F91C
F97C
FA02
FA15
F9C8
F9B5
FA02
FA26
F9C0
F92E
F909
F94F
F988
F98D
F9AF
FA19
FA6E
FA52
F9F1
F9C0
F9C6
F9A2
F937
F8EA
F902
F931
F91A
F8F9
F945
F9BD
F988
F895
F85C
FA84
FEC4
02CF
048F
042A
035E
0354
03AB
0394
031D
02EE
032B
0349
02F9
02A4
02C2
0322
0340
0315
0315
0365
039C
0360
02F9
02E5
0317
0310
02A7
0241
0230
0237
020F
01F5
0253
02F1
031F
02BA
027C
02FE
03B5
03A2
02CD
0254
02B6
02B9
00BE
FCF9
F990
F850
F8DC
F97E
F94D
F8DF
F8F9
F95E
F955
F8DC
F8A1
F8FC
F97E
F9A7
F989
F979
F96C
F91D
F8A5
F87B
F8BD
F8F1
F8B7
F869
F89E
F94E
F9D4
F9D7
F9AF
F9C4
F9E1
F99E
F930
F93C
F9D3
FA34
F9D3
F92D
F918
F97A
F974
F8F1
F94E
FBD2
FFD1
0305
03EC
033C
02B6
0309
037B
0358
02FA
0317
03A3
03EE
03A8
033F
0328
0340
0330
030A
0324
037B
03AC
0390
0370
0387
0393
033B
02AB
0271
02B5
0302
02F0
02AF
02A6
02CE
02CF
0299
027E
0296
0285
022F
0232
0315
040B
034A
0008
FBBC
F8DE
F86B
F928
F95F
F8C7
F85C
F8B7
F94E
F95B
F8ED
F8A6
F8C8
F8FC
F8F9
F8E9
F901
F919
F8E5
F878
F83D
F86B
F8CC
F917
F93F
F954
F951
F933
F92D
F964
F9A0
F984
F91E
F8ED
F934
F98C
F96F
F912
F925
F9B5
F9E8
F93B
F8B1
FA02
FD88
0179
03A1
0393
02C6
02A5
0321
035A
0317
02F9
036C
03FA
03F6
035D
02C7
0299
02B2
02D9
0316
037F
03E5
03FE
03C6
0379
0344
032C
0336
0363
037F
033B
02AD
026F
02EE
03BA
03E5
0335
0284
02A1
0338
034C
02B5
0260
02D9
0317
0177
FDDE
FA35
F877
F8B4
F962
F963
F904
F90B
F970
F984
F90A
F892
F89D
F8F5
F910
F8DC
F8BD
F8E6
F91D
F923
F90C
F90A
F913
F8FD
F8D2
F8C2
F8CD
F8C8
F8B5
F8CE
F914
F926
F8CB
F873
F8C1
F992
FA02
F99B
F911
F95B
FA3A
FA6B
F97F
F8E2
FA6F
FE23
01DF
03A0
036E
02D6
02E0
0337
032E
02E4
02F0
035D
0394
033F
02C6
02B2
02F9
032A
031F
0322
0364
03AC
03B1
037D
0351
033C
031A
02E5
02C7
02D2
02EB
0305
033E
038E
039A
031F
0280
0272
0303
035F
02E1
0219
0223
02F1
02E2
0086
FC8E
F956
F878
F94A
F9F6
F9A7
F90B
F900
F962
F983
F937
F8FA
F916
F93A
F90D
F8BB
F8AF
F8F1
F922
F910
F8F3
F908
F941
F969
F97A
F98F
F9A0
F986
F950
F93F
F963
F97B
F957
F926
F92C
F94B
F935
F902
F924
F9A7
F9D5
F931
F892
F9A4
FCFC
0106
036C
0373
0283
0251
030D
039D
0352
02B7
02A3
0318
0367
033B
02F5
02FF
033A
0345
0312
02EE
0302
0322
0321
0311
0315
031A
02FA
02C1
02A4
02B1
02C0
02BB
02C9
0306
033E
0328
02D9
02A8
02BA
02D1
02C5
02D3
0332
0389
0345
0286
0231
02C0
0332
01E3
FE83
FAC7
F8C3
F8D2
F987
F98D
F901
F8CE
F93B
F9A3
F982
F926
F925
F97C
F9A7
F960
F8F0
F8B8
F8C0
F8DD
F902
F93E
F975
F973
F943
F92C
F952
F97E
F972
F942
F92A
F930
F922
F903
F913
F96D
F9BF
F9B1
F960
F935
F946
F93D
F8F6
F8DA
F941
F9B9
F973
F899
F8A6
FAF5
FF04
02A5
040E
037E
029D
0290
0312
034F
031F
0300
033D
0386
037A
0330
0307
031C
033D
0348
0353
0368
0361
031B
02C1
029D
02B7
02D9
02E6
0300
0342
0380
037D
0347
031D
030F
02F4
02BE
02AA
02DD
031E
0321
0304
0324
0377
036F
02D7
0264
02DA
03B7
0341
0064
FC31
F90C
F853
F932
F9E9
F9B4
F928
F8FE
F922
F91B
F8DB
F8B8
F8D5
F8F1
F8E2
F8DD
F91E
F970
F971
F91C
F8D7
F8E9
F92A
F94C
F94D
F960
F98D
F9A1
F97F
F94F
F944
F958
F96A
F97D
F9A7
F9CA
F9AD
F957
F923
F944
F977
F961
F932
F969
F9FA
FA16
F944
F879
F97A
FCDE
010D
03A8
03DB
02E9
0285
0308
0398
039A
0365
0382
03D2
03D8
0383
0347
0362
037E
033E
02D7
02CC
0332
0392
0386
0339
0315
0331
0348
0329
02F3
02D4
02CE
02CE
02D8
02F6
0312
0311
0302
030D
0327
0321
02FE
030C
0364
0395
032F
028D
02A1
0391
0400
023C
FE47
FA39
F846
F8A1
F99D
F9BB
F914
F8A8
F8DF
F933
F924
F8E9
F8FB
F94F
F96C
F923
F8CC
F8C8
F8FE
F918
F8FF
F8ED
F90A
F938
F94B
F946
F94C
F968
F98B
F9A7
F9B3
F9A7
F985
F96F
F983
F9A6
F995
F94F
F92A
F962
F9A7
F979
F8EF
F8C4
F960
FA10
F9D0
F8D7
F8DD
FB5B
FFA2
0341
0464
0387
0292
02B3
0371
03CF
03A5
0387
03C2
03F2
03B2
0332
02F0
030E
0348
036A
038A
03B7
03C6
0393
0348
032D
0343
0348
0320
02F5
02EF
02FE
0308
031C
034C
0363
0322
02BA
02AF
0328
039F
0391
033B
0341
03A1
039A
02D0
021B
0280
0382
032F
004B
FC08
F8FB
F877
F971
FA07
F99E
F90C
F917
F97C
F987
F920
F8C0
F8B1
F8C2
F8BC
F8C0
F8F9
F942
F957
F93A
F932
F95E
F98D
F98F
F97E
F98D
F9B1
F9B7
F99D
F994
F9AE
F9B5
F98D
F96C
F993
F9D6
F9C7
F955
F8F8
F90D
F950
F943
F8FC
F913
F9A9
F9FE
F97B
F8F3
FA19
FD80
0190
03F5
03FD
030D
02D2
0378
03FE
03CA
0356
0345
0384
0396
0369
035B
0394
03C7
03B2
037E
036D
036C
033C
02EB
02C6
02DE
02EB
02C7
02B8
0303
036D
0386
034A
0327
0350
0378
0356
0327
0355
03BD
03D1
036B
0317
0346
0398
0377
031C
035A
0433
0436
01EB
FDB9
F9DB
F83A
F8A5
F970
F970
F8EE
F8C3
F914
F95C
F946
F910
F911
F93E
F959
F95E
F978
F9AC
F9C8
F9B4
F99B
F99B
F98B
F945
F8F8
F903
F96F
F9DA
F9F7
F9ED
FA04
FA24
F9F0
F963
F8F5
F8FA
F931
F92B
F8F7
F901
F94F
F965
F919
F8FA
F984
FA29
F9EB
F901
F92A
FBD0
0014
0364
0429
0346
02B6
033B
03FE
0419
03BE
039B
03C9
03D2
038F
0361
0386
03B6
0399
0358
0351
0378
0371
0323
02E7
02F7
0316
02FD
02D6
0303
0375
03B0
0371
0313
0309
033F
034F
032B
032F
037D
03B5
0389
0340
0356
03A6
0387
02D9
0276
031A
0401
0350
0023
FBDB
F8EF
F87A
F969
F9FB
F9A7
F92C
F934
F97A
F96D
F911
F8E8
F91E
F954
F93F
F913
F926
F96D
F99B
F99E
F9A6
F9C2
F9C8
F9A3
F98A
F9AB
F9CE
F9A8
F95A
F958
F9BA
FA08
F9E2
F986
F96A
F988
F978
F931
F92B
F99D
FA05
F9E1
F988
F9C1
FA75
FA91
F99E
F8EA
FA5B
FE1A
0211
03FE
03AE
02C3
02A1
032C
0393
039D
03B5
0409
043B
03FE
038F
035D
0379
03A9
03CB
03EC
0400
03D5
0368
030E
030C
0339
0340
0322
0333
0387
03BA
0370
02E3
02A4
02DF
032F
0336
031C
032F
0354
0333
02E0
02E5
036F
03D7
037A
02CA
02E6
03E5
0425
01F0
FDAD
F9CD
F859
F8FD
F9D0
F9AE
F921
F91D
F993
F9BC
F961
F912
F944
F9A8
F9B7
F972
F942
F94C
F950
F92F
F92D
F973
F9B9
F9AD
F974
F978
F9BF
F9E4
F9B4
F980
F99D
F9E1
F9E1
F999
F96F
F990
F9B4
F9A4
F9A7
FA04
FA63
FA2D
F981
F945
F9E9
FA9E
FA57
F972
F9C2
FC7E
009A
03A5
044C
0379
02F5
036B
041D
0439
03E0
03B2
03DB
03F3
03AF
0345
0315
0333
036A
0394
03AF
03B8
03A1
0370
034A
0342
0343
0339
0337
034F
0365
034F
0320
0319
0347
0368
034E
0331
035F
03AD
0398
030A
029D
02D3
034D
0339
0291
0255
0320
03EA
02D5
FF60
FB45
F8DB
F8C1
F99F
F9EB
F975
F909
F91A
F951
F941
F905
F8F8
F927
F95C
F97D
F99C
F9AE
F993
F95D
F953
F994
F9D9
F9D9
F9B3
F9B8
F9E0
F9CC
F969
F92F
F981
FA0E
FA39
F9F1
F9C7
FA09
FA42
F9F1
F962
F954
F9D8
FA1F
F9AE
F931
F98F
FA7C
FAB4
F9D9
F96C
FB3B
FF1B
02D0
045A
03E7
0329
033D
03C9
0400
03CF
03B3
03DB
03F0
03B8
036B
0353
035E
0358
0350
037D
03C4
03C4
0360
02FA
02FA
0341
0360
033E
0334
0372
03A9
037A
030F
02EC
0338
0385
0379
034B
0362
039F
0389
0317
02D4
0319
0370
0340
02D0
0301
03D0
03C3
016B
FD53
F9C8
F88B
F922
F9CB
F999
F923
F93C
F9BA
F9E7
F997
F951
F96C
F9A0
F996
F974
F98C
F9C4
F9C4
F98B
F97D
F9C1
F9F9
F9C6
F958
F931
F976
F9CA
F9E2
F9DF
F9F8
FA16
FA04
F9DC
F9E6
FA21
FA3B
FA10
F9E3
F9F1
FA0B
F9D8
F97C
F976
F9E2
FA24
F9C5
F967
FA69
FD58
010F
03A3
042F
037E
02FB
0342
03D7
0412
03E8
03C0
03CE
03DC
03BE
0393
038D
03A6
03AF
03A0
039F
03B7
03B3
0370
0325
0329
0379
03BA
03B4
0394
0399
03B6
03B1
0383
035A
034C
0343
0342
0374
03D7
03FD
038E
02D5
0288
02DE
035D
039F
03E4
0461
0456
028A
FEE4
FB10
F910
F940
FA34
FA71
F9D7
F93D
F928
F95E
F983
F996
F9B1
F9C1
F9A9
F988
F999
F9D8
FA06
FA04
F9FD
FA24
FA5F
FA69
FA2B
F9D5
F99E
F993
F9A4
F9BB
F9CE
F9D8
F9E2
F9F4
FA0F
FA27
FA2D
FA1E
FA0A
FA15
FA4B
FA87
FA88
FA3B
F9D9
F9B8
F9E3
FA11
FA1A
FA3B
FAAC
FB09
FAA3
F99E
F951
FB0D
FE98
0232
0439
0493
0449
042F
043F
0425
03E6
03B2
038B
035E
034E
038B
03EB
040B
03CF
038A
038B
03BC
03CE
03B3
039F
03B5
03D3
03D2
03C3
03BF
03BC
03A9
0397
039D
03A2
0380
0349
033A
0365
039F
03B7
03B1
03AC
03AF
03A9
0391
0371
0344
0308
02E1
02F4
031E
031D
0306
034B
03E3
03CE
01EC
FE68
FAE7
F911
F914
F9C2
FA05
F9D1
F9A9
F9C3
F9E9
F9F1
F9EA
F9DE
F9C3
F9A6
F9B0
F9EC
FA2F
FA49
FA3C
FA27
FA14
F9F0
F9B9
F991
F99A
F9D0
FA1A
FA61
FA87
FA7B
FA51
FA3A
FA42
FA3C
FA0F
F9E5
F9EB
FA15
FA39
FA53
FA78
FA8F
FA5F
F9F6
F9C3
FA0D
FA84
FAAB
FA99
FAC6
FB19
FAD7
F9E8
F9A3
FB98
FF85
033A
04C8
045B
03A3
03B9
043B
045E
0423
0408
0423
0414
03BF
0381
039B
03D5
03DE
03BA
03A6
03AE
03A6
0383
037D
03BA
040F
0430
040E
03D9
03B8
03AE
03AD
03A7
0395
037C
036C
0370
0382
039A
03B5
03BC
0390
0340
0313
033C
038F
03B1
0397
0399
03D6
03DF
0358
02D3
0344
046C
047E
01FB
FDA4
F9F5
F8A1
F91F
F9C9
F9DB
F9CC
FA09
FA3E
FA04
F9A6
F9B1
FA18
FA5A
FA4C
FA44
FA75
FAA3
FA8D
FA5D
FA63
FA91
FA89
FA2A
F9C0
F9A3
F9CD
FA07
FA3A
FA72
FA9F
FAAA
FA9A
FA8A
FA78
FA58
FA35
FA21
FA19
FA0B
F9FE
FA09
FA2A
FA42
FA42
FA3D
FA3A
FA23
FA06
FA3B
FAE7
FB6E
FAFF
F9F5
F9F9
FC56
0047
0393
04CA
0478
040C
041F
043C
0401
03BA
03C0
03E3
03CC
03A2
03C0
0414
0436
0411
03FA
0421
0441
040C
03AA
0384
03B4
03E9
03E3
03C3
03C2
03D7
03D0
03A8
0384
0380
03A3
03E7
042D
0446
042C
0412
041B
0420
03EB
0395
036E
038E
03B6
03B5
03B3
03D5
03D2
0361
02F6
035A
044D
0435
01CD
FDDC
FAA0
F983
F9EB
FA5E
FA3E
F9FE
FA0E
FA37
FA2D
FA17
FA32
FA50
FA32
F9FE
FA08
FA40
FA4C
FA23
FA19
FA58
FA92
FA78
FA36
FA32
FA6E
FA83
FA3D
F9F0
F9FE
FA4D
FA7E
FA71
FA52
FA43
FA3D
FA33
FA20
F9FC
F9D2
F9CC
FA05
FA56
FA76
FA5C
FA49
FA64
FA75
FA4E
FA36
FA80
FAD1
FA75
F9AE
FA00
FC95
009E
03DE
04F0
0470
03E7
0405
0453
0449
0409
03F3
0405
0405
03F5
03F6
0401
03F8
03EE
0403
0420
041B
040B
0425
0458
044C
03E6
038A
03A1
03FF
041E
03DF
03B1
03E7
0442
0465
0458
0455
0455
042F
03FA
03EA
03F5
03E0
03B4
03C4
0422
046B
044B
0402
03F8
0401
03AA
0332
0367
0430
03FB
016B
FD52
FA1D
F947
F9F7
FA65
F9F7
F97F
F9B0
FA32
FA64
FA50
FA61
FA97
FA93
FA45
FA0C
FA2A
FA74
FA9E
FA86
FA38
F9D9
F99E
F9B6
FA10
FA60
FA6E
FA54
FA4F
FA5E
FA44
F9FD
F9CD
F9DC
F9F8
F9FD
FA0C
FA3B
FA57
FA3A
FA1C
FA3B
FA62
FA37
F9E0
F9EC
FA78
FAE9
FACD
FA9E
FAFC
FB72
FAF4
F9CB
F9F4
FCD7
0135
044B
04D7
0419
03DC
0463
04BF
0486
0449
046D
0484
0425
03BB
03E6
047A
04C0
047F
0425
040F
0418
040C
0402
0420
0448
0442
0419
040C
0426
0430
0416
0410
0439
0458
043B
0410
0418
043F
0451
0448
043B
0423
03F4
03D8
03F3
0418
03F5
039F
0391
03E8
0410
03A1
0347
03F0
050D
0492
015B
FCDF
F9C9
F928
F9C3
FA0C
F9D1
F9C5
FA14
FA40
FA1B
FA17
FA71
FAAF
FA66
F9F0
F9DB
FA16
FA24
F9F7
F9F0
FA33
FA73
FA76
FA68
FA7C
FA8C
FA5E
FA14
FA05
FA2D
FA3D
FA2B
FA51
FAC4
FB07
FAC3
FA55
FA49
FA8F
FAB6
FAA0
FA92
FAA3
FA9C
FA69
FA4C
FA6E
FA85
FA58
FA3D
FA93
FAE5
FA6D
F9A8
FA68
FDB3
0219
0508
0582
04C2
0466
04AD
04DE
04AB
0473
046A
0440
03D5
0397
03D7
0436
0440
0420
0441
0491
04A0
045F
0431
044C
0473
0460
0428
0400
03E5
03B7
0397
03BD
040C
0425
040D
042F
049D
04D0
047A
0411
041D
0467
045E
0404
03E4
0422
0442
03FB
03BC
03F0
0432
03ED
037E
03CC
047A
03B2
0064
FC0F
F95D
F93F
FA4A
FAC5
FA7C
FA3D
FA64
FA8E
FA81
FA80
FAA9
FAA4
FA46
F9FF
FA2B
FA77
FA61
FA11
FA0C
FA61
FA9A
FA86
FA78
FAB5
FB03
FAF8
FA90
FA26
F9F5
F9EF
FA05
FA3E
FA76
FA67
FA20
FA08
FA3D
FA5D
FA35
FA2C
FA96
FB0E
FB02
FA9D
FA90
FAF2
FB11
FA93
FA27
FA7D
FAFA
FA84
F991
FA3B
FDA1
0214
04C7
04E3
03FC
03C2
043D
0483
0449
0412
042A
0449
043E
044A
048E
04AD
0466
0419
0435
047F
0480
0449
0451
04A4
04CC
048C
0443
045B
04B0
04C9
048C
044C
043D
0431
040B
0403
043A
0475
047E
0477
047D
0464
041B
03FE
044F
04AC
0480
03F3
03C1
041F
0452
03E1
038B
0440
0536
043B
0075
FBE7
F968
F996
FAAB
FAF5
FA85
FA4F
FA95
FACE
FAB0
FA83
FA7F
FA66
FA10
F9CC
F9E7
FA2A
FA41
FA42
FA6C
FAA3
FAA5
FA8C
FAA0
FAD3
FAC7
FA6E
FA2D
FA47
FA74
FA4F
F9F8
F9EA
FA39
FA72
FA5B
FA43
FA67
FA7C
FA3D
F9F1
F9F9
FA3B
FA68
FA99
FB10
FB91
FB8B
FB02
FAC1
FB2B
FB71
FAC0
F9FB
FB32
FEFA
0335
0547
04E2
03E8
03D8
046A
04A6
0468
0446
0472
048A
0460
0454
04A2
04E6
04AD
042E
03F5
0420
0458
0466
045E
0454
043F
0429
042E
044B
0461
046C
048D
04C6
04E0
04B5
047C
0488
04BE
04B4
0457
0411
0422
0440
0429
040D
0429
0441
040C
03C7
03E7
0442
042A
0394
0378
0467
052B
03C4
FFEA
FBCD
F9BF
F9DA
FA75
FA73
FA26
FA32
FA7D
FA98
FA89
FAA6
FADA
FAB9
FA42
FA02
FA49
FA9F
FA7B
FA07
F9D8
FA0E
FA4F
FA64
FA79
FAB1
FAE3
FADA
FAA5
FA78
FA6C
FA79
FA98
FAC9
FAEE
FAE1
FAB5
FAAD
FAD6
FAEF
FAD2
FAB2
FABA
FAC8
FABF
FAC5
FAF3
FB02
FAAA
FA41
FA64
FB02
FB35
FA97
FA48
FBF5
FFB4
0383
055F
053E
04A1
0495
04DB
04D5
0485
0454
0463
0479
047F
049B
04D2
04E1
04A5
045C
0450
046E
047F
0480
0493
04A7
048F
0450
0421
041D
042D
043A
0449
0465
047F
0489
0491
04AB
04C4
04B2
047D
0453
0443
0431
0423
0445
0486
0491
0457
043E
0482
04AD
043F
03A0
03DA
04FB
0565
0360
FF4E
FB8A
F9EC
FA0D
FA58
FA20
F9FC
FA5D
FACA
FAAA
FA37
FA18
FA65
FA96
FA59
FA09
FA19
FA6D
FA9F
FA9B
FAA0
FAC2
FAD2
FAC1
FABE
FAE0
FAF9
FADB
FAA0
FA88
FA9A
FAA4
FA8B
FA83
FAB9
FB05
FB0F
FAC5
FA76
FA6D
FA96
FAAF
FAAA
FAC5
FB15
FB3B
FAC5
FA12
FA74
FCF8
00F7
0455
0570
04B2
03DF
0416
04D5
0513
04B9
0487
04D2
050C
04BD
0444
044B
04C2
0507
04D8
049D
04B6
04ED
04DE
0495
046C
0471
045F
0428
041F
0468
04A4
047B
042A
041F
0447
0432
03DC
03D3
0464
050A
0514
0499
044D
046C
046C
03FC
03BC
0452
0505
040F
00AD
FC53
F974
F91F
FA3A
FB06
FAEC
FA91
FA94
FACD
FAC4
FA79
FA52
FA78
FAA4
FA92
FA5D
FA56
FA8D
FAC4
FACD
FABF
FABE
FABD
FA99
FA63
FA53
FA77
FAA2
FAB3
FAC1
FAE1
FAE9
FAAF
FA61
FA5B
FAA1
FAC6
FA84
FA39
FA6C
FB03
FB5D
FB3B
FB18
FB46
FB44
FA93
F9FA
FB31
FEDA
0343
05E1
05E6
04D4
047C
0508
0568
0516
049F
0499
04C1
0487
03FD
03BE
0407
0471
0494
0493
04BE
0502
050A
04CC
049C
04AF
04E0
04FB
0505
050B
04EA
0480
0406
03E8
043C
0496
049E
0484
04AA
04FD
0507
049B
042E
0430
0471
046F
042F
0445
04C8
04A5
0296
FEC5
FB14
F962
F9BE
FA99
FA9F
F9F3
F98E
F9DA
FA5D
FA91
FA92
FAC5
FB25
FB51
FB1D
FAD3
FAB9
FABB
FAA1
FA6F
FA57
FA68
FA89
FAA8
FAC9
FADA
FABD
FA87
FA88
FAD9
FB1C
FAE5
FA5E
FA20
FA64
FAAF
FA90
FA4F
FA7F
FB0F
FB50
FAFB
FAA9
FAF2
FB69
FB37
FA9B
FB29
FDF9
0205
04FD
05A2
04DA
0450
0498
0506
04FD
04B7
04B1
04E5
04F6
04DC
04E4
0522
0545
0510
04B8
0490
0494
0489
046B
0472
04A4
04B2
0472
042F
0444
048E
0496
044A
0422
0473
04DF
04CF
0455
0420
0485
0503
04FB
049C
0491
04EC
04FE
046A
03E6
043C
04D0
03DE
009E
FC8D
FA10
F9F1
FAC7
FAE7
FA35
F9C8
FA20
FA99
FA8D
FA45
FA60
FAC7
FAD2
FA53
F9EE
FA2B
FAB9
FAEF
FAB7
FA90
FAB6
FACB
FA81
FA27
FA39
FAAC
FB09
FB1E
FB27
FB43
FB33
FACC
FA68
FA74
FAC9
FAD4
FA7A
FA4E
FAB9
FB54
FB7E
FB4A
FB44
FB6A
FB0A
FA05
F9B2
FBB3
FFE7
0416
060A
05AA
04A7
0464
04C1
04F2
04CF
04DA
053F
057F
0530
04A5
047D
04C8
04FC
04C5
0473
047E
04D3
04F9
04BA
046A
046C
04B7
04F5
04F7
04D6
04B7
04A1
0499
04AF
04D9
04E6
04B9
047E
0471
0481
0464
0415
03EE
0414
0432
03F6
03C4
0444
052A
04F1
0263
FE42
FADE
F9D1
FA85
FB3A
FB11
FA8F
FA63
FA71
FA4E
FA1D
FA5B
FAFA
FB47
FAE2
FA53
FA54
FAE2
FB56
FB4D
FB00
FAC3
FA99
FA61
FA33
FA3D
FA74
FAA1
FAB8
FAD5
FAEF
FACF
FA7A
FA54
FA9E
FB0E
FB30
FB0E
FB19
FB6B
FB93
FB3E
FACF
FAE5
FB68
FB88
FAE5
FA67
FB82
FE92
0255
0508
05F4
05B8
0556
0536
0520
04E9
04C7
04EE
051C
04E6
0459
0408
0458
04F4
0536
04F2
049D
04A5
04E7
04FD
04DC
04D8
050F
052D
04F1
0491
046F
049D
04DB
04F6
04DE
048C
040B
03A1
03A3
040F
0480
04AD
04BC
04E0
04E0
0470
03F0
042B
0504
0508
02E9
FF2D
FBDC
FA6A
FA6C
FA8B
FA34
F9E5
FA12
FA68
FA64
FA1A
FA03
FA42
FA84
FA8B
FA77
FA7E
FAA1
FABE
FACC
FAD9
FAF3
FB16
FB36
FB3E
FB20
FAEE
FADB
FB0C
FB5B
FB73
FB32
FADC
FAC1
FAD7
FADA
FABD
FAB9
FAEC
FB13
FAD5
FA51
FA2D
FAEA
FC10
FC6A
FB57
F9E3
FA21
FD1B
018D
04EF
05D9
0521
048F
04E2
056F
057A
053B
0541
0581
057D
0521
04E9
051B
055A
052C
04A9
0451
0454
046D
0469
0479
04C7
0514
04F9
047E
0412
040A
0457
04B1
04D6
04A7
0448
041C
0473
0511
0542
04B3
040E
044E
0565
0605
0529
038A
02F3
041A
058F
0519
0207
FDE1
FAE1
F9FB
FA74
FB06
FB17
FAD9
FAA6
FA86
FA57
FA29
FA47
FACD
FB61
FB80
FB18
FA9F
FA89
FAD2
FB26
FB56
FB72
FB71
FB21
FA94
FA59
FAEE
FBEF
FC4B
FB78
FA34
F9C8
FA98
FBC5
FC2E
FB9A
FACA
FA97
FB18
FBA4
FB8D
FAD1
FA23
FA34
FAE6
FB62
FB29
FB08
FC66
FF94
031C
0528
0556
04D3
04BB
04F8
04DA
044E
03F7
043B
04BA
04EF
04DE
04D9
04E5
04CD
04A0
04B6
051A
055B
0510
0467
03F8
0416
0477
0495
0445
03DF
03D8
0454
04FE
054C
04F8
0450
03F7
043B
04C3
04FE
04C7
047D
0474
0495
0485
0432
0404
0467
0514
04F8
0314
FF9F
FC26
FA56
FA7F
FB6B
FBB7
FB2C
FA95
FA87
FAC6
FAE3
FAE4
FAFE
FB0A
FABE
FA4D
FA54
FAFD
FB9F
FB8B
FAF2
FAB0
FB29
FBD6
FC0A
FBC8
FB85
FB6F
FB49
FAFD
FACF
FAF6
FB43
FB5E
FB3E
FB2B
FB5C
FBB7
FBF6
FBEC
FB97
FB14
FAA6
FA9F
FB09
FB6C
FB41
FAC0
FB09
FD2A
00E9
049F
068D
0654
0513
0422
03F1
0429
0486
0511
0599
0597
04E2
043A
0484
0595
0634
058F
0450
03D9
0494
0580
0586
04B7
0400
03F1
0451
04B0
04E9
0502
04E8
048F
042F
041A
0463
04C6
04FD
04F7
04C0
046B
0421
0416
0446
046E
0477
04AB
0528
054B
0408
0116
FD8F
FB0A
FA29
FA44
FA7C
FAAE
FB31
FBE1
FC0C
FB59
FA71
FA51
FB19
FBD6
FB9C
FA9B
F9ED
FA4A
FB33
FB98
FB16
FA5F
FA53
FAFA
FB98
FBA1
FB56
FB57
FBC5
FC11
FBA9
FAAE
F9DE
F9DB
FA9B
FB85
FC02
FBE8
FB7C
FB1F
FB0E
FB53
FBCF
FC2F
FC03
FB25
FA38
FA77
FCB1
0052
03A0
052F
051A
04A0
04B1
0514
0516
049A
0430
043E
0484
049A
0495
04D1
053D
053C
047A
0387
0361
044B
0570
05B0
04CE
03A5
0346
03FA
051A
05BC
0581
04C8
043B
0439
049B
04ED
04DF
0481
042F
0434
0488
04DD
04EC
04AD
0456
042A
044B
04A4
04DD
045F
02A8
FFD4
FCCF
FAC8
FA3D
FAAA
FB2B
FB4C
FB20
FAD6
FA88
FA6B
FAD2
FBAF
FC53
FC0B
FB08
FA56
FAAE
FB9C
FC0B
FB83
FA91
FA0D
FA43
FADC
FB5D
FB8A
FB73
FB47
FB30
FB38
FB44
FB43
FB4C
FB76
FB93
FB5A
FAEA
FACD
FB4C
FBF8
FC20
FB9F
FAF3
FA8E
FA72
FA82
FAF8
FC42
FE73
010E
0372
0536
0625
0632
059B
04EE
0498
049F
04D5
0521
055B
0529
0461
0385
036F
0459
0571
05BE
053B
04C4
04E6
0548
055C
0534
0532
0540
04DB
0400
0374
03E3
04F3
058F
0521
0434
03C8
042A
04C3
04F1
04C6
04D4
053D
0548
03EF
0103
FD97
FB2F
FA6F
FAB3
FAF7
FAE2
FAD1
FB11
FB5E
FB48
FAD7
FA8E
FACC
FB58
FB9D
FB4E
FAAE
FA40
FA48
FAAF
FB35
FBA5
FBDD
FBC0
FB4A
FAC0
FA98
FB08
FBB8
FC06
FBB9
FB47
FB45
FBAB
FBE4
FB9D
FB35
FB42
FBAC
FBB5
FAF6
FA31
FAC2
FD3A
00AB
0378
04CD
0529
057E
0611
0653
05C7
04C9
0443
04B8
05BB
0666
063C
0586
04EA
04CF
0520
0581
05A0
0559
04BC
040D
03B8
0411
04EC
0592
0552
044E
037F
03BC
04CA
0596
0572
04CB
047D
04A8
04AB
0447
042D
04FD
0613
05FA
0413
0162
FF5F
FE49
FD2D
FB68
F9AA
F923
FA0A
FB51
FBC5
FB26
FA1E
F97E
F99D
FA49
FB02
FB43
FAE2
FA3D
F9F0
FA4C
FB12
FBC1
FC11
FC04
FBAF
FB2D
FACA
FAED
FB9A
FC3D
FC3A
FBB6
FB6D
FBB2
FC0E
FBF6
FBA6
FBBC
FC25
FC0B
FB17
FA44
FAE0
FCED
FF27
00BB
0235
0455
068A
075D
0651
04A0
03E7
0480
0579
05DE
0596
0515
04BE
04C4
052F
05C3
060E
05ED
05B3
059F
056C
04CC
041D
041C
04E2
05A1
0592
04DD
044D
0443
0476
04A4
04FC
058F
05D6
054E
045D
040A
04BB
05A7
05AF
0486
02C8
0112
FF5D
FD5B
FB44
F9DF
F9BE
FA86
FB3F
FB43
FAC5
FA73
FAA6
FB17
FB53
FB54
FB70
FBC6
FC02
FBCC
FB46
FAED
FB17
FBA7
FC32
FC4F
FBE9
FB54
FB0B
FB3D
FBA0
FBCD
FBAC
FB7B
FB6C
FB68
FB5E
FB80
FBF7
FC60
FC0E
FAFB
FA1C
FA7C
FC17
FDFE
FF88
00FE
02F5
0536
06B5
06A8
0570
044F
0428
04C8
0566
059F
05A6
05B0
058A
04F8
0452
044D
050A
05B7
056F
046B
03C7
0422
04E2
0520
04CA
0483
049A
04B0
0471
0426
0455
0504
059E
0596
04F5
043D
0406
0499
05A3
063E
059F
03EF
021C
00A2
FF03
FCBE
FA80
F99F
FA73
FBC9
FC31
FB83
FAB7
FA82
FAAA
FAC4
FAE9
FB5C
FBE3
FC00
FBA7
FB48
FB34
FB55
FB76
FB87
FB90
FB91
FB89
FB7E
FB64
FB30
FB0D
FB52
FBF3
FC3B
FB82
FA43
F9E1
FAFA
FC67
FC81
FB26
F9DD
F9F2
FB0D
FC18
FCFB
FEBD
01CD
04EC
065E
05E1
04E7
04D1
0586
05FC
05B8
0543
053F
0587
0584
0515
04BA
04E3
0560
05AF
05A1
056B
053B
0501
04A8
0457
044C
0484
04B8
04A7
044B
03E5
03D8
0459
051E
0571
04D8
03C5
035B
0437
05A3
0645
05A4
0487
03B5
02BA
0097
FD69
FAC8
FA25
FB21
FC08
FBCA
FB06
FAE8
FB86
FBE0
FB55
FA82
FA6E
FB32
FBE1
FBBE
FB12
FABC
FB16
FBA8
FBE5
FBD0
FBB8
FB9A
FB27
FA70
FA26
FAD6
FC0A
FC94
FBDD
FAB1
FA69
FB5E
FC81
FCA0
FBC4
FB04
FB25
FBC3
FBFD
FBBD
FBF5
FDA2
00A4
03B7
0582
05A9
04F6
048F
04E9
0584
05A3
0539
04EF
0531
0598
0577
04CC
044B
0475
04FB
0549
054B
054C
0543
04DB
0443
0442
0517
05CD
054D
03F0
034B
0443
05DE
0663
0569
0429
03E9
049E
0554
0575
053A
0523
055B
057A
04A0
022A
FE93
FB7F
FA4F
FAB4
FB18
FA85
F9BC
F9FC
FB2B
FBE9
FB76
FAAA
FAA6
FB4A
FB9D
FB47
FAE1
FAD6
FAD9
FAA3
FA9F
FB45
FC1F
FC25
FB22
FA2F
FA63
FB76
FC29
FBD1
FAFE
FA94
FAC3
FB13
FB23
FB01
FAEF
FB0B
FB44
FB6A
FB51
FB07
FB14
FC42
FEDA
020A
046C
0551
054E
055C
05A1
0580
04CD
0453
04E2
0617
06A6
05EC
04B5
0447
04DD
059D
05C3
056C
050E
04D2
04B0
04CB
0534
0599
0591
0538
0516
0558
0596
0574
0535
0544
0575
053A
0495
0431
0462
04A9
0496
0486
04E7
0511
03BD
00BB
FD7F
FB9A
FB0F
FAC2
FA3D
FA37
FB21
FC16
FBD8
FA8C
F9AD
FA3C
FB95
FC47
FBB9
FAA5
FA26
FA9D
FB8A
FC2E
FC2D
FBB7
FB4C
FB55
FBC7
FC26
FBFA
FB56
FAC4
FAB4
FB14
FB78
FB8F
FB5F
FB27
FB1F
FB55
FBAB
FBDB
FBA3
FB14
FAD0
FBB0
FDF4
00D1
0309
041A
049E
055B
0632
064F
0576
04A0
04ED
0622
06D6
0634
050E
04CD
059C
0648
05EA
0508
04B6
0504
0510
0483
042E
04BF
0595
0582
0486
03FA
04C7
0619
066B
057F
04A9
04FE
05F7
062F
052F
03F0
03B4
04BF
060E
0627
043E
00EB
FDBF
FBFA
FB78
FB1E
FA59
F9D0
FA58
FB85
FBFE
FB3E
FA4C
FA5D
FB42
FBDA
FBA2
FB27
FAEF
FABF
FA43
F9DD
FA44
FB50
FBE8
FB4C
FA31
FA04
FB44
FCDE
FD4D
FC1F
FA6F
F9D7
FAD9
FC47
FC76
FB1F
F9C5
F9F8
FB78
FC6F
FB9B
F9D2
F935
FAF2
FE3A
0151
0354
04A0
05C0
068B
067C
05AA
04F9
0538
0630
06D3
0675
0594
0530
0587
05FD
061C
0613
060D
05C0
0512
04B0
0541
0643
0663
0543
0428
046B
059E
061D
0553
0475
04AE
0599
0613
05D5
0569
0511
04A8
0468
04D1
059D
058C
03BE
00D2
FE30
FC67
FAFD
F9CD
F992
FAAC
FC15
FC66
FB79
FA6B
FA2B
FAAD
FB4F
FB82
FB1F
FA75
FA18
FA5D
FAF2
FB38
FB05
FAD7
FB27
FBBA
FBF0
FB9A
FB16
FAAC
FA57
FA4A
FACD
FB6C
FB22
F9F4
F97C
FAED
FD11
FD6E
FB69
F947
F984
FBDA
FDD8
FE2A
FE36
0016
03C9
0720
0815
06A0
046E
0367
044A
062C
0752
06D9
058B
04D7
053A
05F4
0622
05BC
0552
0524
04F3
0490
0449
0475
04E8
051E
04D5
044D
040A
0464
0528
059B
0537
0474
045A
0520
05BB
0539
0418
03A6
0451
0527
051D
0437
02FC
015B
FED4
FBD6
F9F2
FA3A
FBDA
FCEB
FC73
FB23
FA4A
FA8A
FB6F
FBFF
FBA2
FAB3
FA16
FA2D
FA75
FA5E
FA29
FA8B
FB7C
FBFF
FB75
FAAC
FAE5
FC00
FC7E
FB99
FA5F
FA3C
FB0F
FB98
FB4F
FAE5
FAF7
FB3B
FB39
FB38
FBAC
FC2C
FBDF
FB04
FB47
FDDB
01C3
04B5
0589
052E
0526
05B1
05EB
0548
0473
0480
0595
06AD
06B6
05B9
04B5
048C
052D
05D2
05D2
0538
049E
048E
0505
0576
055E
04CC
0450
0447
044A
0396
020D
008F
0004
003C
003B
FFA6
FF45
FFD1
00BA
00D5
000D
FF9A
0014
FFED
FCB8
F620
EF04
EB17
EB85
EE32
F022
F01F
EEF6
EDDA
ED42
ED27
EDA8
EEBF
EFBB
EF9A
EE3F
ECE2
ECEA
EE5A
EFCD
F003
EF26
EE5D
EE73
EF2D
EFD7
F00C
EFE9
EFC0
EFC0
EFDC
EFF2
EFF6
EFF4
EFED
EFCE
EF8D
EF5A
EF89
F024
F0BA
F0A4
EFB0
EE56
ED5C
ED56
EE54
EFA9
F020
EF07
ED3F
ECB4
EE3F
F07B
F13F
F012
EE96
EE71
EF6C
F022
EFF9
EFA6
EFC8
F001
EFD7
EFA7
F011
F0D7
F11E
F099
EFE5
EFAA
EFEE
F05A
F0B1
F0D5
F0A6
F033
EFEC
F045
F118
F1BC
F1DD
F1E2
F23C
F2A7
F298
F232
F239
F2F0
F372
F29B
F0B6
F027
F3C0
FBE1
053D
0B3B
0BF4
098F
07A0
07B1
08B2
0920
08C5
083A
07BC
073F
073A
082B
0969
097D
082A
070A
077F
08D9
096E
08D9
0821
07E8
079B
069B
0545
045A
03D1
031A
0243
0213
02CA
0398
03B5
0355
030D
02E6
02B0
029F
02E4
031F
02E4
0284
028A
02CB
029D
020E
0210
0321
0448
0438
032F
02BB
0392
048C
0457
034B
02C0
0333
03E4
040C
03A4
031B
02F2
03A2
054A
074C
089D
08BB
0826
07C9
07F5
0846
0864
086C
0880
086B
0807
07A2
0797
07CE
0806
083C
0886
08BF
08B4
0860
07DD
0773
07BE
0910
0A3D
08B7
02DF
FA55
F328
F030
F09B
F17B
F14C
F0EB
F156
F206
F206
F176
F0FB
F097
F00D
EFD0
F063
F125
F0DF
EF99
EEE0
EFC7
F164
F20E
F190
F126
F15E
F160
F0A6
F021
F0B7
F1A1
F17C
F066
EFD3
F07D
F189
F1DC
F16C
F0EB
F0C6
F0F6
F17C
F245
F2BF
F248
F143
F108
F233
F3A1
F3D0
F2C3
F1E1
F220
F31E
F3ED
F426
F3F9
F3AD
F35D
F31E
F318
F361
F3C6
F3EC
F3AC
F346
F31B
F354
F3BF
F403
F3F6
F3B6
F372
F33E
F33E
F3BD
F4AE
F53A
F48A
F31A
F275
F353
F49D
F4DE
F417
F36A
F376
F3D7
F440
F4EF
F5A3
F510
F2BE
F0F9
F34A
FA4E
0246
06BE
06EB
0581
0504
058C
0603
0616
0636
067D
0689
063C
05F4
05E5
05E3
05F4
0674
073E
077C
06D0
0622
0673
0757
076D
0658
0559
05A4
06C0
0737
067F
057B
050F
0514
0519
0587
0722
0990
0B4F
0B5E
0A71
0A13
0ACD
0BBF
0BDB
0B23
0A68
0A39
0A78
0AD6
0B3B
0B8D
0B84
0B02
0A76
0A63
0AA6
0A9C
0A16
09B5
0A02
0A9B
0AA7
0A0F
09A3
09E4
0A40
09D9
08DA
084A
08A9
095F
09B2
09A3
0966
08A0
06F8
0521
0479
0541
0602
0564
040D
03D1
0519
0635
05AB
043A
03AA
044C
04D2
049C
04B5
05B0
05A0
01D4
FA9A
F3D0
F106
F1E6
F35F
F381
F2FD
F304
F345
F2CF
F1F0
F1D7
F2A1
F304
F240
F145
F14A
F210
F27E
F267
F2A7
F389
F43B
F412
F3A1
F3CF
F46B
F47C
F3E2
F3AC
F474
F54D
F50F
F411
F3BE
F4A6
F5C9
F5F7
F539
F48F
F4B4
F570
F600
F5E3
F543
F4BB
F4D3
F57F
F60E
F5CE
F4EB
F450
F497
F549
F58C
F544
F524
F59D
F635
F609
F4D8
F35C
F29D
F2F1
F3B5
F411
F3E1
F3AA
F3D7
F43E
F48B
F4C0
F516
F57D
F59D
F55F
F534
F56F
F5AD
F550
F480
F40D
F442
F494
F4A3
F4BE
F516
F539
F4EC
F4D5
F56B
F5C4
F4C8
F3A1
F590
FC12
0415
08A4
0873
0713
0832
0B58
0D87
0D94
0D05
0D2F
0D86
0D26
0C85
0C9F
0D3C
0D47
0C9E
0C53
0CE5
0D62
0CF5
0C4F
0C87
0D4B
0D5E
0C78
0BA6
0BB5
0C3F
0C71
0C27
0BEA
0C19
0C85
0CC2
0CA6
0C48
0BCC
0B5D
0B1C
0B02
0AEF
0AE5
0AD9
0A56
08E8
0719
063C
06CC
07A9
078D
06BC
0677
0717
0798
071A
0626
05EF
06B2
0780
078F
0719
06BA
069E
06A7
06DE
0730
073C
06DA
0679
0687
06CF
06ED
06EA
0704
070A
06A1
05FA
05B6
0609
065A
0622
05CD
063A
0794
0945
0AE7
0C5B
0D0C
0C5B
0B2B
0B6D
0D1F
0CF0
079B
FE53
F649
F370
F4CE
F67F
F65D
F569
F526
F56C
F55F
F520
F54E
F5B4
F5AD
F55C
F575
F601
F647
F5E9
F55C
F51D
F51F
F532
F582
F62B
F6AA
F654
F561
F4D1
F514
F573
F534
F4A5
F476
F4A3
F4AF
F48F
F498
F4D2
F4EE
F4DC
F4D1
F4D2
F4A9
F469
F492
F558
F613
F5EE
F516
F490
F4DE
F560
F56B
F542
F56D
F5BF
F5AC
F53B
F4F1
F503
F535
F562
F59D
F5C5
F577
F4AC
F414
F474
F5B3
F6EE
F783
F78C
F75C
F703
F6A5
F69B
F6F1
F741
F761
F7A1
F805
F7F7
F74A
F6D6
F758
F815
F7B6
F677
F63D
F7BB
F8CB
F731
F4BF
F66F
FE7B
08DD
0F4D
0FCB
0DBF
0D17
0E35
0F06
0E85
0DC3
0DEE
0EA1
0EA7
0D81
0BA5
09BF
084F
07AB
07C9
0822
084F
087E
08F6
0976
0991
0960
0959
0983
095C
08AF
080D
0828
08DC
0959
0925
08A7
0870
0881
0886
086F
086E
0899
08E9
095E
09CE
09CF
0929
0854
080E
087B
08EC
08B0
07FF
07E1
0924
0B86
0DD8
0EFB
0EB4
0DC8
0D4A
0DA4
0E3D
0E45
0DC4
0D78
0DB1
0DD1
0D43
0C5C
0BE0
0BFC
0C40
0C67
0CA0
0D00
0D3A
0D26
0D2D
0DA0
0DFE
0D85
0C76
0BDE
0C0D
0C2F
0BC4
0B8E
0C31
0CD9
0C62
0B82
0C1B
0DE2
0D39
06F7
FCE8
F4D3
F288
F43A
F57D
F49A
F363
F39B
F488
F493
F3CE
F392
F443
F4C7
F458
F3C2
F431
F56B
F625
F5CE
F527
F503
F53E
F537
F4DC
F4AF
F4F8
F55A
F554
F4F0
F4B3
F4E6
F543
F55F
F535
F525
F575
F608
F68E
F6E9
F738
F782
F787
F712
F66D
F62D
F67E
F6ED
F705
F6E2
F6F8
F76A
F7E5
F80E
F7DF
F795
F76A
F786
F7EF
F868
F877
F7E0
F71B
F6EA
F76C
F7F7
F80B
F7FC
F852
F8E4
F8FD
F85B
F796
F76D
F7FD
F8BE
F91C
F8DB
F815
F72B
F6A0
F6AE
F6F0
F6DC
F694
F6AB
F71D
F735
F6CA
F6B6
F776
F7FD
F717
F5EC
F7B6
FE17
0660
0BC1
0C38
0A2F
0916
09A8
0A4C
0A05
0981
098B
09DF
09E4
09A8
0992
0994
0959
090B
092D
09A0
0993
08CB
0855
095A
0B9C
0DC1
0EDB
0F16
0EF6
0EA5
0E17
0D83
0D46
0D78
0DBD
0DA5
0D2E
0CD2
0D06
0DB7
0E4C
0E3E
0DB4
0D72
0DF3
0EB4
0ECB
0E1E
0D8F
0DBF
0E40
0E4F
0DDB
0D66
0D33
0D22
0D23
0D51
0D9D
0DD3
0E07
0E81
0EFD
0E72
0C3C
0963
07D5
082B
0906
08F9
0849
0820
08B2
091C
08CF
083A
0800
0825
0854
0871
088D
0892
0863
0844
0891
0915
0934
08C9
0845
07C3
06F5
0641
06CD
088A
08FB
0569
FE53
F789
F478
F4FB
F652
F690
F61F
F61A
F688
F6C6
F6C1
F6D4
F6EB
F6A2
F61A
F5E5
F62C
F67E
F680
F657
F656
F691
F6D9
F6F9
F6DF
F6A2
F67C
F6A5
F70C
F740
F6F6
F696
F6DF
F7D1
F88B
F86E
F7DE
F790
F798
F7A1
F7A3
F7D3
F823
F846
F826
F7E3
F781
F6E9
F64E
F623
F679
F6BB
F676
F61C
F65E
F6FC
F712
F6A1
F6A0
F73D
F753
F694
F71C
FB5A
029E
0916
0B9E
0ABF
0956
0922
099C
09C4
09A6
09AD
09AC
0961
0931
0984
09FF
0A41
0AD9
0C88
0ED1
1034
1009
0F3E
0F0A
0F76
0FB3
0F7A
0F44
0F3A
0ECF
0DD2
0D13
0D4D
0DF8
0E02
0D4E
0CBA
0CCD
0D28
0D45
0D40
0D82
0E0B
0E55
0E01
0D5B
0D11
0D6D
0E09
0E4F
0E20
0DD2
0DA0
0D42
0C38
0A96
092E
089A
0879
0834
0839
0948
0A57
0885
0253
FA28
F47B
F35D
F4CD
F59A
F4F2
F45E
F4FA
F60F
F68A
F688
F6B8
F704
F6C9
F5F5
F51C
F492
F437
F408
F43A
F4B8
F50A
F4ED
F4AF
F4C1
F529
F5A7
F63F
F735
F85D
F8FE
F8A7
F7D4
F755
F75C
F776
F74E
F704
F6E9
F723
F78C
F7C7
F79D
F756
F764
F7BD
F7DB
F796
F787
F835
F929
F958
F887
F7AC
F7A4
F816
F83B
F841
F8CD
F95C
F8C4
F7D1
F9A4
0004
0837
0D32
0CEC
0A36
08FE
0A08
0B37
0B0D
0A4D
0A29
0A6F
0A5F
0A1D
0A39
0A7C
0A4D
09EE
0A30
0B13
0BAA
0B79
0B1E
0B44
0B85
0B0E
0A02
0972
09DE
0A65
09FB
08D9
0827
088F
09C4
0B3D
0CBA
0E06
0ECD
0EF0
0EBA
0E9C
0EC8
0F0C
0F1D
0EE9
0E97
0E3B
0DB4
0D04
0C90
0CBC
0D52
0DA6
0D66
0D14
0D4D
0DCC
0DB9
0D25
0D6D
0F10
0FAE
0BC2
02FD
F9BC
F502
F58F
F7D6
F855
F6D8
F54F
F4D9
F4F3
F4F9
F514
F57A
F5C6
F5A6
F57B
F5AF
F5EE
F5BD
F55E
F570
F5EC
F639
F629
F62D
F679
F69B
F633
F5A3
F596
F5FA
F60A
F580
F524
F5C8
F71E
F80F
F7FC
F734
F650
F5AB
F569
F5A0
F652
F751
F830
F878
F824
F7D7
F82A
F8D0
F8DB
F806
F73A
F770
F860
F8F0
F8D9
F8EC
F968
F929
F7C9
F7E7
FD10
06C6
0F96
1286
105F
0E14
0EA9
1092
110A
0FF6
0F3E
0FA0
101A
101E
1062
10EC
1036
0D84
0AAD
09FC
0B0A
0B68
0A24
08E2
0938
0A66
0AA7
09E1
0998
0A6F
0B2E
0AB9
09CB
09C3
0A86
0ACE
0A31
099F
09CF
0A48
0A58
0A33
0A7F
0B15
0B1F
0A62
09D3
0A50
0B2F
0AE7
0931
07C6
0872
0AEA
0D35
0E01
0DD0
0DAE
0D94
0CEA
0C33
0CCD
0E64
0DD1
0831
FF0E
F7BB
F5E5
F7E6
F957
F84C
F68E
F632
F6D0
F6D8
F638
F633
F70C
F76B
F689
F58D
F5E5
F72D
F7D8
F77B
F730
F7D5
F8DF
F93C
F8A2
F7A0
F6CD
F651
F627
F646
F680
F68D
F664
F649
F64D
F61C
F591
F523
F552
F5E2
F626
F5DA
F567
F55A
F5E7
F6D2
F798
F7D4
F797
F753
F755
F77E
F784
F76A
F77A
F7CB
F811
F803
F7BD
F773
F740
F7D5
FAE3
017B
09C4
0FB0
10EA
0F47
0E67
0F7E
10B7
106D
0F77
0F86
106B
1080
0F61
0E97
0F2B
101B
100C
0F77
0FBC
10DA
1172
10EA
1040
106A
10E7
1097
0F69
0E5D
0E12
0E3E
0E8C
0F0B
0F5F
0E7F
0C23
09AE
08C6
0954
09D6
0980
0900
090F
092B
0884
0785
076C
0866
091B
0890
07B1
081B
09C4
0AF3
0A98
099F
0972
09FD
0A1F
09BD
0A19
0B80
0B99
076A
FF45
F780
F468
F5E4
F81F
F823
F6B5
F63B
F73B
F816
F7B6
F70C
F764
F85C
F891
F7C8
F740
F7BC
F864
F827
F75B
F722
F7AF
F81F
F7E6
F78E
F7B3
F815
F814
F7BB
F7A2
F7F1
F828
F7FE
F7DD
F819
F84A
F7FC
F7A2
F814
F927
F997
F895
F6EA
F620
F6B5
F7B2
F805
F7B2
F779
F79D
F7AC
F757
F6EE
F6D1
F6D4
F6AD
F6A8
F73E
F805
F7D7
F69F
F68C
FA5F
0203
099B
0CF7
0BCC
099F
0988
0B17
0BE2
0B17
0A28
0A36
0A63
0979
0833
0895
0B20
0DF5
0F33
0F1F
0F39
0FE5
1023
0F5E
0E68
0E50
0EF7
0F6E
0F4E
0F0E
0F12
0F11
0EBA
0E53
0E61
0EE2
0F66
0F97
0F5F
0EAE
0DA0
0CD8
0D21
0E73
0FBC
0FF9
0F52
0EBF
0EA9
0E7A
0D96
0C38
0AF8
09F1
0904
0892
0926
0A4B
0A9A
0984
0888
0978
0B91
0B64
0673
FE5A
F780
F4B6
F4E3
F530
F481
F410
F506
F6B7
F798
F73C
F69D
F6B0
F760
F7F6
F7FC
F780
F6D0
F638
F5F3
F61D
F69B
F734
F7C2
F82F
F861
F85D
F865
F8BF
F92A
F8F9
F7FE
F715
F757
F8BC
F9F9
F9E5
F8C5
F7DF
F7F5
F888
F89F
F7F8
F723
F6AE
F6B2
F715
F7E0
F8F4
F9C5
F9D2
F94C
F8E4
F8E4
F8CB
F839
F7DB
F8B3
FA62
FAEE
F91C
F6B9
F771
FCEB
04A7
0A55
0C03
0B53
0AD7
0B3B
0B70
0AD1
0A10
09FC
0A60
0A90
0A82
0AA9
0B0D
0B2F
0AD6
0A61
0A3C
0A4C
0A35
09E7
09A6
09A2
09D4
0A2C
0AAB
0B18
0B0E
0A81
0A1D
0AB0
0C41
0DF5
0EEE
0F14
0EF1
0F00
0F40
0F66
0F60
0F68
0FA2
0FCC
0F82
0EC6
0E0B
0DB3
0DAE
0DB3
0D9D
0D7E
0D62
0D50
0D69
0DC4
0E13
0DC8
0D0B
0D08
0E69
0F80
0D0D
05BA
FC59
F5B7
F42F
F5D8
F727
F692
F53E
F4BF
F539
F5CC
F5FF
F608
F61C
F61F
F5EF
F59B
F544
F51A
F54B
F5CE
F640
F645
F600
F5F6
F662
F6EB
F715
F6DA
F69F
F6AC
F6EF
F74C
F7D1
F866
F89C
F81A
F713
F620
F5B8
F5F9
F6CC
F7E6
F8D3
F93D
F939
F933
F97C
F9F7
FA31
F9C7
F8DC
F815
F807
F88F
F8E5
F881
F7D9
F7DE
F894
F8D2
F818
F843
FC35
0445
0CF3
11F1
1220
0FE9
0E37
0DF8
0E7B
0F12
0FA9
102B
103B
0FAA
0E8F
0CF1
0AE9
0940
090F
0A4E
0B89
0B8F
0AD3
0A75
0A8C
0A46
0982
091F
098C
09F1
0970
08AB
08F7
0A4F
0B11
0A39
08D0
086D
0921
09C8
09EC
0A26
0AC6
0B2A
0AC3
0A0F
09EB
0A43
0A23
0933
0896
09BB
0C78
0EF8
0F9C
0EA5
0DAE
0DCB
0E85
0ED1
0EBC
0F64
10CB
1076
0B7D
0255
F963
F4FB
F551
F712
F77A
F6C1
F68D
F73D
F7BF
F775
F716
F763
F7F3
F7E2
F71D
F654
F5FF
F603
F635
F686
F6DF
F71B
F739
F736
F6F1
F661
F5E4
F5E8
F65F
F6BC
F69F
F646
F620
F632
F642
F673
F71B
F7DF
F7D3
F6D0
F603
F67A
F7B0
F838
F79A
F6CF
F6ED
F7E6
F8CE
F906
F8D8
F8E9
F94B
F951
F86B
F714
F697
F7B0
F958
F9B0
F8B6
F96F
FEF4
0835
101B
12B3
1121
0F7F
0FE8
1100
10E7
0FCD
0F0B
0EF7
0EDB
0E94
0ECA
0F7C
0F99
0EB3
0DE5
0E3D
0F2C
0F70
0EE9
0E6A
0E4A
0E2C
0DE8
0DB9
0D74
0C83
0ADE
0973
0905
0921
08EB
0892
08E8
09A6
098B
087C
0812
0919
0A09
0955
0829
08D4
0AC0
0A1F
0473
FC3C
F693
F5A3
F6E2
F6F0
F598
F500
F611
F754
F73B
F622
F598
F677
F811
F909
F8C8
F809
F7EB
F896
F91C
F8BB
F7D3
F75C
F7B7
F86D
F8FF
F96C
F9C0
F99A
F8C2
F7F8
F843
F95F
F9D3
F8F7
F805
F858
F96E
F995
F856
F713
F724
F81E
F88E
F815
F830
FAB7
FFD5
05A3
09B6
0AFE
0A61
09B0
09E4
0A62
0A1A
093E
090F
09FA
0ACF
0A6D
0962
0921
09F8
0AC3
0A8B
09B2
0940
0997
0A27
0A4F
0A05
09A4
0977
099A
09EE
0A08
09AF
097C
0A5E
0C44
0DF5
0EA4
0ECA
0F1D
0F6A
0F2A
0E90
0E21
0DC7
0D3D
0D19
0E28
0F47
0D39
0631
FD0C
F723
F694
F85A
F8B1
F77D
F705
F7DD
F85F
F7A8
F6F8
F799
F8E5
F959
F8D0
F875
F8C7
F8F0
F853
F78D
F753
F762
F755
F77F
F80E
F833
F746
F612
F5ED
F6CE
F772
F73A
F6E0
F715
F771
F754
F728
F7A1
F82A
F782
F602
F5A4
F70D
F82D
F74A
F63E
F8B2
FF63
06D8
0B4A
0C82
0D11
0E92
1021
106A
0FCA
0F89
0FDB
0FC3
0ED1
0DE7
0E0D
0F1E
0FFB
0FCB
0EC7
0DEA
0DD9
0E38
0E42
0DDF
0DC8
0E7C
0F94
1048
1061
1035
0FE5
0F3A
0E48
0DC0
0E07
0E45
0D13
0A5C
07E6
076F
089E
097D
08E4
07C8
07EC
097E
0A57
07D4
01A3
FA89
F5FB
F4FB
F5AC
F5E4
F57D
F5AA
F6BB
F78E
F740
F683
F68E
F73D
F749
F64F
F582
F5E6
F6E6
F755
F726
F731
F7BE
F831
F810
F791
F71E
F6CA
F680
F65C
F68B
F704
F7A3
F871
F946
F981
F8B9
F7A5
F75C
F7AC
F772
F6C4
F732
F90E
FA17
F8A4
F723
FA3B
02E4
0C54
110B
10D9
0FEF
10B9
112B
0EDE
0B38
097E
0A3E
0B07
0A4F
0956
09C1
0B08
0B59
0A41
0919
090E
09B9
0A0F
09CA
0950
08EF
08D9
0951
0A39
0ADF
0AD0
0A69
0A14
0989
0890
07E0
0858
097F
09EF
0984
09FD
0C8B
0F7E
1008
0E2B
0D15
0E91
0FB5
0BFB
0325
FA24
F5CB
F600
F71B
F6CE
F61C
F6B3
F80F
F869
F784
F700
F7E3
F913
F8E5
F771
F675
F70D
F863
F8EB
F854
F7B5
F7F6
F8A6
F8A4
F786
F606
F518
F4FE
F54E
F59D
F5E9
F65E
F6EE
F742
F71E
F6BD
F6A3
F6DD
F6D1
F623
F594
F633
F793
F7CF
F625
F503
F81A
FFEC
084C
0C51
0B69
0952
0932
0A54
0A60
0942
092C
0B42
0DF9
0F39
0EEA
0E88
0ED6
0F15
0E86
0DA9
0D7B
0E1F
0EE3
0F30
0EFA
0E7A
0E0D
0E08
0E5C
0E9A
0E9F
0EC6
0F30
0F3B
0E62
0D51
0D4B
0E56
0EDF
0DE7
0CBB
0D47
0F07
0F5F
0D59
0B34
0AEF
0AB6
06DD
FF1E
F7CE
F506
F619
F71D
F61E
F4D5
F532
F651
F612
F475
F398
F4AC
F681
F754
F6E1
F62D
F5EF
F603
F61D
F64A
F697
F6C5
F6B3
F6A5
F6D7
F71C
F735
F741
F76F
F79E
F7A7
F7C5
F83B
F8BD
F8C2
F866
F85D
F8CE
F8E9
F81F
F753
F7C7
F8FA
F8F7
F772
F75D
FC09
04D3
0D0B
109F
0FF7
0E93
0EAB
0F6D
0F4F
0E84
0E52
0EF3
0F5B
0ED4
0DBD
0C9E
0B67
0A00
08FB
0907
09E0
0A70
0A21
0971
091B
092B
0947
0960
0996
09C3
09A4
095F
095A
09A2
09DB
09CE
09AC
099A
0964
08F6
08B3
08DC
08DA
080B
0727
07B7
0981
099E
055B
FDCA
F744
F503
F623
F762
F721
F685
F6FE
F81C
F877
F7D2
F745
F787
F81E
F846
F7F4
F79A
F76E
F75B
F76B
F7D1
F87C
F8E4
F894
F7BB
F710
F722
F7DB
F89A
F8BA
F833
F7AA
F7BC
F825
F805
F719
F63F
F654
F6F2
F6F9
F648
F61D
F723
F800
F6FA
F50D
F5D9
FBA2
040F
0A22
0B4F
09A1
08AF
0989
0A89
0A5C
09AD
099D
09F0
09AA
08D7
087B
08F5
097A
0977
09AD
0B27
0D8F
0F47
0F50
0E60
0DD6
0E1B
0E8B
0E96
0E5F
0E50
0E89
0EC8
0EB7
0E49
0DE9
0E16
0EB6
0F00
0E65
0D75
0D4F
0E0A
0E5F
0D85
0CC9
0DE1
0FB0
0E54
077D
FDD2
F6A7
F496
F58A
F61A
F573
F516
F5D6
F6AA
F690
F609
F5FB
F62E
F5E4
F552
F556
F601
F65D
F5D7
F50C
F4EB
F581
F60B
F5F9
F577
F50B
F50B
F582
F627
F66A
F601
F58A
F5EC
F6F0
F748
F672
F5B8
F684
F843
F91B
F893
F830
F8EF
F968
F7E1
F5D5
F77B
FEE8
08DC
0FB2
1108
0F5C
0E65
0F2E
1032
101B
0F42
0EA9
0E91
0E91
0E7E
0E92
0ED7
0EF3
0EB9
0E78
0E8A
0EBC
0E5E
0CF9
0AF4
0963
0910
09A1
0A01
099D
0902
08FD
0965
0942
0844
077C
0814
0995
0A3F
0945
07FB
081C
095F
09CF
08A8
07A8
089B
0A2A
089B
023C
FA01
F4D6
F498
F6BC
F7C4
F6F4
F60B
F63F
F6E7
F6F7
F698
F697
F703
F741
F71C
F6F8
F70C
F713
F6EB
F6E8
F740
F78D
F743
F695
F653
F6DC
F7AD
F81A
F7F6
F777
F6EA
F6CA
F775
F86C
F894
F7A5
F6D1
F735
F822
F7EF
F675
F589
F643
F707
F5D1
F407
F5DF
FD17
05F5
0B05
0AEA
0900
08B5
0A0A
0AF3
0A94
09D7
0992
097D
0936
090C
093C
095C
0927
092D
09E8
0AB4
0A93
099C
08CD
08AE
08F0
0969
0A8F
0C83
0E5A
0F01
0E9E
0E46
0E63
0E55
0DDB
0DAD
0E3D
0EB8
0E51
0DB6
0E16
0F04
0ED0
0D40
0C7F
0E1E
0FE4
0D60
0530
FB60
F58D
F543
F746
F7F1
F6D5
F5DA
F606
F676
F611
F522
F4BE
F536
F5C9
F5CC
F568
F530
F553
F58D
F5A7
F5AF
F5C4
F5E5
F600
F614
F62C
F647
F659
F655
F638
F608
F5D9
F5C3
F5CD
F5FB
F65F
F703
F79D
F7AF
F71D
F692
F6D3
F792
F784
F657
F629
F9F2
01FC
0AAD
0FAB
0FF7
0E4F
0DAF
0E61
0EC8
0E2B
0D88
0DDC
0EAB
0ED7
0E31
0D84
0D64
0DA6
0DDC
0DDD
0DBE
0DA3
0DAA
0DBA
0D8B
0D08
0CAD
0D1F
0E2A
0E88
0D34
0ACC
08FD
088B
08A4
0859
07DC
07C7
07F9
07F0
07DC
084E
08FD
08F0
0825
0807
093C
09B0
064C
FEF6
F783
F3D5
F3FE
F518
F525
F4B7
F500
F5C5
F5E9
F538
F49B
F4C8
F57E
F633
F6CA
F74A
F780
F760
F756
F7A0
F7D7
F794
F73E
F782
F831
F85B
F7B3
F715
F741
F7AC
F751
F69E
F76F
FAD5
FF8F
034D
050A
0567
0534
049C
03C4
0343
0366
0388
0310
02D5
0488
0867
0C54
0DF5
0D51
0C8C
0D29
0E71
0EE4
0E61
0E13
0E87
0EE1
0E3C
0D19
0CC2
0D8A
0E66
0E50
0D72
0CB8
0C9E
0CD2
0CDA
0C98
0C37
0BEE
0C03
0C91
0D19
0C90
0A66
074A
04A1
032A
0284
0216
01EA
0265
0362
0423
0432
03E0
03BB
03DC
0404
0425
045B
0489
045B
03CB
034D
0345
0391
03C8
03C3
039A
0336
025D
0161
0168
036D
0707
0A78
0C34
0C29
0B85
0B69
0C02
0CC2
0D30
0D46
0D28
0CD9
0C5B
0BED
0BE3
0C32
0C5F
0C06
0B5C
0B0A
0B71
0C2D
0C81
0C1E
0B65
0AEE
0B08
0B89
0BDA
0B1D
08C6
055E
0275
015F
01E4
0287
0231
0159
0131
0203
02E2
02FE
02AA
02AF
0323
036C
0335
02E4
02ED
033B
0369
035D
0344
0323
02C5
022F
01B7
0192
01AC
0226
0391
0638
095B
0B9C
0C54
0C19
0BDF
0BE7
0BE3
0BCA
0C01
0C9E
0D0A
0CC7
0C26
0BDC
0C06
0C10
0B98
0AFC
0ACE
0B13
0B58
0B50
0B0A
0A9D
0A1A
09E3
0A84
0BB4
0BEE
09B7
0580
01AF
0060
014B
0254
01FB
00CA
0038
00BA
0173
018D
012F
00FC
011B
0132
0119
011F
0176
01D1
01C9
0171
013D
0169
01B4
01C1
0177
00F2
0072
007A
01C0
0486
07F3
0A74
0B20
0A8A
0A0C
0A51
0ADA
0AEF
0A9A
0A6F
0AAA
0ADF
0AA3
0A1D
09C7
09D8
0A22
0A6B
0A9A
0AA4
0A8A
0A6E
0A78
0A8D
0A58
09E2
09C5
0A59
0AC7
0984
062A
0259
0034
002A
00B4
0066
FF94
FF7A
004F
00F7
00AD
0011
0024
00CB
0119
00C1
0088
010D
01D8
0205
017B
00DD
0083
002B
FFC9
FFCA
003A
005D
FFCF
FFB1
01B0
05B2
0957
0A61
092E
0820
08BA
0A24
0AC0
0A47
09B8
09BD
09FE
09F6
09AF
0964
0907
088B
0852
08C6
099C
0A11
09E8
09A1
0994
0969
08EA
08B2
0947
09BE
0850
049B
0096
FEA8
FF06
FFCF
FF8C
FEBE
FE96
FF17
FF44
FECB
FE6D
FEC2
FF5A
FF8E
FF80
FFB2
FFFD
FFB8
FEF2
FEA4
FF45
FFEC
FF8D
FE90
FE52
FF22
FFBB
FF3D
FED3
007A
0453
081C
09A5
0925
087C
08C9
097E
09AE
0967
0951
099C
09D5
09B0
0969
094B
094B
0946
0950
096E
095B
08E8
087C
08A6
094A
09A3
0951
08EA
091C
096B
0876
059B
01F4
FF55
FE88
FEE6
FF67
FF9F
FF9F
FF68
FEF5
FE83
FE6B
FE97
FE91
FE2A
FDD5
FE0D
FEA1
FEEC
FEB3
FE57
FE20
FDCE
FD30
FCD0
FD5D
FE83
FEF1
FE09
FD22
FE57
020E
0634
0859
0826
0754
0760
0813
0865
0823
0801
0861
08C4
08A9
0853
084A
086F
082B
0779
0717
0778
0815
0828
07C7
07A1
07E9
0813
07CF
0796
07BF
077A
0586
01FE
FEB2
FD4C
FD9F
FE38
FE3F
FE14
FE3A
FE75
FE4E
FDED
FDD5
FE08
FE08
FDB0
FD79
FDAA
FDD9
FDA5
FD69
FDAD
FE35
FE4B
FDEF
FDEF
FE84
FEA2
FD7A
FC49
FD70
0179
05F6
0815
07B4
06FC
0759
07FF
07B2
06D2
06B7
0789
0807
077B
06DE
075D
0882
08D3
07F1
0708
0711
0788
0770
06E4
06D4
076A
07C1
075A
06F0
072D
0723
0530
0154
FDB6
FC62
FD1F
FE05
FDE7
FD54
FD41
FD9D
FDB1
FD56
FD19
FD4A
FD9E
FDCA
FDEF
FE29
FE26
FDAD
FD2C
FD3D
FDAA
FDA6
FD12
FCDA
FD91
FE4F
FDEA
FD05
FDD4
0153
0595
07BA
0744
0666
06F4
0832
084E
0723
0651
06C8
078C
0756
0675
0639
06E7
076C
0717
0697
06BF
0731
0716
069A
06B1
077A
07F0
0784
0714
0782
07D1
05FB
01BE
FD7C
FBB1
FC3D
FD0A
FCD6
FC5A
FCA4
FD6F
FDBD
FD5E
FD0B
FD27
FD3C
FCE9
FC87
FC85
FCA7
FC84
FC57
FC9A
FD12
FCF9
FC50
FC2B
FD2F
FE53
FE14
FCC5
FCB3
FF72
03B7
06AA
0703
0619
05C8
064B
0692
0620
05B1
0610
06FD
07A6
07BD
0793
0765
0715
069D
0648
0643
0653
063C
0639
0698
0715
0711
068E
066E
0724
0793
05EF
01FB
FDD0
FBE2
FC6D
FD79
FD49
FC29
FB90
FC0B
FCB4
FC9D
FBF7
FB95
FBB8
FBF9
FC11
FC38
FC8E
FCCF
FCC3
FCAC
FCD5
FCFD
FCB9
FC32
FBFA
FC1C
FBF1
FB55
FB84
FDE6
0202
0583
0698
05D9
0535
0590
061C
05FB
0586
0586
05E1
05C9
0515
0495
04EA
05AF
0628
0649
066B
067F
0628
0592
056E
05DE
061B
059E
0526
05B3
06A6
05F1
02A4
FE7E
FC22
FC29
FCCB
FC6D
FB82
FB69
FC3E
FCC5
FC47
FB8D
FBA2
FC5B
FCC4
FC87
FC27
FC02
FBD3
FB6C
FB36
FB8D
FC00
FBE7
FB73
FB79
FC0C
FC30
FB73
FB2C
FD2C
0150
0533
06B3
061E
0561
058E
0605
05F6
05A3
05AF
05F2
05C5
0536
0513
05AE
064B
062F
059E
0558
056D
0553
0508
052C
05CC
05F2
050E
042B
04A7
05EC
0594
0250
FDD4
FB0B
FAD8
FB87
FB77
FAF9
FB28
FBDE
FBFF
FB58
FAF8
FB8A
FC49
FC2D
FB75
FB32
FBA2
FBEB
FB97
FB51
FBBC
FC4A
FC18
FB66
FB46
FBE1
FC20
FB73
FB21
FCF6
00D5
0482
0600
0585
04AF
0486
04DC
0536
0580
05B5
059B
052F
04E2
050D
0561
0556
0505
0517
05BE
0645
0604
0553
0502
051A
04DE
0412
03A1
0461
0597
0559
02A4
FEAD
FBB8
FADB
FB3E
FB7A
FB1C
FAA9
FA8A
FA94
FA8A
FA97
FAFC
FB7B
FB7F
FAEF
FA6D
FA95
FB34
FB8F
FB56
FAF3
FAD9
FAFF
FB29
FB55
FB8A
FB76
FAE0
FA89
FBE9
FF82
03BC
062F
0618
04FC
04A9
053A
058F
0528
04B3
04D5
0542
0565
055D
05A0
05F3
059D
0499
03E1
041D
04B9
04CC
0470
0473
04FA
0547
0508
04EA
0555
052C
02E8
FEDE
FB68
FA55
FAF2
FB4B
FABF
FA61
FB00
FBE3
FBED
FB31
FAB0
FAD4
FB06
FACF
FA95
FAD6
FB49
FB57
FB13
FB04
FB31
FB1D
FAB6
FAA1
FB18
FB40
FA56
F958
FA73
FE62
0310
059C
0562
044B
0436
04F9
0549
04D0
0470
04BC
0516
04B7
03EF
03AD
0427
0499
0478
0432
0461
04D6
04E9
048E
0460
049F
04C4
0471
042B
0481
04B4
0327
FF77
FB73
F970
F9D0
FAE5
FB21
FAA9
FA7D
FAD3
FB04
FAC6
FA96
FAD1
FB04
FA9C
F9DD
F998
FA08
FA95
FAB8
FAA1
FAAF
FACD
FAC3
FAB6
FAE3
FAFF
FAA2
FA55
FB74
FE88
022A
0448
0466
03FC
0465
0546
056D
04B3
040E
041D
0464
0449
040E
0446
04C0
04B7
040A
038E
03DD
0475
0480
040A
03D0
040C
0430
03EE
03D1
0445
0472
02CF
FF16
FB0E
F8F9
F958
FAAB
FB38
FAAF
F9F8
F9DD
FA41
FA88
FA6E
FA3D
FA4A
FA81
FA8C
FA58
FA33
FA6B
FADA
FB12
FAE6
FAA2
FA95
FA91
FA39
F9D9
FA88
FD17
00E7
0426
0569
04E4
0400
03D5
0441
0478
0426
03BC
03C4
0432
0487
047C
043E
0414
03F8
03BC
0372
036D
03C3
040A
03DD
0386
03B2
044F
0422
01F1
FE1F
FAAE
F95D
F9F9
FACB
FAA2
F9EA
F9BD
FA4F
FAC9
FA82
F9D6
F98D
F9DD
FA49
FA6C
FA74
FAA5
FAD1
FA8E
F9F8
F9BF
FA4E
FB0F
FAFC
FA00
F97E
FB18
FEDC
02DE
04EA
0490
034E
02CE
034B
03D7
03D1
039A
03C6
042E
042C
03A2
0334
036B
03EB
03F9
037D
0323
0369
03F1
040B
03B9
03B3
0450
04B7
0384
0053
FC73
F9D0
F946
FA0A
FAB6
FAAB
FA5A
FA54
FA7B
FA51
F9D2
F997
FA00
FA9D
FAAE
FA24
F9B1
F9E7
FA7A
FAB7
FA74
FA30
FA41
FA49
F9DB
F96C
FA2E
FCCE
007B
0376
0496
042B
0374
0351
039E
03C0
0383
0348
0367
03B3
03BF
037D
0352
0385
03CA
03B4
035D
034E
03A2
03BB
0326
0277
02BC
03EA
045B
0261
FE44
FA48
F881
F8F9
FA0D
FA5C
F9E9
F97E
F989
F9CB
F9F2
F9FF
FA15
FA21
F9F6
F9A9
F98C
F9C5
FA0C
F9FA
F992
F953
F9A5
FA3C
FA56
F9B4
F951
FAA8
FE19
0230
04C5
04FB
03E1
032A
036A
03E2
03C7
0341
0303
0342
0382
035C
030C
0309
0354
0382
0366
0353
0391
03DB
03B4
033C
0334
03F6
0498
0386
0033
FBF7
F902
F860
F93A
F9F8
F9EC
F99B
F9A9
F9F5
F9F5
F99B
F967
F9A7
F9FD
F9E8
F97B
F949
F98F
F9DD
F9BB
F966
F984
FA2F
FA9A
FA09
F8FA
F90C
FB71
FF90
0354
04F8
047C
0359
02E8
0346
03B3
03B2
0381
0385
03AE
03A1
0356
032C
0359
0390
037B
0346
0361
03C7
03E1
0356
02B5
02DF
03BB
03EB
0216
FE72
FAC1
F8C1
F8AE
F967
F9BE
F981
F938
F949
F983
F989
F95D
F955
F997
F9DF
F9DD
F9A0
F981
F99A
F99A
F945
F8EB
F916
F9B2
F9F5
F968
F8D9
F9D9
FD04
0114
03E2
046D
0398
02F6
0327
0393
038A
032A
0305
0348
0387
0368
0320
031C
0364
0394
0373
0341
0356
0389
0361
02CD
0277
02FF
03E8
03A8
0115
FCDA
F92C
F7E6
F8DC
FA34
FA59
F968
F8A5
F8DA
F98F
F9D3
F970
F8FB
F8F1
F92B
F948
F942
F955
F975
F959
F90A
F912
F9B7
FA50
F9F5
F8DA
F898
FAA9
FEA5
0267
040D
03A4
02B5
027F
02ED
0338
031B
0301
0345
03A3
039C
0334
02F5
0336
039A
0383
02EE
028A
02D8
0376
038E
02F9
0291
0305
0396
0292
FF3E
FB0B
F85B
F830
F951
F9E9
F97D
F905
F951
F9ED
F9E8
F92B
F88F
F8B1
F933
F95E
F91B
F8F2
F92D
F972
F958
F919
F93D
F9B4
F9BC
F8EC
F820
F8EF
FBFD
0019
032A
0411
037D
02E2
02EF
0333
0316
02BB
02B3
031A
0367
0338
02E2
02FC
0377
039F
0316
0275
028E
0346
039A
02FC
0235
0274
0397
03DF
01B6
FD98
F9CA
F82F
F89C
F96E
F977
F8F4
F8BB
F900
F93A
F90E
F8CB
F8E6
F949
F973
F93A
F900
F91B
F94F
F92D
F8C6
F8B7
F949
F9DE
F99A
F89B
F844
F9FF
FDAB
0184
03A1
03A1
02BC
0264
02E4
0375
0363
02E4
02A9
02E7
0324
02FA
02AB
02B5
0304
030D
02A9
0277
02F7
03A0
0367
024B
01A9
0284
03DA
035A
0002
FB77
F872
F80C
F905
F992
F944
F8E6
F90B
F95F
F962
F922
F910
F94A
F979
F956
F913
F90C
F948
F96B
F930
F8D2
F8D0
F94C
F9C0
F97E
F8B9
F8CB
FB01
FF03
02BB
0438
0390
028D
0296
034C
0373
02C5
0236
0280
031D
031D
0281
0229
0287
0303
02E9
0274
026D
02F8
034B
02D9
023F
0289
039D
03E2
01D5
FDCD
F9E2
F808
F85B
F957
F99A
F91F
F8CA
F910
F979
F96D
F911
F902
F964
F9A3
F951
F8D4
F8EB
F996
FA00
F99C
F8F5
F8F1
F982
F99B
F8B3
F7E1
F8FE
FC94
00F6
03B5
03E9
02CF
023A
02B4
0354
0330
0286
0241
02B4
032F
0300
0269
023E
02B2
0318
02E5
0277
0286
0301
031E
0295
023A
02E4
03F1
038C
00AD
FC75
F935
F83C
F8E3
F99F
F999
F91B
F8D0
F8F1
F933
F94E
F94B
F95A
F981
F993
F972
F93B
F91F
F922
F913
F8ED
F8F7
F95B
F9AD
F94C
F876
F88B
FABB
FE8C
0201
037A
032C
0292
02AB
0325
033D
02E0
029F
02C7
0302
02E9
0296
027C
02C9
0326
0321
02C1
0283
02BD
0320
0317
02A3
027B
0315
039D
0277
FF0C
FAE1
F85B
F857
F970
F9CC
F91F
F889
F8D1
F97B
F9A3
F939
F8E3
F907
F956
F968
F94A
F947
F95E
F952
F921
F90A
F930
F95D
F93C
F8C2
F87E
F965
FC09
FFCD
0301
0432
0385
0287
0281
0333
0379
02F1
0268
028F
0301
02F1
0268
0229
0283
02EA
02E3
02C2
030A
037A
034E
0280
021D
02E6
0401
0396
00CA
FCBA
F979
F841
F8AE
F974
F9A0
F93A
F8E2
F8F9
F946
F95D
F933
F923
F960
F997
F96B
F911
F916
F97C
F997
F906
F86B
F8A5
F978
F9B7
F8EC
F861
F9E6
FD97
0172
0354
0311
0239
022A
02CF
033E
030D
02A9
029A
02D2
02E1
02A1
026B
0296
02F8
0316
02C8
027D
02AB
031D
0322
028D
0222
02A5
0377
02DA
FFDD
FBC9
F909
F8B9
F9A6
F9F6
F93E
F893
F8CB
F970
F99B
F947
F92F
F996
F9DE
F97C
F8C6
F888
F8EF
F961
F95D
F922
F935
F980
F95E
F898
F804
F8EB
FBBD
FF74
0257
035F
02FD
026D
0271
02C5
02C4
0261
0227
0271
02E0
02E9
0298
0283
02EB
0352
032C
02A9
0277
02CB
0318
02E0
027C
02AD
036F
0388
01AC
FDFF
FA44
F857
F886
F97B
F9BE
F91D
F895
F8E7
F9AD
F9F2
F97C
F8F7
F8F5
F92B
F90E
F8BD
F8D2
F960
F9AC
F93C
F8A9
F8DD
F9A4
F9C3
F8C6
F810
F980
FD32
012B
0354
0365
02B7
028F
0301
0359
0329
02A9
0252
0262
02BB
030E
0324
030B
02F6
02F0
02D6
02A1
0282
0298
02B6
02B1
02BF
0321
0366
026E
FF98
FBD2
F906
F850
F902
F9A6
F98E
F922
F8ED
F8EB
F8D9
F8BD
F8D9
F92B
F960
F941
F900
F8F2
F920
F946
F93A
F924
F942
F988
F995
F925
F8A1
F912
FB47
FED0
0217
03AC
0381
02BD
027B
02D7
033B
033C
0300
02D5
02C6
02B5
02A5
02B7
02E6
0303
02F0
02CA
02C6
02F5
0322
030A
02C0
02B7
031C
0333
01BA
FE55
FA68
F80A
F7FF
F90A
F977
F8F7
F893
F8EB
F972
F972
F926
F937
F999
F9A7
F934
F8D8
F8F7
F92A
F901
F8D6
F936
F9B8
F96A
F892
F905
FC00
003E
0319
0371
02A9
0296
035D
03D2
035F
02B0
0289
02C2
02D4
02B9
02BC
02C8
0292
0246
0269
02F5
0337
02D0
0267
02CE
039F
0349
00C9
FCFC
F9DC
F898
F8C1
F929
F925
F8D9
F8B0
F8D9
F939
F993
F9B3
F988
F938
F914
F949
F9A0
F9B0
F955
F8F0
F8EB
F929
F91B
F89D
F889
FA19
FD75
0127
0351
037D
02DA
02B7
0329
0364
030F
02A9
02AF
02E3
02C2
024F
020A
0225
0256
026E
02A9
0319
034A
02E9
0287
02F1
03BA
0326
001C
FBD8
F8E8
F883
F96D
F9BD
F91C
F89F
F8F1
F970
F954
F8E4
F8EE
F97B
F9C9
F97C
F928
F95A
F9B9
F9A7
F945
F937
F975
F92F
F84D
F842
FAA1
FEE9
02A1
03D9
0316
024E
0287
031E
032D
02D2
02AF
02DB
02E1
02A3
0287
02BC
02DD
02A0
0267
02A6
030F
02F6
0273
0279
035F
03E6
0252
FE8B
FA8B
F873
F883
F94E
F990
F949
F919
F934
F94C
F935
F91F
F92B
F935
F924
F927
F963
F997
F96B
F90C
F904
F965
F97A
F8CD
F83B
F95E
FCB2
00AC
0318
0345
0272
0227
02A2
031B
0315
02E3
02EA
0307
02F2
02C9
02D5
02F6
02CE
026E
0262
02D5
0337
02FF
0295
02D7
0399
0357
00D0
FCC3
F96D
F85A
F901
F9B8
F995
F905
F8D0
F90C
F93E
F92B
F911
F933
F979
F9A6
F9A5
F983
F93E
F8EB
F8D5
F934
F9B3
F99B
F8D2
F877
FA09
FDAB
0197
03B3
0396
02AC
026F
02EC
034C
0330
0300
0312
031C
02CF
0276
0287
02DC
02E7
02A1
02A3
031D
0365
02F5
026A
02B9
037D
02F0
FFFC
FBD4
F8E6
F84D
F8FD
F960
F91A
F8DA
F900
F93D
F94D
F960
F996
F9A7
F964
F928
F963
F9CD
F9AD
F8EA
F868
F8D9
F9A6
F9A0
F8C6
F8B9
FAFC
FF0B
02A9
0418
03A0
02DE
02DC
034C
036D
0324
02DF
02D2
02CA
02B1
02BC
02F9
030E
02BF
0273
02B3
034A
0368
02DC
028E
0334
03D0
026E
FE9B
FA61
F843
F897
F983
F972
F8B8
F88D
F92E
F9B6
F991
F928
F911
F930
F92E
F92E
F984
F9E9
F9C7
F937
F910
F9A6
FA11
F96F
F882
F947
FC9A
00DE
038D
03D6
031B
02F5
0377
03AD
0333
02A7
02AA
0307
0332
0310
02F4
02F7
02DD
02A3
02AD
0318
035C
02FB
026E
02A8
038F
0383
0111
FCE0
F95B
F83B
F8E7
F989
F948
F8DB
F90A
F988
F997
F937
F915
F96D
F9BE
F9A4
F973
F999
F9D4
F99C
F91B
F916
F9AE
F9FA
F95A
F8D2
FA39
FDE8
01EE
03F5
03A3
02A7
0294
0351
03C6
0383
0318
0312
0339
031B
02C8
02AB
02D2
02E3
02C3
02CA
0324
0363
031E
02B7
02E7
0363
02AC
FFC2
FBC5
F917
F8DA
F9CF
FA16
F95E
F8D0
F923
F9AB
F98C
F90D
F90F
F9A5
FA00
F9C1
F987
F9D1
FA1F
F9BF
F910
F90F
F9C3
FA0A
F968
F93A
FB45
FF40
02CA
03F9
0356
02C1
030F
0383
0360
0300
0310
0372
0383
0325
02DF
02EE
02E5
0284
024E
02CF
0388
0378
02A1
024C
0337
0419
02BF
FEC4
FA6A
F850
F8BF
F9C4
F9BE
F8FF
F8C4
F94D
F9BC
F98B
F93C
F966
F9CC
F9DD
F9AD
F9C5
FA23
FA26
F9A3
F959
F9CC
FA3A
F998
F87B
F903
FC55
00DD
03CF
0427
035A
032C
03B2
03E5
0370
030A
032D
0363
0322
02BB
02C9
032A
0337
02D9
02B2
030B
0349
02E2
0269
02E4
0414
042A
01B2
FD75
F9E5
F8A1
F913
F994
F95B
F8EE
F8F9
F95E
F997
F98A
F98D
F9BF
F9D6
F9AE
F996
F9CF
FA07
F9D2
F971
F992
FA2E
FA4A
F95C
F898
F9FA
FDDC
021A
042E
03D5
02F2
0310
03C9
03EC
035C
0304
0350
03A1
0361
02E5
02D1
0310
0313
02D7
02EC
036A
0394
0302
0284
0311
0404
0366
0039
FBF8
F92B
F8CF
F9A5
F9FF
F992
F932
F958
F99A
F988
F95E
F986
F9E5
FA09
F9E6
F9D9
F9FC
F9EB
F96F
F90F
F968
FA1C
FA1D
F94C
F942
FBA8
FFF3
0386
046D
0363
02A2
032B
03F5
03D5
0325
0307
0392
03C7
0336
02AE
02EF
037E
0376
02FF
02FC
0388
03B2
030C
0293
0334
03E8
0283
FE89
FA3C
F83D
F8BB
F9C2
F9DE
F96F
F961
F9AD
F9B1
F96A
F975
F9F3
FA33
F9C7
F940
F95A
F9DE
F9FE
F9A3
F992
FA1A
FA6A
F9C0
F8E5
F9B5
FCF7
012D
03FC
0484
03DD
037A
039B
03A4
0355
031E
0357
03B3
03BF
038D
037F
0399
037D
0323
0305
0363
03B2
0354
02B2
02E1
03E4
040F
01B9
FD71
F9BC
F87E
F927
F9CC
F98B
F927
F96F
F9FB
F9EC
F950
F900
F957
F9BF
F9AC
F969
F98A
F9F3
FA08
F9B7
F997
F9E6
F9F9
F953
F8E2
FA5C
FE1C
0246
0487
0467
0377
0348
03DC
0437
03F2
0391
038C
03AE
0395
0361
0371
03B2
03BA
037E
036E
03AF
03C8
0366
0319
0395
044A
0382
0051
FC12
F93A
F8D3
F9A0
F9E5
F95B
F8F5
F937
F9A0
F9A3
F97A
F99D
F9E8
F9D7
F970
F946
F991
F9C7
F980
F935
F98A
FA27
FA0B
F92E
F927
FB81
FFAF
0352
049D
0406
0351
0370
03DF
03E2
0395
0386
03B6
03B2
0367
0350
03AC
0409
03ED
0397
039B
03EC
03E3
035C
032B
03D6
044F
02C0
FEDB
FAAA
F891
F8DE
F9D7
FA03
F998
F98B
F9F5
FA1B
F9B2
F957
F98B
F9F5
FA00
F9C5
F9BD
F9DD
F9A6
F923
F917
F9D3
FA76
FA01
F914
F9AB
FCD8
0134
042E
04AA
03C9
033C
0370
03BF
03B8
03A0
03C0
03E0
03B9
037C
0382
03B0
039A
034A
034E
03D4
0434
03D1
0324
033E
0419
0412
01A8
FD7B
F9F0
F8C4
F96C
FA1F
F9FD
F991
F989
F9B7
F9A8
F97F
F9AC
FA0E
FA12
F99F
F956
F99C
F9F7
F9CD
F971
F9AB
FA58
FA56
F943
F8AC
FA91
FED5
02F9
04A8
040B
0323
034A
03FC
041D
0396
033C
0380
03F3
040E
03E7
03D9
03E6
03D2
03A7
03AF
03E3
03CC
0341
02E3
0362
0434
03AA
00BE
FC8C
F97B
F8DE
F9C8
FA62
F9FC
F968
F97A
F9EA
F9F1
F97E
F93B
F97C
F9D4
F9CF
F99F
F9AB
F9DE
F9DE
F9C1
F9ED
FA4C
FA3C
F9AC
F9CE
FBF1
FFB0
02FB
0432
03C2
0348
038E
0400
03FB
03BD
03D3
041C
040E
03A9
0388
03E5
042D
03E0
0363
036C
03DA
03D8
033D
02FF
03C0
0461
02EF
FF13
FAEC
F8F3
F963
FA5B
FA4B
F993
F96C
FA01
FA62
FA0D
F995
F99E
F9E1
F9CF
F98F
F9B1
FA22
FA29
F99F
F95C
F9EF
FA85
FA05
F91F
FA00
FD98
0200
046F
043E
0337
0317
03C3
041C
03CF
0380
039C
03D4
03CE
03B3
03BB
03C3
03B8
03D5
041C
0410
0380
0323
0399
0410
02C7
FF42
FB4A
F92D
F94E
FA14
FA20
F9B1
F9A2
F9FC
FA30
FA18
FA02
FA09
FA03
F9F9
FA0E
FA1C
F9E2
F999
F9C8
FA55
FA63
F9AE
F992
FBC1
FFDF
036A
047E
03D0
0359
03D0
045D
0448
03DC
03A2
039F
039D
03AE
03DD
03D8
036B
0312
036A
040E
0406
0368
0363
042D
03F6
0117
FC98
F95D
F8E8
F9F7
FA86
FA29
F9CF
F9F4
FA13
F9D4
F9A6
F9DB
FA0B
F9E5
F9CE
FA20
FA6B
FA3A
F9FC
FA44
FAA4
FA47
F9A8
FA90
FDDD
01F8
0464
0476
03B9
03A3
03FE
03F7
03A1
038C
03AE
03A3
038A
03C3
0419
0402
0397
0381
03DA
03EF
036D
032C
03D1
0437
025C
FE39
FA5D
F912
F9D2
FA7F
FA30
F9BD
F9E5
FA49
FA4D
FA07
F9E2
F9DD
F9C5
F9C3
FA17
FA6E
FA41
F9DA
FA04
FA9E
FA87
F9A9
F9D7
FCA2
00F0
03F8
046E
039A
0348
03B4
03FA
03D2
03C8
040A
0414
03C2
03B2
041E
044B
03BF
032D
0351
03B3
037F
0312
0370
0441
0394
004F
FC01
F968
F963
FA57
FA94
FA23
F9E2
F9ED
F9DF
F9C8
F9EF
FA19
F9E8
F9A8
F9E7
FA6B
FA76
FA09
FA0F
FAD7
FB46
FA75
F9A0
FB14
FF0C
02ED
0459
03D3
036F
03E7
044A
0403
03AE
03DB
0418
03DB
037C
03A1
0414
0417
03B0
03A1
03F8
03D6
0319
02ED
03CB
0402
01A1
FD55
F9FD
F952
FA28
FA67
F9BB
F965
F9FB
FA9A
FA77
FA04
F9F7
FA2B
FA27
FA12
FA42
FA6F
FA34
F9EE
FA34
FAAC
FA73
F9CD
FA76
FD90
01CE
0492
04D3
03F9
03B9
041F
044A
0408
03D9
03E3
03D5
03AE
03BB
03F0
03ED
03AE
039F
03D9
03D9
036A
0342
03F3
0477
02E9
FF0B
FB12
F944
F98D
FA30
FA27
F9DA
F9DC
FA09
FA10
FA0D
FA2D
FA3D
FA07
F9E1
FA31
FAA5
FA8F
FA1E
FA31
FACE
FACD
F9D1
F98D
FBE7
0049
03F2
0500
043B
0399
03D9
0442
0434
03FC
03FD
0405
03E0
03D2
03FF
03FF
03A0
036D
03CC
0423
03C2
032A
0372
0456
03E4
00CE
FC69
F972
F90F
F9E1
FA39
FA04
FA11
FA6E
FA81
FA36
FA0A
FA20
FA26
FA0B
FA25
FA7D
FA9C
FA54
FA33
FA98
FAD7
FA32
F988
FADF
FEB7
02E7
04EC
04A5
03E9
03EB
0437
040F
03A9
039F
03DE
03E0
03A0
0398
03DB
03EE
03B0
0399
03D2
03D4
037A
0386
044C
0474
0248
FE1B
FA61
F91D
F9D7
FA9C
FA71
F9FB
FA03
FA5B
FA80
FA7C
FA8B
FA85
FA42
FA19
FA56
FAA2
FA91
FA6A
FAA5
FAEC
FA71
F986
F9F4
FCFF
016F
0488
04F9
0407
0388
03C3
03EA
03BA
03A7
03D6
03F1
03DC
03DD
03FC
03E6
0395
0382
03D5
03F1
0366
02F7
03A3
04AA
03D0
0035
FBE1
F98D
F9A2
FA63
FA7C
FA3C
FA54
FA96
FA80
FA38
FA42
FA7D
FA55
F9EA
FA03
FAAF
FAFA
FA7B
FA21
FAA4
FB32
FABF
FA23
FB79
FF41
0348
050F
0485
039E
03A5
0414
040B
03BD
03C1
03F9
03F8
03DD
03F8
040B
03C1
0375
03B4
042F
0408
034D
0323
03F4
042C
01E5
FD9D
FA1B
F941
FA15
FA8D
FA38
FA15
FA8B
FAE3
FA9E
FA2F
FA27
FA63
FA7C
FA7A
FA95
FAA4
FA69
FA3B
FA97
FB06
FA94
F9AA
FA53
FDB8
0226
04C2
04BB
03C9
03A9
0433
0454
03E4
03A8
03EF
042C
0406
03E3
0408
0406
039B
0350
0393
03E6
03C4
03AD
0447
04BF
033C
FF55
FB28
F940
F9D1
FAD9
FAD5
FA3C
FA1D
FA6E
FA81
FA4C
FA49
FA7A
FA7F
FA61
FA80
FAC8
FABB
FA54
FA30
FA84
FA93
F9E6
F9B4
FBD4
0028
0417
0552
0453
0355
0381
0424
0448
03FC
03D6
03FE
0425
041C
03F7
03C9
039C
039F
03EC
0422
03DD
038D
0404
04DD
0443
011A
FCC5
F9E2
F979
FA4C
FABC
FA88
FA61
FA85
FA90
FA60
FA54
FA86
FA8B
FA42
FA2C
FA87
FAC9
FA8C
FA47
FA7D
FAB5
FA48
F9E5
FB38
FEBF
02B3
04CB
04AF
03EE
03C9
03FD
03E8
03B9
03DF
041C
03FF
03C6
03F3
0453
0449
03DD
03BE
0417
0441
03E6
03BB
0449
046F
025A
FE28
FA6B
F958
FA55
FB2D
FAE0
FA43
FA3D
FA95
FAAC
FA7D
FA61
FA68
FA62
FA60
FA8D
FAB0
FA71
FA1C
FA52
FAD3
FAA1
F9D1
FA3A
FD4A
01C5
04D1
051A
0400
0381
03F4
0455
041B
03D1
03F1
042D
042B
0425
044F
0453
03FD
03C5
0408
044F
0411
03C1
041D
0497
037E
0021
FC20
F9D7
F9CB
FA79
FA93
FA54
FA6E
FAB1
FA90
FA3E
FA43
FA83
FA7F
FA43
FA50
FAA6
FAB3
FA5C
FA40
FAA9
FAD1
FA23
F9C8
FBAE
FFD3
03AE
0507
0464
03D5
0426
047D
0436
03D9
0409
0478
0487
0442
0429
0442
0429
03EE
040E
046A
044A
03BD
03D5
04C4
04C0
0200
FD68
F9ED
F94E
FA65
FAFF
FA83
FA00
FA2D
FA83
FA64
FA1A
FA25
FA5F
FA70
FA78
FAA8
FABA
FA7B
FA5B
FAB7
FAF0
FA48
F979
FA78
FE15
0289
051F
0527
0445
040C
0456
045E
0439
0463
04A5
047A
041F
0435
04A0
04A3
041D
03D0
0426
047A
0430
03E0
045D
04D0
0337
FF2F
FB13
F965
F9FD
FACA
FAA6
FA37
FA4F
FAA9
FAA8
FA5D
FA44
FA65
FA67
FA50
FA74
FAB4
FA92
FA31
FA4F
FAE9
FAF6
FA38
FA50
FCE0
0116
044B
0504
0453
0407
046F
049B
0435
03F3
043F
048D
0467
0435
0463
0491
0452
040B
0438
0475
042A
03C5
042B
04EC
0429
00DB
FC8D
F9E3
F9B0
FA6A
FA8E
FA4B
FA65
FAAA
FA83
FA2C
FA4B
FAB8
FAC1
FA60
FA42
FA9E
FAD5
FA93
FA72
FAE8
FB34
FA74
F9A0
FAF9
FF0C
036C
0561
04E5
040B
041B
0495
04B2
0495
04A9
04C5
0489
042B
0421
044E
042F
03DC
03F1
0465
0468
03E1
03E2
04CD
0503
02A7
FE4F
FAB8
F9B4
FA6B
FAEA
FA8E
FA2B
FA4D
FA7D
FA50
FA25
FA56
FA94
FA98
FABE
FB3C
FB74
FAE7
FA3C
FA62
FB05
FAF2
FA2E
FA90
FD85
01DB
04D0
0533
046E
0446
04BC
04D4
046F
0442
0482
04B0
048E
0466
045F
0437
03E6
03E0
044F
0497
0436
03CB
0442
04FD
03F9
0062
FC15
F9B1
F9B4
FA78
FA98
FA4B
FA52
FA9A
FA94
FA48
FA48
FAB1
FAF4
FAC0
FA87
FABD
FB1C
FB2B
FAF5
FABB
FA63
F9EC
FA2F
FC4F
001A
03B5
0547
04D6
0407
0420
04D0
0517
04B4
044B
0453
0489
047D
0434
0406
041B
0433
0408
03C0
03E1
0483
04C5
0361
001B
FC65
FA33
FA1A
FAE3
FB07
FA5B
F9E1
FA3C
FADF
FAF9
FA93
FA54
FA78
FA9A
FA78
FA6B
FAD7
FB6E
FB6D
FAA6
FA13
FB21
FE3B
0226
04E7
0576
048C
03CB
0411
04C0
04CD
042E
03CD
0426
04A1
048B
042D
0447
04C5
04C0
03EC
0354
0405
0547
04F3
01E0
FD67
FA20
F957
FA24
FADC
FAC4
FA55
FA46
FAAC
FB0E
FB0A
FAC2
FA99
FAAA
FABB
FAA4
FA9E
FAE5
FB2C
FAD8
FA07
FA15
FC68
0097
045D
05BB
04F2
03E9
03EB
048C
04C0
045F
041B
044F
0488
0452
03F8
040A
0471
0487
0412
03B5
041F
0502
0507
0305
FF44
FB7F
F983
F9A9
FABA
FB48
FB06
FAAD
FAD0
FB1E
FB02
FA96
FA81
FAF4
FB4C
FB04
FA86
FA90
FB06
FAFF
FA32
F9D0
FB73
FF2E
032D
0564
0570
0497
042E
0462
048B
0449
03F4
0408
0477
04B9
047F
0419
0402
0437
0443
0409
040F
04BC
055D
046C
013B
FD0D
FA2C
F9BE
FAC6
FB73
FB12
FA69
FA5B
FACE
FB0B
FAD3
FA94
FAA4
FAC9
FAB5
FA9B
FAEF
FB92
FBBD
FAF8
FA01
FA63
FCFA
00EC
0440
0587
04F8
0403
03D1
0457
04C6
04A9
0458
0457
049D
04B2
0476
044D
0478
0497
043A
03B4
03DA
04B8
04EF
0303
FF31
FB90
FA0A
FA80
FB42
FB17
FA5E
FA1E
FA8B
FAF4
FADE
FAA6
FAD7
FB44
FB47
FAC2
FA6D
FADD
FB96
FB86
FA7E
F9DC
FB53
FF01
0304
052F
0515
042C
0404
04B2
0532
04EE
046A
0460
04B2
04B0
0433
03E0
0430
04A6
0486
03F5
03F0
04D9
0590
0466
0104
FD01
FA7A
FA23
FAEA
FB52
FAE8
FA55
FA55
FADC
FB49
FB40
FB01
FAF8
FB1E
FB20
FAF1
FAEA
FB28
FB2B
FA7F
F9C1
FA74
FD6C
0191
04A3
055C
0487
03E1
0431
04D0
04E4
0477
042B
043F
0452
0411
03BC
03C3
041D
0451
0430
0426
049E
052F
04A8
0232
FE60
FAFE
F995
FA13
FB05
FB25
FA86
FA26
FA88
FB1A
FB1F
FAB2
FA94
FB07
FB66
FB1E
FA8F
FA8A
FB0D
FB31
FA92
FA55
FC15
FFE1
03C3
05A2
054E
045C
0433
04B8
04F7
0494
0421
0433
0495
04B0
046A
043E
0480
04DD
04D4
0472
0455
04C6
0502
03BD
008E
FCB7
FA34
F9E8
FADA
FB63
FAEC
FA4B
FA6E
FB20
FB6F
FB09
FA97
FAB6
FB1F
FB30
FAF6
FB18
FBAD
FBE0
FB19
FA38
FB01
FE28
0240
050D
059D
04E2
045C
048D
04E9
04D5
0477
0462
04C8
0536
052A
04B6
0462
0470
0483
042E
03BC
03EC
04B1
04A4
0252
FE2D
FA8E
F96B
FA53
FB32
FAD9
FA15
FA28
FAEE
FB2C
FA6F
F9B4
F9F8
FAD0
FB15
FA98
FA54
FAEB
FB9A
FB3C
FA14
F9E4
FC19
001D
03CE
0580
0551
049B
046C
04C2
0502
04ED
04D6
0506
053E
050D
0489
0447
0485
04BD
045D
03BF
03DD
04EB
0594
042F
00A8
FCD7
FAB0
FA7D
FB05
FB23
FAC8
FA7C
FA79
FA86
FA77
FA73
FAA5
FAEA
FAFB
FAD4
FAC3
FB08
FB72
FB7D
FAEE
FA68
FB2D
FDF2
01CF
04BC
056C
048C
03E4
0456
0522
0533
04A6
0478
04F8
054F
04D0
040D
040C
04C6
0526
04A6
0423
049F
058E
0516
0230
FE0E
FAFE
FA28
FABD
FB3E
FB10
FAB0
FAB2
FAFC
FB0C
FABC
FA7B
FAB2
FB26
FB41
FAE3
FA9A
FAE3
FB57
FB1C
FA45
FA4A
FC96
00AB
0443
0593
0502
0452
0479
04E7
04D3
0470
0478
04EE
0512
0491
041B
046C
052E
0563
04C6
0434
048A
0569
055D
0348
FF95
FBF8
FA0A
FA0D
FAEA
FB62
FB28
FAE6
FB22
FB85
FB60
FAC4
FA81
FAF4
FB72
FB3D
FAA6
FAA1
FB40
FB6E
FA8D
F9D1
FB3C
FF22
036B
05AD
058D
04B1
048C
04FE
0516
0493
0423
0459
04EB
0524
04D4
0482
04A3
04FD
04FD
048F
0455
04D4
056D
049C
0193
FD79
FA97
FA1A
FB02
FB84
FB1A
FAB0
FB09
FBA7
FB9C
FAF6
FAA0
FB00
FB61
FB14
FA82
FA94
FB42
FB7C
FAAE
F9D0
FA9A
FDA6
01AE
04AC
0598
0504
043F
0417
0467
049A
0476
044D
0473
04BA
04B4
0469
045F
04D2
0530
04E1
0442
0453
052F
055E
0345
FF36
FB76
FA00
FA94
FB5F
FB2E
FA7A
FA4D
FAD0
FB45
FB31
FAF0
FB0C
FB65
FB62
FAD9
FA62
FA95
FB34
FB65
FADB
FA89
FBDD
FF2B
02FD
0549
055C
046B
0420
04D8
058C
0556
0493
0448
04B4
0513
04C4
0436
0441
04E6
0546
04E9
047F
04D6
055F
046F
0136
FD16
FA6E
FA36
FB2F
FB8D
FAF0
FA62
FAAD
FB56
FB76
FAFE
FAB7
FB11
FB88
FB62
FABA
FA63
FAC3
FB3D
FB04
FA66
FADB
FD77
0175
04B0
05A7
04E5
0438
049B
0551
0534
045D
03F6
0483
0526
04E4
0417
03E8
049C
052B
04C9
0428
047C
057F
0559
02C9
FECD
FBA8
FA87
FAAF
FAD6
FA9E
FA80
FAC6
FB1A
FB12
FACB
FAB8
FB05
FB60
FB68
FB23
FAFC
FB3E
FB98
FB64
FA96
FA54
FC08
FFB0
0374
055D
053C
0491
049D
0521
0530
04B2
0479
04EB
0562
0524
0482
0465
04FA
0572
0524
047B
0477
0554
05EE
04BA
015D
FD4B
FAA2
FA55
FB69
FC13
FB93
FAC2
FABF
FB6B
FBB1
FB2A
FAAD
FB06
FBBC
FBC5
FB1E
FAD2
FB57
FBB4
FAEA
F9C8
FA73
FDD8
024E
052D
0578
0473
03DC
0438
04DC
0514
04DC
04A0
049E
04B6
04AE
0485
046D
0483
04A7
04AA
04AD
0505
0582
050D
029D
FEB5
FB64
FA57
FB21
FBE2
FB82
FAB0
FA95
FB2D
FB79
FB0E
FAA4
FAF5
FBA1
FBBD
FB28
FAA8
FAC0
FAFD
FAB6
FA2E
FA93
FCC9
0053
0395
0532
0526
0491
0482
0503
054F
04F7
0476
0484
04FA
0500
044A
03AD
0400
04E0
0525
048E
042F
04D5
0586
0452
00B9
FC99
FA52
FA60
FB47
FB89
FB14
FABB
FAE0
FB1D
FB03
FAC5
FADC
FB57
FBBA
FBA4
FB47
FB27
FB60
FB6D
FADE
FA48
FB1F
FE3A
0280
058C
05ED
0490
039E
041B
051F
0556
04B9
044C
0490
04E9
04B1
043F
044F
04CF
04F1
0477
0435
04E4
05C4
0514
020B
FDFC
FB27
FA94
FB57
FBDD
FB8B
FAF9
FADD
FB2C
FB58
FB23
FAEB
FB15
FB79
FB97
FB4D
FB01
FB0B
FB23
FACD
FA4C
FACB
FD38
00FD
043E
0590
053A
049B
0493
04D3
04BC
0465
046F
0501
0574
052F
047C
042F
0493
0516
051C
04DA
050D
05C6
05E6
041C
0071
FC95
FA70
FA6D
FB4F
FBA7
FB3F
FAE7
FB20
FB78
FB4C
FAD0
FAC7
FB5C
FBC9
FB72
FAD2
FAD4
FB5C
FB4C
FA3C
F994
FB33
FF12
02F4
04BF
0499
043F
04AD
053D
0511
0481
048A
053D
059E
0515
0451
0446
04CA
04F0
0489
0487
0570
0615
049C
00C8
FCA6
FA8E
FAD1
FBC3
FBDD
FB38
FAD9
FB1F
FB71
FB4D
FAF7
FAF1
FB2E
FB44
FB31
FB5E
FBCD
FBCC
FB04
FA7A
FBD1
FF53
033B
055D
054E
047D
044F
04BF
0500
04E2
04EB
0544
0560
04F0
048D
04E0
0580
0566
0480
0407
04C6
0592
0455
00A4
FC8A
FA70
FAA1
FB7D
FBAA
FB5C
FB53
FB85
FB58
FAD3
FAB1
FB36
FBA6
FB57
FAC5
FAEA
FBB5
FBF3
FB1D
FA85
FC13
FFDF
03C6
05A1
0559
048E
046E
04B1
049A
0440
0451
04E8
0556
0527
04C8
04D0
0515
04F6
0479
0468
050C
0543
038D
FFF5
FC5E
FA9D
FAB6
FB3D
FB3C
FB07
FB3D
FBAB
FBA4
FB22
FAD4
FB0F
FB52
FB1C
FAD0
FB15
FBA7
FB8B
FAAD
FA9B
FCE6
0107
0488
0590
04B1
03E4
042D
04E3
0515
04CA
0495
048D
045D
041D
045D
0525
0598
0518
0453
047A
0563
0545
02BB
FEA9
FB7F
FAA7
FB4C
FBB5
FB49
FAC4
FACB
FB17
FB29
FB27
FB80
FC0B
FC15
FB74
FAE0
FAFB
FB5B
FB23
FA84
FAF8
FD99
018C
04A4
058C
04F2
0463
048B
04E6
04EB
04CE
04F4
052E
050B
04AC
04AE
0528
0561
04DF
0450
04B5
05A7
0548
025C
FE18
FB22
FAC4
FBC5
FC25
FB6B
FAAD
FABC
FB22
FB1D
FACE
FAD6
FB34
FB3E
FACF
FAA2
FB29
FBA3
FB21
FA3C
FAE4
FE1D
0270
054A
059F
04AF
043A
0491
04E4
04C9
04B0
04F7
053A
0507
04AF
04D9
0571
05A6
051F
04A0
04FE
05AA
04FB
021C
FE3A
FB75
FAC8
FB59
FBC6
FB9D
FB5F
FB6A
FB80
FB4C
FAF8
FADC
FAE9
FACC
FA8F
FA9F
FB0E
FB40
FAC1
FA53
FB76
FEA4
026B
04B6
04EA
044B
0439
04B2
04D3
0462
041E
048D
0535
055F
0529
053D
05A2
05A8
0521
04E9
0595
0614
0495
00DD
FD02
FB47
FBAB
FC4B
FBE2
FB19
FB1F
FBD5
FC1F
FB9B
FB17
FB3B
FB8A
FB48
FAC0
FAD6
FB84
FB99
FA8D
F9CA
FB5A
FF5A
0380
0573
051D
0448
044D
04D5
04EB
047E
0453
04C4
0547
0552
0521
0535
056E
0541
04BF
04C5
05AC
063B
04A1
00AD
FC83
FA92
FB12
FC12
FBE6
FAEE
FA97
FB45
FBEB
FBA8
FAF1
FABC
FB12
FB2A
FAC8
FA8F
FAD5
FAE4
FA30
F9C1
FB6D
FF74
03AA
05A0
0533
0451
046A
04FE
04F0
0455
0431
04CA
0548
050B
049A
04B8
052A
0529
04D1
0527
0656
06BC
048A
0023
FC0E
FA66
FADE
FB9D
FB8B
FB20
FB31
FBAA
FBD7
FB7A
FAFE
FAC1
FAB6
FACD
FB2F
FBCF
FC03
FB33
F9FA
FA06
FC82
0099
040C
054F
04DD
0452
0490
051D
0536
04E4
04BF
04FF
0540
053F
053C
0569
0560
04C4
0429
049C
05FE
0677
043F
FFDD
FBF1
FA85
FB1F
FBC9
FB88
FB07
FB11
FB57
FB2A
FAC0
FAD2
FB56
FB71
FADE
FA8A
FB31
FC01
FB8F
FA2C
FA1C
FCF7
016B
0486
04F5
0421
0400
04C0
0531
04DC
04A2
0537
05FF
05FC
0551
04FD
0541
0549
0498
0415
04D3
062B
05ED
02DA
FE59
FB31
FAB2
FBB1
FC43
FBD1
FB24
FAE7
FAE4
FAB4
FA8E
FADC
FB64
FB74
FAF0
FA99
FAF7
FB67
FAF5
FA0E
FA8B
FD9D
0204
0516
057A
046A
03F8
04B0
057C
0586
0545
057C
05EF
05D4
0526
04C2
0510
0564
051E
04CE
0560
064B
0598
023E
FDCC
FB00
FAE4
FBFD
FC60
FBC3
FB1D
FAE9
FAB4
FA3B
FA0F
FAAA
FB78
FB8D
FB01
FAC3
FB20
FB30
FA5C
F9C2
FB4A
FF33
035B
055D
0502
0412
040C
04C2
053B
053C
0547
0591
05AB
055A
051A
055E
05BD
057B
04C9
04C7
05DD
06A1
0518
0110
FCB3
FA67
FA81
FB64
FB9E
FB44
FB24
FB58
FB4A
FAD6
FA9C
FAFD
FB65
FB1C
FA76
FA72
FB2F
FB85
FAB5
F9FB
FB75
FF75
03AB
0589
0505
0449
04DC
0603
0635
0558
04AC
04E4
0544
0503
0493
04E1
05B7
05F2
054C
04F2
05B4
0645
0472
000E
FBB7
FA1D
FB1D
FC42
FBDB
FAA6
FA42
FAF1
FB92
FB6E
FB02
FAF2
FB08
FACA
FA80
FADB
FBA1
FBB1
FAB5
FA2F
FC0E
003B
044F
05F5
0542
043D
0472
0588
063D
060F
0583
052B
0506
04E9
04EE
0534
056E
0534
04C4
04D5
0577
0572
035F
FF6B
FB94
F9D6
FA53
FB7A
FBD6
FB58
FAD1
FAB3
FABF
FAB0
FA9B
FA99
FA85
FA63
FA9F
FB72
FC35
FBF5
FAF6
FB05
FD98
01D3
0515
05B9
04B5
042D
04E7
05DE
0605
05AA
05A7
05FE
05FE
0586
0545
0584
058C
04D5
0425
04A7
05E2
05A9
0293
FDF6
FAAA
FA0E
FAE7
FB51
FAEF
FAA3
FAD1
FAD9
FA50
F9CC
F9FA
FA80
FA8C
FA2E
FA6B
FB98
FC78
FBBC
FA26
FA44
FD9E
02B0
0648
06C2
056B
04AD
0566
067B
06AC
0610
0592
05A3
05EC
061E
0655
068F
065A
0585
04C8
050C
05DA
0547
0210
FD74
FA3E
F9D7
FAEE
FB56
FA96
F9F0
FA40
FAD4
FAAE
FA0E
F9F1
FA67
FA74
F9C5
F971
FA61
FBAE
FBAD
FA85
FA9A
FDC2
02BF
065B
06E5
05B0
0501
0578
0608
05EF
0599
0597
05BA
059E
0592
061E
06F9
0720
0647
0570
0589
05D6
047D
00D9
FC95
FA16
FA0B
FB02
FB47
FAAD
FA40
FAA1
FB41
FB46
FAA9
FA21
FA22
FA62
FA73
FA5B
FA5E
FA75
FA65
FA86
FBE1
FF0D
0319
0617
06EB
0646
05A4
059F
05AF
0551
04D4
04D2
0547
05B1
05D7
05F1
0607
05CE
0558
0554
0609
0656
0494
009C
FC6A
FA36
FA3B
FAE1
FADE
FA77
FA8D
FB22
FB7B
FB43
FADF
FAA4
FA68
FA23
FA5A
FB4F
FC2B
FBBA
FA36
F9A8
FBDA
0037
043D
060B
05FE
05AB
05DD
0615
05B8
0509
04BC
04F9
054D
0567
0579
05AD
05B9
054D
04C8
04F0
05C1
05EA
03ED
FFE7
FBD2
F9C0
F9E1
FAB0
FAD2
FA6C
FA64
FAEE
FB5A
FB30
FAE0
FAFD
FB59
FB57
FB02
FB01
FB7A
FBA0
FB00
FAB1
FC66
004D
046D
0696
068D
05DE
05D0
063C
0664
062F
0605
05FC
05BF
053B
04C8
0487
0438
03E6
043D
0599
06E5
062E
02C1
FE45
FB36
FA80
FAF3
FB09
FA81
FA14
FA20
FA37
F9F2
F9A4
F9E3
FAB2
FB77
FBCA
FBDB
FBF3
FBEB
FB7E
FB13
FBBF
FE33
01B5
0493
05B7
059E
058B
0600
066C
0644
05DA
05CE
0607
05DC
0537
04DA
0541
05BD
0570
04C5
04E5
0565
039E
FD6D
F45D
ED03
EAA8
EC39
EDF6
EDA2
EC36
EBAB
EC55
ED0C
ED22
ED16
ED6F
EDD6
EDC3
ED67
ED68
EDDB
EE25
EDF5
EDD7
EE79
EFAF
F099
F0A8
F021
EFA1
EF6F
EF75
EF9A
EFE8
F056
F0A4
F091
F030
EFE9
F005
F04E
F047
EFD3
EF81
EFE9
F0B1
F092
EEE9
ED2B
EE29
F351
FAD8
010B
0384
02EC
01B2
017D
021F
0294
0260
01D3
016B
015C
0185
01A3
0193
0190
01F7
02BA
034B
0366
03A6
04EB
06FF
086F
081C
06B6
05FA
0699
077B
0766
0699
0641
06CA
0779
0796
0750
0728
071E
06E6
0698
0678
064B
058E
0479
03DF
037F
0156
FBBC
F403
EE00
EC61
EE0F
EFB3
EF6F
EE45
EDFE
EEA7
EEE5
EE19
ED41
ED9E
EF17
F067
F08F
EFDC
EF72
EFFD
F106
F197
F15C
F0F9
F129
F1D2
F22A
F1C8
F135
F132
F1BF
F236
F255
F272
F2B0
F2A2
F20F
F184
F185
F196
F0F4
F00C
F040
F1B3
F258
F084
EE1E
EF73
F63B
FEDE
03F0
03E3
01F4
01AB
02F9
037C
025D
015D
0210
03B4
0471
03E2
033E
0372
0424
04BD
056B
06A1
0812
08DD
08AB
081E
0807
0884
091F
0978
0990
097F
0949
08F2
0892
084F
0843
0859
0840
07C3
073D
074C
07C7
075F
0515
020D
010E
0331
0598
03B9
FC69
F3AE
EEB3
EE9D
F041
F07D
EF7B
EF40
F053
F130
F0BC
EFD6
EFDD
F0BE
F14F
F119
F0D0
F11C
F1C7
F23C
F250
F239
F21B
F202
F215
F266
F2A6
F284
F24D
F29F
F365
F3B7
F31C
F243
F210
F26B
F2A6
F29E
F2B6
F2DE
F28A
F1E1
F201
F337
F3CE
F224
EFF0
F186
F8C8
01FD
0748
06CC
0406
031A
045E
0559
04CB
040B
047A
0564
054D
045C
042C
059C
07CC
094B
0991
091D
08B6
08C9
0930
0964
090A
0869
083B
08CC
0988
09C0
099C
09C7
0A3C
0A3E
09B3
0983
0A23
0A7D
0946
06E8
050E
0463
03F5
0333
0341
0503
066F
03D8
FC81
F472
F076
F109
F289
F203
F040
EFB3
F0E2
F204
F1B2
F09D
F050
F12E
F259
F2FC
F2FB
F2A5
F262
F29C
F35A
F401
F3E9
F33D
F2E7
F370
F44F
F49B
F42B
F3A3
F385
F3BC
F40F
F474
F4BA
F472
F39F
F2F4
F2F2
F328
F2F3
F2AA
F328
F41B
F3E4
F20F
F119
F454
FBB8
031D
0674
05D7
049A
0502
0641
0691
05C7
0517
052E
05BB
06A8
085E
0A97
0BFD
0BBC
0AAE
0A32
0A68
0A74
0A25
0A3B
0AF6
0B70
0AEE
0A2F
0A68
0B58
0B7C
0A54
094B
09BE
0B08
0B58
09EC
07A3
05B8
04CD
04F7
05BF
060D
0500
0369
037A
05CD
074F
03E1
FB79
F31C
EFC1
F13B
F370
F392
F273
F202
F263
F290
F282
F32C
F484
F527
F45E
F355
F36F
F45F
F4D6
F491
F471
F4DD
F529
F4C7
F43B
F44F
F4E8
F538
F4E9
F473
F453
F467
F464
F448
F41B
F3B3
F32B
F2FC
F344
F371
F32F
F326
F3E9
F493
F3A4
F198
F193
F64C
FE75
057C
0821
076A
0687
06DE
0754
06F3
06A4
07C9
0A1C
0BE3
0C0A
0B4A
0B12
0BD6
0CE0
0D57
0D0F
0C5D
0BB7
0B72
0B9E
0BF4
0C0B
0BBA
0B36
0ADD
0AE3
0B2B
0B50
0ACE
0970
07B5
0690
0674
06BA
0665
0584
052E
05DC
0677
05BB
0450
044E
0615
06B3
02BF
FAC2
F36D
F0D2
F259
F448
F468
F3D5
F44F
F578
F5B9
F4E8
F476
F50E
F596
F515
F463
F4E1
F653
F72F
F6C8
F600
F5BC
F5B3
F535
F47A
F447
F4AF
F506
F515
F55B
F5E3
F5CE
F4AD
F361
F2F4
F335
F351
F32E
F355
F3C2
F3E9
F3DB
F447
F4F8
F47C
F2A6
F282
F79E
0100
08DE
0AA2
07E5
05F1
076D
0A56
0BD8
0BDF
0C10
0CDF
0D5D
0D52
0DA8
0E86
0EA6
0D62
0C10
0C30
0D24
0D28
0BEA
0ACD
0ACB
0B57
0BA2
0BCB
0C2A
0C23
0AC5
0857
064D
057D
0566
0579
05FB
06F8
077C
06DC
05F5
05FA
068C
0661
05A7
0618
07F0
0838
03C7
FBB5
F4FA
F319
F4A8
F5EF
F596
F522
F5B9
F677
F649
F5BD
F5FC
F6D1
F6E9
F5E9
F505
F541
F612
F659
F5F0
F57D
F540
F4FE
F4CE
F511
F5A3
F5C8
F534
F48A
F479
F4CC
F4D6
F481
F441
F424
F3D4
F395
F42A
F55D
F5BB
F4A5
F3B6
F4BA
F6C9
F71B
F54B
F506
F9F5
02A6
0988
0B3F
0A0A
0A11
0C1A
0DAB
0D63
0CC9
0D7F
0EB3
0E8B
0D1D
0C53
0D13
0E08
0DBC
0C99
0BF2
0C07
0C24
0C16
0C5A
0CF9
0D33
0C78
0B02
095A
07D7
06C4
0687
070C
0783
0746
06E0
0744
081B
0810
06FD
0665
070F
0798
06B9
05DE
0758
0A1D
0985
02AB
F8D7
F2A6
F2EC
F639
F7C6
F6DC
F611
F6BF
F785
F700
F5E2
F5A8
F66C
F701
F6C2
F63B
F61D
F64E
F65C
F642
F642
F66D
F6BB
F72F
F783
F710
F5A7
F41D
F375
F3B6
F424
F46C
F4EF
F5BB
F60C
F55B
F46C
F472
F558
F5CE
F562
F54E
F66D
F75E
F633
F3F1
F4BC
FB70
05BC
0DDC
1045
0EA3
0D10
0D63
0E42
0E13
0D48
0D3A
0DFB
0E60
0DE8
0D70
0DBF
0E3E
0DDD
0CB9
0C1C
0CD8
0E3A
0EC6
0DAC
0B57
08E6
0755
0708
07A4
0856
088A
0873
0892
08DD
08C4
082F
07B8
07C0
07E5
07CB
07CC
0831
0855
0778
0664
06E9
08F2
0941
04B2
FC95
F617
F4B9
F6D0
F84A
F7A5
F68A
F66F
F6B5
F66C
F62E
F6EF
F7F0
F772
F570
F41C
F50D
F733
F862
F807
F72B
F68F
F607
F576
F531
F53F
F50B
F45F
F3FF
F4C1
F641
F73C
F713
F65B
F5CF
F581
F55E
F59C
F62D
F680
F670
F6B1
F780
F7AF
F652
F531
F7F0
FFDF
098B
0FB5
1091
0EE0
0DF1
0E19
0DDC
0D05
0CD7
0DB5
0E5B
0DD6
0CFC
0D1C
0E04
0E5F
0DC8
0D42
0D70
0D58
0BCA
0950
07AE
07A8
0839
082A
07A2
07A1
0875
0959
0995
0959
093E
0960
0959
08F3
0875
0855
08B9
0935
0918
0851
080A
09C9
0D43
0F57
0C67
0440
FB2A
F612
F5D2
F721
F706
F5F5
F5F6
F71F
F78A
F659
F514
F578
F703
F7C7
F716
F626
F606
F644
F61B
F5C9
F5E3
F610
F591
F4B8
F4B4
F5E6
F737
F765
F678
F58E
F582
F62F
F6DF
F6FD
F679
F5E3
F625
F76C
F87F
F818
F6F6
F729
F8DB
F96E
F731
F4F0
F79D
0054
0A56
0FF5
105B
0F1C
0EF0
0F0B
0DF5
0C8F
0CA3
0DDB
0E2B
0CF3
0BE2
0C89
0E42
0F09
0DC8
0B3F
0910
085A
0915
0A43
0AAE
09F3
0900
08F8
09A3
09B3
08C4
07FE
084E
091B
0985
09EB
0AFD
0BFC
0B67
0970
0844
0944
0B0C
0B76
0AEF
0BF3
0ED5
0FED
0B6D
023C
F979
F553
F587
F6E8
F728
F695
F6A7
F7B0
F867
F7AC
F63D
F5FB
F785
F926
F8AB
F61E
F3ED
F40D
F5A9
F681
F613
F5FB
F71D
F81C
F786
F629
F5DC
F6BE
F72F
F64C
F527
F516
F5EE
F69B
F6CF
F713
F76A
F724
F64B
F60B
F701
F821
F830
F780
F749
F7E9
F8C0
F950
F994
F95D
F86E
F74F
F721
F816
F8DE
F86D
F7B1
F843
F994
F94F
F74A
F73A
FCAF
0614
0D93
0F1A
0C35
0979
0961
0AA6
0B01
0A21
0972
09CB
0A79
0A6F
09A3
08FF
0941
0A3B
0B00
0AE7
0A3D
09DE
0A11
0A45
0A04
09AD
09E4
0AC3
0BF3
0D48
0EB8
0FDA
0FFC
0F03
0DE1
0DB7
0E9E
0F93
0FAE
0F05
0E41
0DC7
0D96
0DA2
0DDB
0E1D
0E4D
0E69
0E51
0DD1
0D11
0C83
0C28
0B5C
09CB
0852
0826
0913
0974
0874
078E
08AE
0AEC
0A97
0555
FD44
F705
F501
F5B4
F659
F60E
F5DC
F68A
F770
F780
F6C3
F641
F69C
F75A
F7A5
F76A
F75C
F7F6
F8C1
F8D1
F7E4
F6C2
F653
F685
F6A6
F696
F6F7
F7FB
F8D4
F8C2
F81E
F7C6
F7F1
F829
F836
F855
F891
F87B
F7E9
F778
F7AB
F7EA
F74A
F62E
F610
F75E
F8A7
F88C
F78E
F70F
F749
F762
F707
F6C7
F6DF
F6CE
F68E
F719
F8AD
F983
F7EF
F5D6
F7E3
0013
0A62
1097
10BC
0E5E
0DAA
0F0A
102C
0FD1
0F20
0F7E
1089
10E8
1048
0F9A
0F7C
0F6F
0ECE
0DE7
0D9F
0E33
0EB7
0E05
0C13
0A37
09C3
0A92
0B47
0AF6
0A04
0951
0923
093B
096C
09A5
09A6
0938
08A6
0895
0937
09FD
0A4C
0A30
0A04
09B8
0929
0900
0A30
0C63
0E07
0E54
0E33
0E97
0F04
0EAD
0E22
0E76
0F2C
0EA5
0CFC
0CB4
0F15
10F4
0D75
0447
FADC
F678
F6D3
F800
F7EF
F7BE
F863
F8B2
F76D
F583
F4E6
F5D2
F6A6
F653
F59D
F59E
F63E
F6D3
F751
F7DF
F809
F75C
F65A
F5D3
F5C1
F5A3
F59A
F639
F755
F7EA
F77D
F6E2
F725
F80D
F878
F807
F79C
F7E1
F851
F835
F7C4
F797
F7B1
F7D1
F824
F8DD
F98C
F995
F914
F8B0
F8BE
F909
F95D
F9AD
F9B1
F907
F811
F7F5
F8E5
F92F
F790
F63A
F95A
0199
0A11
0D5C
0B8A
093A
098C
0B13
0B21
09D2
0955
0A4D
0B15
0A98
09E2
0A04
0A35
0965
0889
0986
0C48
0E9B
0F04
0E68
0E7A
0F7F
105B
1051
0FC7
0F61
0F2C
0EF9
0EE0
0EF9
0EF6
0EA6
0E68
0E98
0EE7
0EE3
0ECB
0F22
0F95
0F0E
0D1C
0ABF
0964
0954
0997
0963
0918
097C
0A59
0A95
09AD
088A
086D
094A
09CC
091F
083C
08C9
0A8C
0AB8
06AB
FF2B
F815
F493
F468
F542
F5CF
F68A
F7E7
F919
F91F
F83D
F794
F791
F79A
F757
F748
F7C3
F82F
F7F1
F78C
F7F3
F907
F9A5
F93A
F88A
F88C
F90B
F900
F806
F6DF
F666
F691
F6C4
F6C3
F6C0
F6D7
F6E2
F6E6
F715
F762
F76F
F712
F6B0
F6CD
F75B
F7BC
F785
F6FF
F6BF
F6DE
F700
F71A
F7B7
F918
FA68
FA91
F9C2
F965
FA34
FAEA
F9EE
F82E
F933
FF5E
0897
0FD5
1215
10E3
0FAE
0FC5
0FF1
0F1D
0E04
0DED
0EE3
0FD1
0FDC
0EFD
0D76
0B88
09D0
0920
098B
0A1E
0A03
0995
09BE
0A99
0B50
0B39
0A85
09D2
0984
09A8
0A23
0AB8
0B09
0AD6
0A51
09F1
09FC
0A6A
0B43
0C96
0E0C
0EEA
0EE7
0E85
0E57
0E3B
0DCA
0D36
0D27
0DD3
0E9F
0ECB
0E45
0DB2
0DBE
0E68
0F02
0ED9
0DFF
0D73
0E08
0EB9
0CAB
060F
FD01
F650
F4B6
F644
F73D
F680
F5E4
F6B7
F7BD
F747
F5EC
F5B4
F70F
F833
F7C1
F697
F633
F696
F6D1
F6D7
F75A
F82F
F847
F763
F6B8
F758
F8A5
F92D
F8A0
F7FF
F7F7
F80F
F7DA
F7D7
F86D
F8E3
F852
F729
F6A7
F71A
F78B
F751
F70C
F795
F8A6
F943
F921
F8DE
F8CA
F86B
F7A1
F752
F81B
F900
F880
F6E1
F63F
F7D1
F9F8
FA03
F7CC
F6A9
FA10
0196
08F6
0C42
0B8B
09FE
09FB
0AEC
0AFA
09FC
09B6
0B68
0E0D
0FAA
0FC1
0F84
0FD0
1017
0FA1
0EE9
0EDB
0F56
0F56
0E94
0E0B
0E91
0F9E
0FFE
0F68
0EB4
0EA2
0F1E
0FC4
1052
1040
0ECA
0C10
098D
08B0
0944
09F5
0A18
0A2F
0A9F
0AD6
0A3A
094E
090E
0977
099D
0942
0934
09BF
09E2
08F5
0820
08DB
0A83
0AEA
0999
0902
0B68
0F32
0FD0
0A97
01D4
FA60
F6F9
F6A9
F71F
F74D
F78E
F83A
F8E0
F8CD
F7FF
F738
F723
F77B
F772
F6DB
F686
F72D
F857
F8B2
F7AE
F63E
F5B2
F615
F656
F5ED
F58A
F5E9
F6B2
F714
F6F1
F6CA
F6F1
F747
F7A1
F7DC
F7AF
F6FA
F63F
F641
F6F3
F746
F693
F5D1
F67B
F865
F9BF
F97C
F893
F855
F8AA
F8D0
F8EB
F97B
F9E9
F912
F77A
F753
F974
FB69
FA58
F777
F7AC
FDE1
0744
0E66
10E1
107A
0F9B
0EB3
0D45
0BC6
0B31
0B78
0B8A
0ADE
0A1A
09EB
0A01
09BF
0955
096C
0A15
0ABA
0AF7
0AF1
0AEF
0B15
0B6F
0BC9
0BA3
0AAF
096D
08F3
09F2
0BF9
0DDE
0ECB
0EE8
0EF4
0F60
0FEB
0FFE
0F51
0E4B
0DC2
0E0B
0E7F
0E4B
0DB6
0DC2
0E8D
0EEE
0E20
0D0B
0D0B
0DFB
0E6D
0DA3
0C66
0B91
0ACE
09A5
08F7
09E0
0B18
0943
02E1
FAE6
F5F8
F5A2
F75E
F80E
F71E
F604
F5D4
F64C
F6C7
F71A
F74D
F734
F6C7
F686
F6F1
F7CB
F857
F831
F79B
F70A
F6D2
F716
F7B9
F862
F8BD
F8AD
F836
F778
F6D9
F6D6
F76F
F80A
F810
F7A0
F749
F751
F778
F788
F7B6
F81D
F843
F7C5
F73C
F7A1
F8BE
F93D
F88B
F7B4
F7B5
F80F
F7D3
F754
F799
F873
F889
F791
F710
F807
F8E3
F789
F542
F679
FD94
077C
0EAA
10C4
0FEB
0F2D
0F78
1005
1037
1017
0FBF
0F2D
0EAE
0EB1
0F12
0F27
0EB5
0E68
0ED3
0F91
0FE5
0FD0
0FDA
101B
1015
0F58
0DED
0C3F
0AE9
0A4F
0A31
09EC
0960
0931
09DD
0AE5
0B54
0AF5
0A83
0A84
0A8E
0A1F
09B9
0A23
0AE4
0AAE
0977
08B8
0925
09A0
094B
0949
0B01
0DBF
0F7A
0FAD
0FA9
1008
0F99
0DDA
0CE1
0E82
1039
0CE6
0388
F9AB
F565
F6A4
F897
F843
F70E
F71E
F7FF
F807
F736
F6E3
F74E
F73F
F644
F599
F613
F699
F5E4
F4A2
F46C
F552
F5E9
F58B
F51E
F582
F65F
F6D3
F6B8
F6B6
F73F
F7F8
F820
F782
F6B2
F67D
F727
F825
F890
F820
F7AE
F83A
F973
F9FF
F95A
F893
F8B4
F96E
F9E2
F9E5
F9BA
F947
F878
F7E3
F82A
F8E3
F8FF
F873
F85D
F911
F917
F785
F6B2
FA42
0214
095D
0BF3
0AD5
09EA
0AB9
0B8C
0B0B
0A3A
0A5D
0AC6
0A24
08EA
08CC
0A0D
0AF6
0A6D
0974
0941
095D
08FB
08E9
0A88
0D62
0F80
0FF3
0FB9
0FD7
0FD6
0ED8
0D58
0CE2
0E0C
0FB0
106C
1030
0FC8
0F91
0F5D
0F3F
0F7D
0FF5
1033
1013
0FDA
0FC5
0FC6
0F87
0E87
0C99
0A66
0912
091E
09F2
0AB4
0B26
0B5F
0B18
0A05
08E3
0908
0A1E
0931
03B0
FB54
F52F
F428
F60B
F6F2
F619
F59F
F696
F788
F720
F643
F694
F7DB
F878
F7F8
F7AB
F867
F938
F905
F848
F809
F81D
F7B7
F70F
F720
F808
F8E2
F933
F983
FA23
FA50
F935
F764
F674
F711
F832
F88A
F803
F75D
F708
F701
F750
F7D4
F801
F77A
F6B2
F65D
F687
F6B4
F6B1
F6B7
F6E4
F702
F6FB
F71D
F7A5
F842
F881
F883
F8B4
F8DC
F851
F745
F6FD
F81E
F99C
FA19
F9AD
F983
F9FD
FA3D
F996
F892
F844
F8F3
F9DD
FA35
F9DD
F93A
F8B0
F87F
F8BB
F91F
F954
F96B
F9AD
F9E2
F982
F8D5
F8DD
F9B7
FA07
F8F7
F827
FA4C
FFE3
0645
0A75
0C11
0CBA
0D51
0D31
0C16
0B33
0B90
0C79
0C94
0BD1
0B31
0B20
0B16
0ABF
0A79
0AAB
0B46
0C44
0DDD
0FD4
1107
108E
0F22
0E7D
0F2C
0FF6
0FD2
0F56
0F85
1010
0FF9
0F4B
0F03
0F67
0F87
0EC7
0DF2
0E22
0F18
0F89
0EF7
0E50
0E5E
0E82
0DAB
0BFC
0AAB
0A69
0AB2
0ABA
0A5A
09FA
09FB
0A54
0AA9
0AB6
0A93
0A9A
0AEE
0B4B
0B4D
0AE2
0A4E
09DE
0996
095B
0931
0919
08E6
089F
08E6
0A57
0C5E
0D98
0D87
0D28
0D6A
0DE6
0DD0
0D71
0DA8
0E53
0E53
0D6A
0CEB
0DB7
0E89
0DB5
0C18
0C34
0DEC
0D6A
07B9
FF02
F85D
F617
F61B
F5D6
F577
F666
F815
F866
F6D5
F54B
F55B
F637
F668
F613
F636
F6AC
F682
F5D7
F5CE
F6A9
F744
F6C4
F5D9
F5AB
F629
F64A
F5BA
F548
F577
F5C2
F5C0
F5F6
F6CD
F796
F79D
F775
F833
F9A4
FA74
F9FF
F913
F8B8
F8E9
F8FD
F8CA
F8BF
F8F4
F8F2
F891
F851
F874
F87B
F80B
F798
F79F
F7C7
F78E
F731
F73B
F77E
F75D
F6E4
F6DA
F797
F860
F854
F797
F710
F731
F7A4
F823
F8CA
F961
F93C
F85D
F7C4
F80D
F891
F878
F805
F7ED
F82C
F844
F848
F8A6
F91F
F8F9
F874
F8DF
FA6C
FB08
F930
F76C
FA74
0328
0C8E
114B
1160
10B4
1148
118D
1017
0E59
0E75
0FFD
10A6
0FA4
0E5F
0DCC
0D10
0B91
0A7B
0AD4
0B78
0ABE
0930
08DB
0A3D
0B9B
0B7C
0A6C
09C4
09BB
099A
0945
095C
09E7
0A06
0974
0927
09BF
0A5C
09FD
0944
09A4
0B46
0CE1
0D81
0D78
0D8D
0DFF
0E85
0ED3
0EC0
0E33
0D4D
0C9F
0CC5
0DA2
0E64
0E77
0E17
0DC6
0DBF
0E09
0E8E
0ECF
0E41
0D50
0D14
0D93
0D4E
0B49
08CA
07ED
08EB
09EA
0995
08C6
08F0
09C9
09C3
0892
079C
07CA
085E
088E
08C5
095B
0972
0874
077E
07D7
08AE
083B
06E5
0745
0A0D
0BAC
07F3
FF9E
F815
F54D
F5F3
F683
F618
F63A
F766
F838
F7DD
F74B
F788
F82B
F844
F7E1
F7B9
F7C5
F758
F690
F69C
F7F9
F96A
F97B
F85C
F75A
F709
F6E5
F681
F617
F604
F651
F6D4
F741
F73D
F6B5
F626
F63B
F70C
F7F2
F84A
F837
F83D
F860
F82A
F79F
F76E
F7D9
F829
F7BC
F706
F6EC
F782
F81A
F84B
F84A
F863
F8A1
F8EA
F925
F931
F8FF
F8C6
F8D8
F924
F91C
F86C
F7A2
F78C
F80B
F843
F806
F811
F8AA
F8F3
F857
F79A
F7B9
F866
F89F
F854
F84E
F88F
F805
F661
F530
F5EA
F797
F7F0
F6C8
F66E
F7FD
F94E
F82B
F657
F816
FEDC
072C
0C4D
0CE6
0B2E
09B5
0957
0A02
0BBD
0E17
0FB9
0FB9
0EDF
0E9D
0F26
0F6F
0EF2
0E66
0E93
0F3A
0F8E
0F53
0F0A
0F1B
0F48
0F27
0ECD
0EA6
0ECD
0EE3
0EA7
0E55
0E35
0E11
0D57
0BDB
0A5C
09EB
0AAE
0B79
0B0D
09A4
08A4
08C5
0947
093A
08CF
08CF
0935
0939
08A0
0838
08A3
0948
0923
0855
07F9
0876
08FA
08F3
0923
0A76
0C8C
0E26
0EB9
0EB2
0E77
0DF9
0D62
0D53
0E04
0EAA
0E68
0DA4
0D82
0E2C
0E88
0DF5
0D4A
0D7B
0E20
0E38
0DD4
0DDD
0E6C
0E71
0D46
0BAB
0A92
09B4
086B
0772
0843
0A42
0A10
0503
FCBC
F5F9
F3CE
F508
F667
F645
F56B
F502
F4F5
F49E
F40E
F402
F4CC
F5E0
F67C
F655
F5BE
F568
F5DA
F6E3
F79D
F762
F697
F644
F6D1
F78A
F793
F707
F6C5
F72C
F7A9
F79B
F745
F75D
F80E
F8C8
F8FE
F8AF
F82F
F7D4
F7D0
F82A
F8A0
F8C6
F863
F7C1
F75E
F75C
F76B
F73E
F6EF
F6BA
F6AA
F6B0
F6D0
F70E
F73A
F71E
F6C8
F67B
F664
F684
F6C0
F6EA
F6D3
F67D
F631
F655
F704
F7F4
F8BD
F92D
F931
F8B7
F7FC
F7B3
F853
F939
F944
F86A
F7DC
F855
F909
F8F9
F881
F8BF
F9A8
FA08
F981
F94E
FA22
FA6C
F8A9
F6FA
F9D9
0243
0B35
0EC2
0C8E
0956
08CA
09FC
0A43
095F
0928
0A37
0B0F
0AAE
0A01
0A09
0A30
09A0
0906
097A
0A69
0A4C
0913
0858
08F6
09D2
09A9
0918
09CA
0BF9
0DF6
0E62
0DCF
0D94
0DED
0E2C
0E14
0DF7
0DDF
0D82
0D01
0CDC
0D37
0DA0
0DAB
0D6D
0D40
0D55
0D8C
0DA4
0D8A
0D70
0D9B
0E04
0E07
0CC2
0A3B
07EE
076F
0877
0932
08B6
081A
0895
099F
09DD
092E
08A1
08BF
08EC
089C
0831
082F
0849
080A
07F0
08C3
09EE
09D8
085E
0785
08EA
0B92
0D5E
0DB0
0D8B
0DB7
0E0C
0E54
0E97
0E86
0DA4
0C89
0CC0
0E4F
0E1E
08D5
FF7D
F779
F4E4
F66F
F7E9
F76F
F65C
F62B
F67F
F68D
F699
F733
F7E5
F7B7
F6C3
F629
F669
F6C4
F696
F651
F684
F6CF
F6A0
F64A
F665
F6A6
F653
F599
F565
F5F9
F679
F628
F573
F549
F5CC
F63C
F624
F5FA
F64A
F6E6
F746
F755
F75A
F76D
F77E
F79C
F7CC
F7DB
F7AE
F784
F789
F780
F731
F6F0
F740
F801
F86F
F812
F760
F72B
F7A0
F82A
F841
F7E2
F739
F676
F606
F661
F73D
F7AA
F75F
F737
F7D3
F868
F7BA
F5EC
F48C
F4B2
F5D2
F6A9
F6B8
F65E
F5E9
F560
F515
F56F
F602
F5E7
F559
F5CB
F7A6
F916
F887
F7B2
FA6C
01F8
0AC3
0FD0
0FD1
0DE1
0D70
0ECD
1011
102C
0FC0
0F8D
0F62
0ED5
0E26
0DE4
0E31
0EBB
0F3A
0F90
0F83
0EB3
0D17
0B57
0A56
0A50
0AA0
0A90
0A22
09CD
09BF
09AF
0987
09C8
0AFA
0CD0
0E4F
0EE2
0EED
0F08
0F03
0E63
0D8D
0D8F
0E85
0F26
0E73
0D36
0CFA
0DF3
0ECB
0E99
0E0A
0E24
0E9E
0E61
0D5D
0CCD
0D5C
0E20
0E05
0D60
0D3E
0DA2
0D92
0CC3
0C39
0CDF
0E2C
0EB8
0DE1
0C6B
0B79
0B73
0C08
0CC5
0D5D
0D95
0D6C
0D28
0D01
0CDB
0C9C
0C77
0C92
0CAD
0C6F
0BFE
0BC6
0BCB
0B99
0B0E
0AD6
0BA1
0CE2
0CDE
0A54
060C
0256
0103
01E9
0353
03AE
02D6
01EB
01ED
02A9
0321
02EC
029B
02C5
0327
0321
02AA
024E
0248
0236
01E3
01CF
0274
0345
0336
0252
0217
03CA
06EA
09CB
0B6A
0C03
0C37
0C30
0BD6
0B48
0AE6
0AED
0B59
0BF3
0C5B
0C28
0B5A
0AA3
0ACB
0BB4
0C63
0C45
0BE6
0C0A
0C84
0C8A
0BF6
0B73
0B49
0AA5
0891
056B
02C8
01CE
0211
0250
01EA
0141
00E0
00D0
00C7
00A7
009C
00D6
0146
01A4
01BA
019A
0182
0181
0172
014A
0146
0190
01D0
018A
0102
017D
03FA
07C7
0AD9
0BE0
0B85
0B4F
0BBB
0C05
0B9C
0B13
0B3B
0BE9
0C2B
0BAE
0B2B
0B55
0BCA
0B99
0A97
099F
098B
0A42
0AEE
0AF0
0A75
0A1D
0A23
09E9
0865
053C
0177
FEEA
FE9E
FFD2
00CC
00A6
FFF9
FFC4
0025
007E
0091
00C2
0147
01A4
0151
009B
005F
00F1
019E
0198
00FA
0093
00CD
0132
0132
0113
01D8
042E
0783
0A54
0B79
0B24
0A7D
0A60
0AA6
0AAF
0A4C
09E1
09C0
09C2
09AA
09A1
09F3
0A70
0A87
0A14
09AA
09C1
0A0B
09EC
0976
0960
09F3
0A5F
0967
06B0
033D
0092
FF7C
FF99
FFE9
FFCB
FF74
FF8B
003C
00DB
00A8
FFD3
FF48
FF6A
FF95
FF29
FE8C
FE92
FF2B
FF68
FEF4
FEBD
FF9E
00DC
00EB
FFC0
FF6D
01CC
061F
09BF
0AEA
0A39
096C
0971
09EB
0A2C
0A0F
09E4
09DF
09E5
09C9
097C
091E
08E9
090D
097D
09F8
0A3E
0A35
09C7
08FC
083C
0832
0900
09A9
08BF
05CF
0201
FF2F
FE4B
FEC0
FF49
FF3B
FEE0
FEC9
FEFD
FF04
FE8E
FDE7
FDAE
FE1B
FEBC
FEFE
FEE4
FEDE
FF1B
FF52
FF54
FF54
FF68
FF2B
FE71
FE0C
FF55
0291
0643
087A
08B9
0835
0827
087E
086F
07D1
0763
07C3
08AB
0950
093E
08B3
083A
0808
07D8
076B
0702
071D
07CB
0874
0894
0876
08CB
096A
08EC
0624
01DA
FE72
FD88
FE5B
FEF1
FE63
FD7D
FD4D
FDC6
FE14
FDD6
FD7C
FD8D
FDF3
FE33
FE25
FE11
FE2F
FE50
FE33
FDF2
FDF6
FE69
FEE2
FEC5
FE27
FE11
FF9C
02AC
05DC
07C2
0822
07C1
0766
074D
075E
0784
07AA
07B8
07B0
07BD
07F8
082D
0811
07BB
0797
07DC
0848
087B
0858
07F5
0794
07AA
086D
0915
0811
04AF
0061
FDAE
FDA8
FEE8
FF5F
FEAE
FE1A
FE67
FECA
FE53
FD68
FD2A
FDC2
FE3B
FDFB
FD8F
FDC1
FE6B
FEAD
FE24
FD74
FD6F
FE04
FE4E
FDBA
FCEA
FD4C
FFC2
0397
06DC
0805
0747
0634
0601
0685
06F7
0716
0732
0772
07A5
07B2
07CB
0805
0811
07B2
0733
071E
076B
076E
06C5
05FF
0609
070E
0819
07CA
0565
0184
FDEB
FC44
FCAC
FDAF
FDDF
FD3F
FCCF
FD02
FD3B
FCE8
FC7E
FCC7
FD92
FDD6
FD40
FCB6
FCF5
FD74
FD42
FC99
FC96
FD84
FE37
FD8B
FC0A
FB99
FD87
0140
04EA
06FE
0740
0683
05DF
05EA
0666
06B4
06A8
06AE
0713
077A
0756
06B3
061E
05EC
05F7
060D
0643
069E
06BA
0636
0575
056E
066E
0752
0679
0372
FF90
FCC9
FC1C
FCEC
FDBE
FDA1
FCE3
FC72
FCAC
FD0B
FCF8
FC97
FC72
FCAA
FCD6
FCC9
FCE4
FD63
FDAD
FD0B
FBE7
FB8F
FC72
FD55
FCEE
FBE3
FC5E
FF77
03C3
06C5
076D
06C2
0649
0671
06AC
068D
0642
0610
05F2
05C5
0592
0588
05B7
05F7
0615
0610
0625
0682
06E5
06CD
0622
058E
05D9
06CB
0701
0529
0188
FDF3
FC1E
FC2A
FCDE
FD1D
FCC9
FC66
FC4A
FC5B
FC62
FC5A
FC5A
FC5F
FC50
FC34
FC39
FC6F
FC95
FC58
FBD2
FB9D
FC30
FD24
FD71
FCA8
FBD7
FCC8
000F
0430
06E7
074D
0670
05E3
061D
0670
064A
05F7
0613
069E
06F7
06B3
0618
05B0
05A3
05B2
05B1
05CB
0629
0683
0659
05A2
0509
052F
05A9
051C
029E
FEE8
FBE6
FAF3
FBA0
FC6B
FC6C
FC07
FC02
FC61
FC80
FC14
FB93
FB8D
FBF2
FC48
FC65
FC86
FCBA
FC9D
FBF2
FB43
FB69
FC6A
FD34
FCCF
FBBE
FBC7
FE2D
0239
05C2
071E
0685
0585
054E
05C2
0603
05A8
051C
04F7
0544
059A
05C0
05E0
0610
0607
0587
04E8
04DC
0585
0620
05E1
0510
04D0
059E
0659
0539
01C3
FD90
FADC
FA7B
FB5C
FBF5
FBCC
FB81
FBA2
FBF5
FBF0
FB90
FB51
FB6E
FB8C
FB44
FAC9
FAB6
FB36
FBC0
FBCB
FB7D
FB6E
FBB3
FBAA
FAF5
FA62
FB70
FEAE
02D5
05C1
065B
0575
04B3
04E2
0574
0584
0502
04A6
04EF
0585
05AE
0540
04C4
04C3
051F
055E
0552
053F
0547
0525
04AE
0459
04C1
0590
0550
02D2
FEB0
FB12
F9B8
FA6F
FB99
FBF9
FBA9
FB60
FB4C
FB13
FAA0
FA75
FAF3
FBB0
FBE3
FB65
FAE9
FB0D
FB86
FB8B
FAF1
FA73
FABA
FB62
FB6B
FAAD
FA71
FC3B
0004
03EC
05EC
05AA
0487
0402
0450
04A4
047B
043C
047D
0514
0540
04B4
040A
040B
04A6
050D
04C3
043B
042D
0499
04DB
04AF
04AA
054A
05D1
04AF
014C
FD14
FA58
FA16
FB33
FBE9
FBA2
FB27
FB46
FBBD
FBB9
FB04
FA53
FA58
FAF2
FB6A
FB5C
FB15
FB07
FB31
FB3D
FB12
FAF4
FB02
FADE
FA38
F99A
FA46
FCF3
00CF
03FB
0538
04EE
0475
0496
04F7
04F7
04A0
0488
04E9
0553
054B
04F5
04CE
04E9
04CD
0437
03A7
03D7
04B7
0551
04EF
0417
03FD
04E5
0569
03C7
FFE6
FBC6
F9A7
F9EE
FB0B
FB58
FAB5
FA32
FA7F
FB27
FB59
FAFA
FA94
FA80
FA81
FA4F
FA1B
FA45
FAAB
FABF
FA4F
F9E9
FA22
FAC2
FAEF
FA66
FA23
FB87
FEC4
026B
04B1
0513
048E
045C
04B6
04EF
0497
0415
0417
049E
0503
04D7
0479
0490
051E
056F
0505
0444
03F2
0431
045D
03FF
038A
03BB
0455
03FD
019F
FDDE
FABC
F9C4
FAA7
FBCA
FBFC
FB61
FAD2
FAC0
FAE7
FAE5
FAB3
FA76
FA35
F9E8
F9C4
FA09
FA92
FAC5
FA47
F98A
F95E
F9EA
FA67
FA24
F99A
FA24
FC91
0024
032C
0484
0461
03C6
0376
0385
03B5
03E4
0418
0449
0453
0428
03FB
041C
0495
04F8
04CC
0427
03B1
03E7
046C
0471
03D9
0384
0423
04E7
0409
00E1
FCF4
FA81
FA30
FAB7
FAB2
FA36
FA31
FACF
FB2C
FAAF
F9ED
F9CB
FA3D
FA61
F9C4
F8F5
F8C2
F93E
F9D5
FA09
F9E2
F9B0
F9B3
F9F9
FA4F
FA4B
F9B9
F92D
F9DA
FC6B
0016
0329
0485
0473
03F8
03C1
03D6
0403
0429
042D
03F4
03A6
03A7
0412
0477
0464
0402
03DF
041B
0439
03EC
03A0
03E0
045D
0437
034B
02B3
0362
0488
0402
00C3
FC4F
F95E
F91B
FA41
FAD3
FA44
F98E
F98C
F9FB
FA19
F9C6
F98D
F9C4
FA20
FA38
FA0A
F9D6
F9B8
F9A3
F99A
F9A5
F9A9
F993
F990
F9D2
FA19
F9D9
F92E
F94E
FB6D
FF26
028D
041C
0414
03C0
03BD
03A6
0338
02FC
036E
0421
043C
03B3
034A
0374
03BF
03B6
039C
03DF
043A
0413
0390
0379
03FE
0444
03B2
0312
0393
04C0
047A
0179
FD1B
FA11
F977
FA12
FA3F
F9CE
F99E
FA08
FA70
FA47
F9C3
F968
F957
F96A
F9A3
FA0D
FA60
FA48
F9F2
F9E8
FA45
FA78
FA21
F9B7
F9DF
FA4E
FA0E
F918
F8F0
FB1C
FF18
029B
03ED
0388
0314
0357
03B6
0388
0319
0315
037D
03BF
039D
0374
038F
03BB
03B4
03A1
03C1
03DF
0398
0324
0331
03D8
0436
039F
02BD
02C9
03AB
0399
011C
FD08
F9D0
F8F2
F9B0
FA53
FA24
F9A8
F967
F94C
F924
F91A
F95C
F9AC
F9AF
F97B
F96D
F98C
F97B
F930
F922
F98F
F9F6
F9CF
F974
F9AD
FA63
FA78
F96C
F89C
FA0C
FDEF
0212
0417
03D4
0305
0305
0397
03DC
03B3
039E
03C9
03CF
037C
0332
0350
039F
03B3
038D
0381
0397
038E
036A
038C
03FD
041C
0378
02B9
02F8
0417
0456
022B
FE28
FA8F
F906
F932
F9A6
F9A7
F98E
F9D0
FA39
FA56
FA17
F9C0
F982
F96A
F991
F9FD
FA58
FA37
F9B7
F979
F9CD
FA37
FA1B
F9AC
F9B9
FA5D
FA93
F998
F864
F90D
FC6F
00E6
03D4
0433
034E
02F8
03A2
045D
045C
03D2
0360
033B
0325
0306
0313
0365
03BC
03CD
0392
033E
02F4
02C9
02D8
0324
0366
0355
031F
0350
03EB
03DE
01E9
FE2E
FA72
F888
F89C
F95F
F9A5
F964
F933
F944
F94D
F929
F90A
F912
F911
F8EC
F8DF
F91D
F964
F950
F8F2
F8BE
F8E3
F918
F932
F979
FA14
FA62
F9A7
F878
F8C3
FBD3
0083
040B
04BC
0386
0298
02EC
03A5
03A6
0305
02AB
02F6
0356
032F
02AF
0278
02C5
0334
0351
0315
02D6
02E1
033D
03A3
03AE
032D
027D
0259
0300
0391
029A
FF9F
FBE0
F951
F8BE
F946
F99B
F967
F939
F971
F9C6
F9DF
F9DC
FA06
FA3D
FA22
F9BF
F985
F9A1
F9B8
F97F
F93B
F94E
F98E
F98A
F951
F968
F9D5
F9DB
F92D
F900
FB0C
FF43
034D
04D3
03F4
02D8
0309
03F7
043B
0393
02FB
031D
037D
0357
02C1
0273
02C7
0369
03D9
03EA
03A7
032F
02C2
02AE
02F6
0338
0336
0348
03C7
0413
02CF
FF73
FB5C
F8B1
F848
F904
F95E
F909
F8C2
F8F3
F92F
F90A
F8C7
F8E2
F949
F984
F97C
F98A
F9C5
F9C2
F93E
F8B3
F8C6
F960
F9CF
F9C6
F9B0
F9C9
F98E
F8AC
F830
F9DA
FDF5
0278
04D8
0499
0376
0320
0384
0386
02D4
0244
0284
0332
0379
031F
029F
0269
0277
0299
02BD
02CF
02B4
0289
029C
02F1
0311
02B7
026E
02F0
03C6
0337
0022
FBAF
F875
F7DA
F8CB
F956
F8E7
F876
F8CD
F979
F9AA
F95F
F93B
F975
F9A5
F997
F9A1
F9F5
FA28
F9DB
F96E
F981
F9F2
F9F6
F952
F8CA
F8F9
F951
F905
F8B4
FA22
FDE2
021C
0452
0413
0322
0321
03D6
0419
03A0
0331
0356
03A6
0393
032E
02D2
0289
0241
023C
02B2
0335
0317
026B
0215
0293
033F
034A
0301
0358
041D
0394
0084
FC16
F8DE
F827
F8D8
F926
F8A1
F831
F87C
F917
F94B
F90A
F8D0
F8DE
F90F
F941
F977
F99A
F980
F942
F945
F9AA
F9FD
F9C6
F941
F921
F988
F9A6
F8E3
F81E
F92C
FCC0
013B
0414
045F
037B
033D
03F5
0486
0425
0349
02DE
0312
0354
0345
030A
02D8
02AD
029D
02E7
036D
0395
0311
0276
0287
0317
0339
02AD
025C
02DE
0316
013A
FD50
F9A6
F84B
F8D6
F953
F8D8
F839
F861
F8F6
F919
F8C6
F8B0
F90D
F957
F943
F937
F974
F991
F93D
F8F5
F94D
F9DA
F9B9
F901
F8D1
F9A4
FA5F
F9D7
F8CF
F986
FCF1
014D
03F0
0417
0332
02D9
033D
03AA
03BC
039D
0383
036A
0349
0333
031D
02E0
028F
0287
02EB
034A
0324
02A6
0281
02F2
0368
034C
02E7
0307
03BE
03D1
01D5
FDE8
F9F6
F801
F843
F939
F96B
F8D2
F86C
F8C9
F96C
F993
F931
F8D5
F8D8
F906
F916
F908
F8FD
F8FD
F916
F95E
F9AD
F99C
F917
F8B0
F8F3
F97C
F95D
F8A8
F8F8
FBBA
0016
036D
0427
0351
0301
03C9
0477
0410
0319
02A4
02EA
0349
0358
033C
031C
02DD
02A4
02E0
0383
03BF
0317
0244
025E
0347
03CA
0351
02CC
0330
03B4
0273
FEE9
FAEB
F8B3
F885
F8DF
F89A
F80A
F803
F88B
F8F9
F8EF
F8B3
F8AB
F8EB
F954
F9BF
F9E0
F96F
F8A4
F844
F8CC
F9B1
F9F6
F970
F8FE
F944
F9A9
F931
F827
F84A
FAF5
FF58
0311
046D
03CB
02CB
0285
02E7
0365
03BF
03FB
03FC
0397
02EF
0277
0276
02C0
02FD
0319
032C
032E
0309
02DC
02E7
0314
02F7
0284
0266
0326
03FD
031D
FFB5
FB49
F871
F837
F932
F978
F8C6
F84C
F8BA
F95A
F93B
F87D
F811
F872
F92E
F9AD
F9C8
F996
F925
F8BA
F8CE
F96C
F9E1
F98E
F8DF
F8CE
F96F
F9B6
F912
F8BA
FA74
FE34
01C6
033A
02EB
0296
0307
0386
035C
02E9
02E3
032E
0329
02CE
02C1
033B
03A0
0366
02E8
02C4
02E4
02C0
0264
0269
02E6
0317
0285
01FB
0282
0399
0344
0055
FC1C
F926
F899
F956
F9B5
F957
F8F8
F90E
F93E
F91B
F8D5
F8DB
F92A
F961
F953
F92A
F90B
F8EB
F8D3
F8FF
F972
F9C5
F99D
F941
F947
F9AE
F9BD
F921
F8D3
FA3F
FD8B
011F
032C
036F
030F
030C
0349
033F
02F3
02D4
02F6
02F2
029F
025E
028A
02ED
0311
02EF
02E0
0300
0303
02CE
02BE
030C
0350
030C
028B
0295
0319
02BD
0054
FC8C
F98B
F8AE
F938
F978
F8D5
F82D
F85A
F912
F97D
F968
F95E
F9B2
FA06
F9EA
F97E
F92F
F91E
F91A
F91D
F958
F9B6
F9C6
F94B
F8A7
F866
F88B
F8C8
F951
FAE1
FDAF
00C2
02C7
036B
0372
0393
03B2
0373
0303
02E0
030C
0308
02AB
0268
0291
02C8
029A
0246
025F
02E3
0336
0317
02FF
034C
038B
0326
0286
02B6
03AE
03C8
0182
FD78
F9F6
F890
F8C9
F91E
F8D4
F86B
F890
F927
F98F
F96B
F8F9
F8B2
F8D6
F949
F9B4
F9D3
F9B5
F9A2
F9B3
F9AF
F962
F8F9
F8CB
F8EF
F92C
F948
F933
F8F4
F89F
F890
F966
FB7D
FE61
0100
029B
034D
03A2
03DE
03E6
03A5
0342
02F4
02DD
02FB
0330
034C
0338
030E
02F5
02EA
02CD
02A3
02A9
02F8
0345
0346
032B
0359
039F
034F
025F
01D2
0278
0374
02C9
FF96
FB50
F863
F7D3
F896
F922
F909
F8E1
F918
F974
F985
F92C
F8A9
F862
F896
F923
F997
F9AA
F97F
F966
F967
F94E
F910
F8EE
F916
F956
F973
F994
F9E7
FA12
F992
F8EC
F9AF
FCB4
00BC
037D
03FB
034D
02FD
034F
037C
032D
02F5
034D
03CD
03CB
0352
02F8
0306
033B
0352
034A
0333
0306
02BD
0277
025D
0283
02DC
0336
0345
02E2
026A
0283
032D
032E
0117
FD1F
F96C
F809
F8D8
F9F1
F9DF
F8EF
F851
F889
F917
F95E
F956
F944
F938
F917
F8F9
F91C
F985
F9E9
FA04
F9DA
F9A7
F995
F98F
F959
F8F9
F8DD
F952
F9DF
F9A4
F8A6
F862
FA71
FE95
0299
0466
0400
031F
0302
0354
0339
02BC
029A
0314
03A0
03AA
033F
02CD
02A5
02C9
0309
0338
033F
0326
030C
0305
0314
0334
0366
0383
0345
02BE
0299
0349
03E1
0292
FEC2
FA45
F7BD
F7F9
F969
FA27
F9DF
F975
F970
F972
F92A
F8F8
F949
F9C9
F9D7
F966
F8FC
F8F0
F913
F921
F921
F945
F998
F9DE
F9CC
F960
F90B
F944
F9E2
FA12
F959
F894
F986
FCED
013B
03DC
03D6
02A5
024C
0320
03F6
03F3
036D
0319
031C
0323
0304
02E5
02EC
0306
0314
0317
0319
0312
02FF
02F5
0302
0322
0353
0378
0342
0298
0217
028C
0390
0364
00C9
FCB1
F983
F894
F906
F93D
F8D5
F89E
F90B
F980
F96B
F924
F94A
F9C6
FA0D
F9FB
F9DE
F9CF
F9A0
F94D
F90E
F906
F919
F92D
F94B
F973
F994
F9BE
FA18
FA65
FA01
F8E7
F88F
FAC2
FF37
033D
047E
0375
027E
02E3
03C3
03D1
0314
027E
0279
0291
026E
0267
02D4
0362
038B
035C
0348
0373
038F
0360
0305
02CB
02DC
0318
031B
02B6
0261
02D2
03D0
03E3
01B1
FDBC
FA34
F8D9
F952
F9F1
F9CC
F96C
F97F
F9CA
F9C5
F992
F9A4
F9EA
F9ED
F999
F94D
F942
F953
F958
F962
F97E
F989
F96F
F95A
F96E
F989
F97D
F979
F9A7
F9A0
F8F7
F87E
F9F5
FDD7
022F
0469
0414
02F6
02B5
0331
035E
02F6
02A0
02CC
0320
032E
0315
0325
0342
0324
02DF
02BE
02D5
0307
0348
038B
03A8
0398
038D
0384
0337
02B5
02AF
0389
0445
0317
FF70
FB1D
F89F
F89F
F98F
F9E2
F9A5
F9A0
F9D5
F9BA
F959
F952
F9CF
FA41
FA27
F9A6
F934
F90F
F92C
F96A
F9A5
F9AF
F978
F93F
F944
F969
F96F
F984
F9EE
FA44
F9C6
F8E3
F96D
FC70
008B
0339
0392
02E7
02C7
034B
039A
0367
032D
0330
031A
02BD
0280
02B8
0318
034E
0386
03E9
0414
03B4
0325
02EF
0300
02F2
02CB
02DD
030F
02F1
02A9
02F9
03E6
03E7
016B
FD20
F9AB
F8BA
F958
F9B2
F974
F985
FA1A
FA69
FA02
F976
F966
F9A7
F9AC
F95E
F921
F92C
F956
F97D
F9B5
F9E4
F9C4
F96A
F94F
F991
F9C0
F9AE
F9C3
FA08
F9C8
F8D8
F89C
FABC
FED9
0291
03F5
0376
02E3
031E
0384
0361
0304
02F9
031B
0308
02EA
031C
037A
03A7
03A8
03AC
0390
0326
02B8
02B7
0311
0347
0333
0332
0366
0365
0302
02F7
03DB
0498
0321
FF26
FAFC
F917
F964
FA05
F9E9
F99F
F9CE
FA23
FA0A
F9AD
F9A3
F9FD
FA2F
F9E8
F96E
F920
F905
F923
F9A7
FA66
FAC2
FA75
F9F2
F9A7
F96D
F920
F927
F9B3
FA0E
F983
F8D5
F9D9
FD3D
0156
03B9
03C9
02F8
02B3
02E7
02EC
02D1
0311
038F
03C3
0390
0351
0339
033B
035A
039E
03C5
0386
030B
02CF
02F9
0323
0307
02FE
0363
03CC
0393
0315
035D
0441
03E8
0101
FCC2
F9C2
F921
F9C1
FA16
F9D3
F99C
F9C3
F9EF
F9CB
F977
F93F
F93C
F966
F9B4
F9EE
F9D6
F997
F9AE
FA18
FA3E
F9E5
F99D
F9CB
F9F7
F9A8
F952
F9A6
FA3B
F9EB
F8C9
F8B4
FB49
FF95
02E2
03C4
035E
0360
03E4
03F7
0375
0328
0372
03D0
03C0
0366
0333
0352
03A3
03EE
03F6
0392
02F7
02B7
0324
03CB
03F0
0391
0358
0376
0360
02F6
02FB
03C3
0403
0216
FE35
FA94
F91A
F991
FA53
FA48
F9B9
F966
F97B
F9AE
F9CC
F9D1
F9C0
F9AF
F9C8
F9E6
F9A8
F90B
F8A6
F8E2
F96B
F9BA
F9D8
FA0D
FA32
F9E4
F952
F931
F9A0
F9C3
F911
F8B1
FA84
FEA1
02B1
0464
03DF
0312
032D
03AC
03A6
032B
02FA
0368
03FF
0419
039A
030F
030F
03A3
0430
040B
0341
02AA
02FC
03D8
0439
03D2
035A
035E
0380
0359
0364
0429
04D8
03A9
0007
FBAC
F90C
F8E0
F9BE
FA0D
F9A4
F952
F974
F9AA
F9A3
F984
F988
F9B2
F9E1
F9F9
F9E8
F9B5
F989
F98C
F9C3
FA0C
FA44
FA42
F9E5
F943
F8D3
F915
F9E1
FA44
F992
F8A4
F963
FCAB
0107
03FD
0478
0392
030B
037B
041D
0415
0377
030A
0343
03BD
03C8
033F
02C2
02F7
03C2
045A
0431
03A3
036E
03B4
03DD
038C
0327
0328
035E
0354
032B
0372
03FC
038A
0115
FD49
FA2B
F91D
F99B
FA1B
F9D5
F947
F932
F99B
F9F3
F9E8
F9B8
F9C4
FA09
FA23
F9D9
F969
F943
F97F
F9CB
F9E4
F9E2
F9FC
FA18
F9EA
F988
F982
FA26
FACB
FA72
F93A
F8CE
FAD3
FEFD
030F
04F4
0499
0396
034D
03AD
03D4
036D
0307
033D
03DF
0440
040E
039C
035C
035B
0353
032D
031B
0336
034C
032A
0305
033D
03D1
043B
0417
03B5
03BE
042E
0406
0233
FECF
FB46
F927
F8D4
F96A
F9D8
F9D3
F9C1
F9EC
FA18
F9F6
F99F
F97F
F9BE
FA0D
FA12
F9E1
F9DB
FA22
FA6A
FA5C
FA0E
F9E6
FA17
FA68
FA80
FA4B
F9FA
F9B7
F97A
F93F
F970
FAC2
FD81
00EF
039E
049E
0447
03B5
0399
03BC
03AA
0378
039B
0414
0450
03EF
0359
0330
0376
039F
0365
031E
032B
0362
0353
02F9
02D5
0339
03BF
03BF
0339
02EB
0367
0420
03B4
013D
FD6B
FA1D
F8C0
F916
F9C0
F9DD
F9B5
F9DD
FA34
FA29
F9B6
F985
F9F9
FA8A
FA78
F9D5
F96F
F9B7
FA3F
FA76
FA6B
FA83
FABC
FAB9
FA68
FA27
FA3B
FA73
FA7F
FA5D
FA3D
FA23
F9F7
F9F2
FAB7
FCB9
FF9F
0266
0421
0490
042D
03BB
03B7
03F8
03FE
039C
0339
0347
03AA
03E3
03B1
0350
0319
031D
032E
0334
0347
037B
03B6
03D3
03BC
037A
0334
032C
0370
0398
0338
029E
02A4
0372
03D1
024C
FEF5
FB93
F9D6
F9C2
FA1E
FA20
FA0D
FA4A
FA8D
FA57
F9D1
F99F
F9F8
FA72
FAA5
FAA3
FAAA
FAB5
FA90
FA34
F9E4
F9DB
FA09
FA30
FA3C
FA53
FA8E
FAC6
FAC0
FA88
FA6B
FA91
FAA5
FA36
F9A1
FA42
FD1A
0146
0466
04ED
03AC
02AF
02EC
03A0
03C7
0372
035B
03A7
03C8
037F
0344
0381
03E7
03F2
03B5
039F
03BF
03C1
038D
036B
037B
0374
0322
02D2
02F3
0362
0390
0358
0357
040F
04DB
044A
01A4
FDDC
FAD7
F9C2
FA2F
FAB9
FA84
F9EA
F9C1
FA2E
FA91
FA79
FA31
FA2E
FA5C
FA57
FA1B
FA0E
FA4D
FA64
F9FF
F987
F9A0
FA39
FAA5
FAA4
FAAB
FAF7
FAFF
FA5C
F9AB
F9D0
FA89
FA9C
F9AD
F939
FB02
FED5
0283
042E
0412
03AD
03CB
0401
03CD
0371
0379
03EC
044C
0439
03D7
0391
039A
03CC
03F2
0401
0403
03EB
03A9
0362
0359
039E
03E6
03E3
03A7
038D
03AC
03AB
0361
0354
0406
04C2
03DE
00A4
FC87
F9DF
F98A
FA55
FAB1
FA55
F9FB
F9FD
F9F6
F9AC
F987
F9DB
FA45
FA3A
F9E6
F9E1
FA3D
FA64
FA07
F9A3
F9D0
FA61
FA9C
FA39
F9C3
F9D3
FA42
FA73
FA48
FA45
FAAE
FAF2
FA69
F981
F9BE
FC2C
FFFB
0306
03F0
036E
033D
0403
04D3
04B6
0408
03D5
0454
04AF
0444
0384
0348
03A8
040B
041B
041C
043A
0424
03A9
0343
0379
0407
0425
03A7
033B
0361
03B4
0397
034A
03A2
0495
04BB
02BC
FF08
FB9B
FA06
FA10
FA6E
FA51
F9F6
F9DE
FA03
FA09
F9DA
F9C9
F9FB
FA2A
FA10
F9DB
F9EC
FA36
FA49
FA00
F9CC
FA17
FA9E
FAC1
FA67
FA27
FA69
FAC8
FAAD
FA45
FA49
FAC2
FACE
F9F6
F951
FA94
FDFC
01C2
03E6
0421
03B4
03AD
03EC
03EB
03C2
03EE
046B
04A5
0458
03F7
0403
0455
0461
040B
03CC
03F6
0435
0406
0386
0359
03C4
043A
0417
037F
032F
0371
03C3
03A6
0372
03D2
0485
0426
01A2
FDB4
FA71
F94E
F9D9
FA86
FA6D
F9E5
F9A6
F9D1
F9FA
F9D9
F999
F98A
F9BD
FA09
FA42
FA54
FA3E
FA19
FA1A
FA5A
FAA8
FAB6
FA7E
FA59
FA91
FAF1
FAFC
FA99
FA3D
FA58
FAA3
FA74
F9D3
F9EB
FBEE
FF92
0302
048E
0441
0386
0382
0415
0480
048B
049A
04DF
04FD
04A3
0418
03E3
0415
0448
0435
03FF
03DA
03B4
0371
0342
0372
03E6
0423
03EA
0399
03AA
03FD
040A
03B8
03A1
041C
044F
02D4
FF6C
FBB4
F9BA
F9EB
FAC9
FABD
F9CF
F92F
F977
F9F9
F9E4
F96A
F954
F9D0
FA43
FA49
FA42
FA9F
FB13
FAFD
FA66
FA0F
FA5B
FAC2
FAA4
FA3C
FA39
FAA6
FADB
FA8A
FA3B
FA6E
FABC
FA6A
F9D7
FA8F
FD8F
01C1
04CC
0563
0463
0396
03CC
0470
04AA
0466
041F
0419
0421
040E
0408
042D
0441
0401
039B
038D
03F1
0452
044F
0419
0415
042F
0400
038A
0368
03E8
0468
041E
035E
034C
0415
0424
01D7
FDAD
FA15
F8E4
F990
FA41
FA0F
F9AD
F9F1
FA97
FABE
FA36
F9AB
F9B0
FA1D
FA80
FAAF
FAC2
FAB6
FA6F
FA06
F9C9
F9E0
FA18
FA2C
FA2B
FA56
FAA8
FAC9
FA95
FA70
FABD
FB31
FB02
FA11
F999
FB2F
FEED
02F8
052B
052C
0474
045D
04C4
04BD
0420
03B3
0401
0496
04BB
0470
0441
045C
045D
040B
03CC
0406
0470
047A
041E
03E7
0419
0456
0435
03E4
03D5
0400
03EC
0385
036F
0419
04BE
03D8
00CA
FCDB
FA1F
F984
FA24
FA80
FA1A
F9A7
F9DA
FA6A
FA95
FA33
F9DC
FA00
FA56
FA5C
FA17
F9F0
FA08
FA0B
F9D1
F9BB
FA28
FAD0
FB0D
FAC0
FA6F
FA7B
FAA1
FA8E
FA7A
FABC
FB03
FA9D
F9C5
F9F8
FC76
008F
03F8
050B
0452
03A0
03FB
04CE
0513
04A1
041F
040B
043A
0447
0428
041C
043A
0457
0453
0447
0448
043A
03FF
03C9
03DF
042F
044A
03F9
0398
039D
03ED
0400
03C3
03D0
046E
04A0
02EB
FF3F
FB7F
F9BB
FA14
FADB
FAAA
F9D0
F972
F9E0
FA65
FA75
FA67
FAB6
FB23
FB0C
FA6E
F9F3
F9FD
FA31
FA16
F9DA
FA00
FA8C
FAE9
FAC9
FA9D
FAE7
FB6C
FB76
FAE9
FA79
FA9F
FADA
FA74
F9E4
FABF
FDE0
0203
04C6
0513
041A
03BC
046B
050F
04BC
03E8
039D
0412
048C
047B
042D
042D
047A
04A1
0481
0468
047C
0473
0418
03AF
0399
03B9
03A6
0363
036A
03E8
044F
041D
03C1
0419
04FD
04DA
0259
FE2B
FAA9
F983
FA36
FAF4
FAB8
F9FF
F9B2
F9F3
FA44
FA61
FA7B
FAB1
FAC6
FA8E
FA43
FA2E
FA33
FA03
F9B5
F9C6
FA5D
FAF3
FAF6
FA97
FA93
FB20
FB92
FB4D
FAA4
FA66
FAA2
FA8B
F9DC
F9C3
FBC8
FFC3
0390
0521
0493
03BF
03F5
04BC
04E6
0449
03CA
0403
0481
0491
0440
042D
0488
04D9
04BB
0467
0443
0449
0436
0417
0437
0482
0470
03D8
0362
03BD
0495
04D3
041B
0368
03C2
048B
03D8
00AB
FC66
F995
F964
FAAC
FB77
FB09
FA2B
F9DC
FA2B
FA81
FA83
FA59
FA3A
FA24
FA0D
FA15
FA55
FA9C
FAA9
FA89
FA8C
FAC9
FAF3
FACB
FA8B
FA94
FAD1
FAD5
FA8F
FA82
FAF3
FB4E
FADB
FA1A
FAB0
FDA1
01CD
04CE
0558
0461
03BD
0416
04A9
04B0
0462
046F
04EF
0552
0529
04A7
0443
042C
0440
045E
0477
046F
0438
0407
042C
0497
04BD
0438
0369
0324
03B0
0457
044A
03C0
03BC
0488
04D8
0303
FF13
FB24
F959
F9C5
FAAB
FA9C
F9D5
F96D
F9BC
FA21
FA1E
FA07
FA55
FAD4
FAF1
FA99
FA58
FA85
FAD0
FAC4
FA6F
FA39
FA49
FA62
FA61
FA72
FAB6
FAF1
FAE8
FADB
FB23
FB84
FB48
FA59
F9E6
FB6A
FEFC
02E4
0521
0543
048A
0454
04C5
0519
04DC
046C
044B
0471
047C
0458
044F
0481
04AF
04A4
0498
04D1
0519
04F7
046E
0422
0479
04FB
04F4
046D
041B
044A
046B
03FB
036F
039B
043D
03DC
016C
FDC8
FAED
F9FE
FA60
FAD3
FAD7
FABD
FAC3
FAAE
FA50
F9EF
F9F1
FA4D
FAA0
FAB7
FAAF
FAA7
FA8D
FA60
FA57
FA8A
FAAB
FA5D
F9D3
F9BE
FA63
FB1A
FB08
FA49
F9F0
FA9B
FB7B
FB51
FA45
FA22
FC65
0062
03D1
051B
04AE
0406
03EC
0410
0406
03FD
0445
04B1
04D8
04B7
04A6
04C8
04DF
04BF
0497
0493
0488
043C
03E2
03ED
0462
04B9
049B
0463
0499
0517
0534
04BA
043A
0445
049F
04A3
0441
0416
045F
043D
0285
FF37
FBC6
F9CC
F9A7
FA77
FB2C
FB53
FB05
FA83
FA1E
FA29
FAB6
FB59
FB81
FB16
FA97
FA7E
FAAF
FAB5
FA70
FA32
FA37
FA4D
FA31
FA05
FA25
FA96
FAEB
FACB
FA5D
FA10
FA1D
FA77
FAFD
FB76
FB6C
FA90
F982
F9BE
FC45
004D
03BB
051B
04DC
0479
04BC
052E
0520
04A7
044C
0434
0411
03D2
03D5
044F
04D4
04CC
0438
03B9
03CE
044E
04C0
04EF
04F7
04F7
04EF
04E0
04D5
04B8
046C
0415
0410
0470
04B4
0460
03D0
03EC
04CF
051F
034F
FF82
FBBB
F9E7
FA10
FAB5
FABD
FA69
FA7C
FAF6
FB33
FAED
FA8D
FA87
FAC2
FAE5
FAE6
FAF1
FAFA
FABE
FA4A
FA0F
FA4F
FAB1
FAAF
FA4F
FA19
FA55
FAB2
FACB
FAA4
FA89
FA89
FA89
FAA6
FB24
FBCB
FBDA
FB0A
FA69
FB96
FEEF
02D1
051E
053A
045C
03F3
0443
04A9
04BC
04AB
04A8
048F
0449
041E
0453
04AD
04B2
045A
042B
0478
04EE
050A
04CA
049C
04AE
04BA
0485
0447
044E
0490
04BC
04B9
04A3
0476
0412
03C3
042D
0549
05BD
03EF
FFEC
FBCF
F9CA
FA10
FAF2
FAF9
FA48
F9E7
FA3B
FAB8
FAD8
FAC2
FACF
FAF5
FAF2
FAD0
FAD9
FB10
FB19
FAC8
FA78
FA93
FB01
FB46
FB27
FAE0
FAB9
FAAD
FAAA
FACC
FB24
FB5A
FB0C
FA6E
FA2F
FA82
FAB2
FA35
F9DF
FB55
FF09
033F
059E
0591
049F
0467
04E7
0518
049B
042B
046C
050A
0549
0502
04A4
0470
043D
0400
0405
046A
04C3
04A0
043C
0432
0497
04D2
0475
03DA
03A3
03E2
0429
0447
0475
04B5
049C
040E
03C7
0470
054A
047C
012D
FCDA
FA12
F9E4
FB09
FBA0
FB2E
FA87
FA57
FA5E
FA3A
FA25
FA87
FB27
FB50
FAC8
FA27
FA0D
FA62
FA9E
FA95
FA95
FAD7
FB2F
FB64
FB7C
FB96
FB93
FB52
FB04
FB00
FB3D
FB55
FB2E
FB2F
FB8A
FBAB
FAFF
FA32
FAFB
FE2D
0260
0515
0543
0438
03D7
0485
0534
0516
0493
047A
04DF
0532
0524
04F9
04F4
04EC
04A2
0438
0409
0430
0471
0497
048F
0454
03F2
03AC
03D9
0460
04B0
0462
03DE
03DE
0462
04A7
0449
0404
04A2
0579
04AD
0159
FCF5
FA0E
F9AD
FA92
FAFD
FA96
FA46
FAA1
FB30
FB46
FAEB
FA9B
FA8B
FA97
FAB7
FB0D
FB78
FB87
FB14
FA9F
FABA
FB45
FBA4
FB92
FB61
FB56
FB44
FAFB
FACA
FB11
FB79
FB46
FA83
FA33
FAF1
FBD9
FB9F
FAA0
FAF2
FDF4
0258
055D
05C4
04D9
046F
04BF
04D9
0475
045F
0505
0598
0525
0404
0378
0407
04E4
051A
04B7
045E
0442
041B
03EE
041A
04A3
04EF
04A1
043A
0473
0522
0568
04EE
045C
044B
0463
041A
03DB
0482
05A1
053B
01F6
FD28
F9D5
F97F
FABE
FB45
FA99
FA14
FA9D
FB6D
FB5F
FA9B
FA3D
FAA9
FB18
FADF
FA76
FAB0
FB73
FBDF
FB8D
FB09
FAEF
FB20
FB29
FB0A
FB16
FB3B
FB07
FA79
FA36
FA9A
FB1E
FB13
FAA8
FA9B
FAF5
FAF8
FA84
FAE9
FD7F
01A5
04FF
05EF
0537
04AC
04F3
0533
04CC
0450
048B
0539
056D
04EC
0477
04A4
0510
0512
04BF
04AE
04FF
052E
04E6
047F
046B
0494
049B
0483
049B
04D9
04CB
0455
0400
043B
049F
0480
040B
0421
04DB
04DC
02BA
FEEB
FB95
FA48
FA89
FAD5
FA9F
FA88
FAF3
FB3C
FAB5
F9D4
F9A6
FA5A
FB03
FAF2
FA97
FAB6
FB3D
FB73
FB24
FADC
FAFB
FB22
FAE5
FA94
FAC1
FB48
FB65
FAEB
FA97
FAF1
FB71
FB54
FADF
FAF9
FB9B
FBA2
FAAE
FA54
FC8D
00FE
04E1
05F7
04E4
03FF
046A
053C
0556
04F5
04FB
0570
058C
050D
04A3
04D0
0518
04C3
0408
03C7
043E
04BD
04B6
0480
04A8
0504
04FB
0493
047E
0504
0576
0526
0471
0435
0488
04A8
044E
043B
04D7
04F0
02C8
FE90
FACD
F9C3
FAF1
FBEA
FB57
FA44
FA50
FB62
FC00
FB63
FA5B
F9F9
FA3D
FA7B
FA95
FAF8
FBA1
FBE6
FB69
FAB6
FA8A
FADD
FB12
FAEB
FACF
FB02
FB35
FB21
FB15
FB77
FBFA
FBF4
FB5D
FAE9
FAF7
FAF9
FA7D
FA59
FC11
FFCC
03A5
0583
053F
047B
047A
04E4
04CB
043B
041C
04D4
05A7
05BD
052B
04B5
04BF
04F3
04E5
0494
043F
03FF
03DA
03F3
0462
04E8
0519
04DF
048B
0464
0455
043B
043C
0479
04A3
0454
03D0
03EF
04D8
0540
0389
FFB9
FBE0
FA20
FAA5
FBCE
FC26
FBA2
FB0E
FAD0
FAB2
FA81
FA5A
FA61
FA7C
FA97
FAD7
FB48
FBA3
FBA4
FB76
FB78
FB9C
FB70
FAE0
FA7E
FACD
FB7D
FBC5
FB74
FB2D
FB67
FBC4
FBB2
FB62
FB78
FBD6
FB92
FA72
F9E9
FBCA
FFEB
03E4
0574
04C3
03D2
03F8
04B4
04E7
0479
0436
0481
04DD
04D9
04BB
04EF
0542
052F
04BE
0483
04BF
04FC
04BD
0435
03E9
03EC
03EC
03E4
0436
04D4
0503
0452
0374
0374
0440
04B8
0457
0406
04AC
055F
041A
0061
FC5A
FA92
FB35
FC30
FBE4
FADA
FA7F
FB10
FB7A
FAFE
FA24
F9D5
FA2B
FA97
FAD1
FB0A
FB52
FB5E
FB19
FAF1
FB49
FBDF
FC20
FBF1
FBCA
FBF2
FC1A
FBDD
FB65
FB1E
FB0A
FACF
FA7E
FAAD
FB7C
FC11
FB9F
FAE5
FBC8
FF1E
034D
05C4
05B2
04A4
0471
052F
05A4
0541
04C7
04FE
058F
059C
0509
0485
0487
04C8
04D5
04A2
0454
03E0
034F
0313
0398
047A
04C6
0439
03B3
0412
04FD
0564
04F4
0464
044C
0458
0414
03E8
0474
051C
041E
00B0
FC5F
F9B4
F990
FA8C
FADB
FA37
F997
F9A1
FA08
FA4F
FA83
FAEA
FB64
FB93
FB79
FB7E
FBD4
FC30
FC36
FBF5
FBC0
FBC4
FBF5
FC44
FC99
FCA0
FBFA
FAD3
FA0B
FA5E
FB77
FC3D
FC17
FB91
FB75
FBAB
FB94
FB67
FC6A
FF68
034A
05ED
065F
05BE
05A3
0643
0694
05FC
0523
04E4
0524
052C
04C0
0451
043A
044F
0442
041B
0401
03E4
03A6
0381
03C7
0452
04A1
0491
048C
04C7
04CC
043B
03A0
03DA
04BD
0519
0451
0360
0392
0477
0404
0103
FCC5
F9CB
F931
F9EE
FA7D
FA7B
FA6D
FA99
FAB7
FA96
FA7E
FABE
FB30
FB7C
FB95
FBA3
FBAA
FB8E
FB71
FB9D
FC0B
FC3F
FBEE
FB7A
FB84
FC04
FC48
FBDA
FB26
FADE
FB0F
FB3A
FB41
FB9E
FC6A
FCBE
FBD2
FA8E
FB20
FE99
0353
0671
06C8
05BF
054D
05C4
0615
05AF
052F
0532
0560
051D
049D
049C
0533
059F
0553
04AA
0447
042E
0400
03CA
03FF
049F
04F6
049C
041B
042D
04A6
04BC
0445
03F7
0455
04E1
04DC
0465
043A
047E
0476
03CB
0353
03E5
04C0
03FB
00CF
FCC8
FA45
FA0A
FAD8
FB37
FAFE
FAEB
FB40
FB7B
FB45
FB04
FB31
FB8F
FB77
FAD0
FA4F
FA9E
FB8E
FC4E
FC56
FBD6
FB53
FB18
FB23
FB54
FB85
FB90
FB6D
FB49
FB58
FB80
FB7F
FB50
FB44
FB84
FBBE
FB9A
FB57
FB86
FC20
FC55
FBA8
FB06
FC0D
FF32
02F8
0567
05EC
0579
051E
050B
0501
0510
056A
05CE
05A9
04E9
0437
042E
049F
04EC
04D8
04AF
04B9
04E9
051F
055E
059B
0592
0520
049B
0485
04E1
052B
050E
04D3
04D6
04EA
04A9
0444
0467
052A
05B0
0531
0438
0411
04EA
0523
0300
FED6
FAED
F92F
F972
FA35
FA86
FAA1
FAEE
FB36
FB15
FABA
FAA8
FAEA
FB00
FAAE
FA62
FA8A
FAEE
FB0B
FADD
FADF
FB2B
FB37
FAA7
F9FB
F9FE
FAAF
FB48
FB4E
FB1E
FB34
FB5D
FB1D
FA9B
FA90
FB2F
FBC9
FBCC
FBA6
FC0C
FCB5
FC9F
FBBC
FBA3
FDDF
01DB
053B
0655
05C7
0547
058B
05E3
05A5
0525
0508
054A
056A
0548
0540
057A
05A8
0598
0597
05DC
05FF
0577
0494
0446
04E0
058A
0559
0494
0448
04CA
054E
0525
04B7
04BB
0500
04B4
03C6
032C
0383
0413
03DD
0331
0345
0427
0411
017A
FD40
F9F5
F91B
F9D5
FA75
FA85
FAB3
FB41
FB82
FAF8
FA38
FA1F
FAA2
FAF3
FAAA
FA3A
FA2A
FA6C
FAAD
FAE5
FB2C
FB46
FAD9
FA1E
F9DA
FA67
FB2B
FB61
FB25
FB3C
FBE4
FC6C
FC3E
FBD0
FBF4
FC98
FCCE
FC37
FBAB
FBFA
FC98
FC4A
FB2D
FB28
FDCD
0234
05B4
06AC
05F4
0560
059B
05F8
05E2
05A1
0595
0584
050E
0478
046C
04F7
056C
054F
04EC
04C1
04C8
04B6
049B
04C2
0511
0518
04BD
0476
048B
0497
0429
03A3
03D4
04B0
052B
04A1
03CB
03BA
0442
0447
037B
02F6
039E
047F
03A3
0076
FCA3
FA57
FA16
FAC6
FB51
FB92
FBBD
FBA8
FB22
FA84
FA67
FAC6
FAF6
FA8D
FA08
FA26
FADF
FB65
FB35
FABF
FAC8
FB5C
FBCD
FB9B
FB08
FAB1
FAD3
FB3B
FBAA
FC00
FC15
FBC2
FB45
FB2F
FBA9
FC09
FB8E
FA83
F9FF
FA6F
FAFD
FAE0
FAD2
FC70
000E
03F2
061A
0653
05F6
05EF
05D8
0538
0498
04C2
0565
0571
04A5
0400
0469
0570
05ED
0585
04F7
04F9
055A
0580
0552
052D
0537
0537
0505
04B4
045E
040F
03F9
0463
0535
05D3
05C2
054B
052F
059B
05D5
053B
0444
03FE
048E
04A9
02E4
FF66
FBE9
FA12
F9F7
FA6F
FA84
FA54
FA71
FAE3
FB2F
FB1F
FB14
FB5A
FBA4
FB72
FAD2
FA59
FA6D
FAD7
FB2E
FB58
FB71
FB6E
FB34
FB0A
FB58
FBEC
FC06
FB56
FA8F
FA81
FAF9
FB13
FA8C
FA22
FA76
FB24
FB6C
FB5F
FBA4
FC28
FC07
FB2B
FB27
FD91
01CC
0554
065B
0574
0477
0453
048E
0490
0485
04D4
0553
0590
058A
0598
05C2
05AC
053B
04D7
04D1
04F4
04D5
0481
0472
04D9
0550
0558
0504
04D6
0500
0533
0521
04FB
0522
058B
05BF
0573
04EB
049F
04AF
04E6
0532
05A2
05D7
04DD
021F
FE75
FBA1
FA9C
FAB5
FAB3
FA55
FA43
FABA
FB14
FAC8
FA5A
FA9A
FB58
FB88
FACC
FA10
FA43
FB0E
FB6A
FB15
FABC
FAD9
FB1E
FB1D
FB03
FB2D
FB6B
FB47
FADB
FAC3
FB16
FB29
FAA9
FA54
FAF0
FBFD
FC3B
FB62
FA8F
FAB2
FB45
FB38
FAC4
FB72
FE1F
01B8
045E
056B
05A6
05CC
05B6
0526
04AC
0514
0631
06D4
0635
04F8
0470
0506
05D4
05D2
050A
0461
046B
04E2
0535
052F
04FB
04BB
0472
0432
0418
041C
0415
0418
0482
0566
0635
0646
05C0
056E
05AD
05FA
05D2
057F
0572
0525
0362
FFEA
FC48
FA63
FA80
FB38
FB5D
FB1A
FB24
FB72
FB77
FB26
FAFF
FB25
FB1D
FA97
FA0B
FA17
FAA4
FB14
FB32
FB63
FBD2
FC0F
FBC3
FB58
FB65
FBB4
FB88
FAB6
FA01
FA0B
FA7B
FA91
FA44
FA47
FAEB
FBA6
FBE6
FBE4
FC13
FC1D
FB41
F9DA
F9AE
FC24
005F
03DB
0506
04B5
04BE
05AB
066C
0616
052B
04C5
051A
056C
0543
0500
050B
051D
04D2
047F
04D9
05D5
067E
062C
056E
054B
05DE
064A
05FF
0575
0554
057C
0559
04E4
04B2
050A
057A
0587
0554
053D
0524
04B4
0434
0453
04ED
049B
0230
FE6F
FB8A
FACC
FB54
FB70
FAB4
FA2A
FA9F
FB7F
FBB1
FB18
FA8F
FAA0
FADE
FAA6
FA1E
F9FE
FA95
FB64
FBC3
FB95
FB2F
FAD9
FA9D
FA76
FA65
FA66
FA6E
FA8A
FACC
FB16
FB27
FB06
FB1B
FBAC
FC5D
FC86
FC19
FBB1
FBA6
FB7D
FABA
FA11
FB02
FE1B
0202
04B1
0575
0548
0547
0582
0578
052C
0515
0538
0503
0442
03A4
03ED
04E6
0593
056E
04F6
04E8
054B
05A1
05BC
05E1
0622
0614
0574
04B8
0493
0512
0581
0556
04D1
0494
04CF
0529
055B
0570
0569
0514
048E
0484
055D
0630
0545
0203
FDFA
FB80
FB52
FC15
FC41
FBD3
FBBE
FC37
FC5F
FBB0
FAD4
FAA2
FADB
FAA1
F9E4
F992
FA39
FB29
FB6C
FB23
FB3B
FBF1
FC64
FBE4
FB07
FAD6
FB60
FBB9
FB53
FAAA
FA79
FAC5
FB0A
FB10
FB0F
FB29
FB36
FB2A
FB2F
FB2D
FAB4
F9DB
F9DB
FC04
0001
03AC
0515
0469
0386
03CF
04E3
0590
056C
051F
053E
058F
058C
053B
0518
055E
05BD
05DB
05C4
05BE
05CE
05B4
0559
04F9
04D3
04D5
04CF
04D0
04FE
053A
0545
053C
0589
062F
067B
05DC
04C9
045C
04E4
0579
054B
04D0
04EE
0530
03E4
0069
FC86
FAA5
FB1A
FC0C
FBEA
FB17
FACB
FB1F
FB27
FA94
FA3E
FABE
FB65
FB3A
FA6D
FA0F
FA9B
FB80
FC0A
FC25
FC07
FBB2
FB23
FAB7
FAD2
FB40
FB67
FB28
FAF8
FB06
FAD9
FA3A
F9EE
FAC7
FC44
FCED
FC26
FB0B
FAFC
FBD9
FC59
FBFB
FBFA
FDD2
0149
0482
05FB
05DF
0566
0558
0590
05A3
058E
0592
05B6
05B6
057E
0559
057F
05A5
055C
04C5
0487
04E7
0559
0530
0480
0408
0440
04DD
054F
0572
0573
055B
051F
0502
054F
05B5
0584
04BD
042D
0426
03E6
02E5
0224
02FD
0481
0366
FD88
F502
EE89
ECB5
EDD7
EEC7
EE7B
EE0A
EE32
EE63
EE14
EDBC
EDFB
EE99
EEF6
EF14
EF73
F017
F061
F019
EFDD
F033
F0AB
F08D
EFF0
EF84
EF88
EF9C
EF7E
EF6D
EFAE
F021
F075
F093
F08F
F063
EFF5
EF69
EF16
EF1C
EF44
EF5C
EF75
EF9D
EFB5
EFC8
F021
F0B7
F0E0
F018
EEDE
EE4F
EED8
EFB3
EFCF
EF03
EE20
EDEA
EE57
EED2
EEFE
EEF3
EEF5
EF1E
