0000
0000
07c0
1ff0
3ff8
3ff8
0ffc
03fc
00fc
03fc
0ffc
3ff8
3ff8
1ff0
07c0
0000
