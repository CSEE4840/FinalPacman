0000
0000
03e0
0ff8
1ffc
1ffc
3ffe
3ffe
3ffe
3ffe
3ffe
1ffc
1ffc
0ff8
03e0
0000
07E0  
0000  
0000  
