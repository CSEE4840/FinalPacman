0000
0000
03e0
0ff8
1ffc
1ffc
3ff0
3fc0
3f00
3fc0
3ff0
1ffc
1ffc
0ff8
03e0
0000
